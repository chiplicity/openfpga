magic
tech sky130A
magscale 1 2
timestamp 1606477073
<< locali >>
rect 7665 18819 7699 18921
rect 12817 18071 12851 18377
rect 15761 18071 15795 18309
rect 16129 17663 16163 17833
rect 12725 17527 12759 17629
rect 4537 17119 4571 17289
rect 18613 15351 18647 15657
rect 16773 14399 16807 14501
rect 13277 13855 13311 14025
rect 18521 13719 18555 13821
rect 16221 13379 16255 13481
rect 19533 13175 19567 13345
rect 6009 12223 6043 12393
rect 11069 12155 11103 12393
rect 8033 11543 8067 11713
rect 14657 10999 14691 11169
rect 18705 10999 18739 11237
rect 14565 10455 14599 10761
rect 19257 10455 19291 10761
rect 14507 10421 14599 10455
rect 3893 9911 3927 10217
rect 5365 10115 5399 10217
rect 16221 9979 16255 10217
rect 8401 8279 8435 8517
rect 10057 8415 10091 8517
rect 7757 7871 7791 8041
<< viali >>
rect 2053 20009 2087 20043
rect 14933 20009 14967 20043
rect 16589 20009 16623 20043
rect 17141 20009 17175 20043
rect 17693 20009 17727 20043
rect 18521 20009 18555 20043
rect 19625 20009 19659 20043
rect 20177 20009 20211 20043
rect 20729 20009 20763 20043
rect 1869 19873 1903 19907
rect 2421 19873 2455 19907
rect 2973 19873 3007 19907
rect 8677 19873 8711 19907
rect 8769 19873 8803 19907
rect 10241 19873 10275 19907
rect 11345 19873 11379 19907
rect 11437 19873 11471 19907
rect 13277 19873 13311 19907
rect 14197 19873 14231 19907
rect 14749 19873 14783 19907
rect 15853 19873 15887 19907
rect 16405 19873 16439 19907
rect 16957 19873 16991 19907
rect 17509 19873 17543 19907
rect 18337 19873 18371 19907
rect 18889 19873 18923 19907
rect 19441 19873 19475 19907
rect 19993 19873 20027 19907
rect 20545 19873 20579 19907
rect 8861 19805 8895 19839
rect 10333 19805 10367 19839
rect 10517 19805 10551 19839
rect 11529 19805 11563 19839
rect 13369 19805 13403 19839
rect 13553 19805 13587 19839
rect 16037 19737 16071 19771
rect 19073 19737 19107 19771
rect 2605 19669 2639 19703
rect 3157 19669 3191 19703
rect 8309 19669 8343 19703
rect 9873 19669 9907 19703
rect 10977 19669 11011 19703
rect 12909 19669 12943 19703
rect 14381 19669 14415 19703
rect 1961 19465 1995 19499
rect 3433 19465 3467 19499
rect 6101 19465 6135 19499
rect 8585 19465 8619 19499
rect 16957 19397 16991 19431
rect 9321 19329 9355 19363
rect 9505 19329 9539 19363
rect 14381 19329 14415 19363
rect 15485 19329 15519 19363
rect 17601 19329 17635 19363
rect 18337 19329 18371 19363
rect 1777 19261 1811 19295
rect 2329 19261 2363 19295
rect 3249 19261 3283 19295
rect 3985 19261 4019 19295
rect 5917 19261 5951 19295
rect 7205 19261 7239 19295
rect 10425 19261 10459 19295
rect 12449 19261 12483 19295
rect 14105 19261 14139 19295
rect 15853 19261 15887 19295
rect 16129 19261 16163 19295
rect 18061 19261 18095 19295
rect 19257 19261 19291 19295
rect 19993 19261 20027 19295
rect 20545 19261 20579 19295
rect 4629 19193 4663 19227
rect 7472 19193 7506 19227
rect 10692 19193 10726 19227
rect 12716 19193 12750 19227
rect 19533 19193 19567 19227
rect 2513 19125 2547 19159
rect 8861 19125 8895 19159
rect 9229 19125 9263 19159
rect 9873 19125 9907 19159
rect 11805 19125 11839 19159
rect 13829 19125 13863 19159
rect 14841 19125 14875 19159
rect 15209 19125 15243 19159
rect 15301 19125 15335 19159
rect 17325 19125 17359 19159
rect 17417 19125 17451 19159
rect 18797 19125 18831 19159
rect 20177 19125 20211 19159
rect 20729 19125 20763 19159
rect 2697 18921 2731 18955
rect 4261 18921 4295 18955
rect 7389 18921 7423 18955
rect 7665 18921 7699 18955
rect 9137 18921 9171 18955
rect 12173 18921 12207 18955
rect 16865 18921 16899 18955
rect 18521 18921 18555 18955
rect 6561 18853 6595 18887
rect 12541 18853 12575 18887
rect 13452 18853 13486 18887
rect 15730 18853 15764 18887
rect 17386 18853 17420 18887
rect 19042 18853 19076 18887
rect 1777 18785 1811 18819
rect 2513 18785 2547 18819
rect 3065 18785 3099 18819
rect 4077 18785 4111 18819
rect 5457 18785 5491 18819
rect 6285 18785 6319 18819
rect 7205 18785 7239 18819
rect 7665 18785 7699 18819
rect 8024 18785 8058 18819
rect 9945 18785 9979 18819
rect 11437 18785 11471 18819
rect 11713 18785 11747 18819
rect 17141 18785 17175 18819
rect 18797 18785 18831 18819
rect 7757 18717 7791 18751
rect 9689 18717 9723 18751
rect 12633 18717 12667 18751
rect 12817 18717 12851 18751
rect 13185 18717 13219 18751
rect 15485 18717 15519 18751
rect 1961 18649 1995 18683
rect 3249 18649 3283 18683
rect 11069 18649 11103 18683
rect 5641 18581 5675 18615
rect 14565 18581 14599 18615
rect 20177 18581 20211 18615
rect 1961 18377 1995 18411
rect 2513 18377 2547 18411
rect 8217 18377 8251 18411
rect 12817 18377 12851 18411
rect 12909 18377 12943 18411
rect 15669 18377 15703 18411
rect 15945 18377 15979 18411
rect 16957 18377 16991 18411
rect 18245 18377 18279 18411
rect 20821 18377 20855 18411
rect 11529 18309 11563 18343
rect 3065 18241 3099 18275
rect 4905 18241 4939 18275
rect 7573 18241 7607 18275
rect 8861 18241 8895 18275
rect 9505 18241 9539 18275
rect 1777 18173 1811 18207
rect 2329 18173 2363 18207
rect 2881 18173 2915 18207
rect 4629 18173 4663 18207
rect 8585 18173 8619 18207
rect 9229 18173 9263 18207
rect 10149 18173 10183 18207
rect 7481 18105 7515 18139
rect 8677 18105 8711 18139
rect 10394 18105 10428 18139
rect 12449 18105 12483 18139
rect 15761 18309 15795 18343
rect 18613 18309 18647 18343
rect 13461 18241 13495 18275
rect 14289 18241 14323 18275
rect 13369 18173 13403 18207
rect 13277 18105 13311 18139
rect 14556 18105 14590 18139
rect 7021 18037 7055 18071
rect 7389 18037 7423 18071
rect 11805 18037 11839 18071
rect 12817 18037 12851 18071
rect 16497 18241 16531 18275
rect 17509 18241 17543 18275
rect 19257 18241 19291 18275
rect 20177 18241 20211 18275
rect 16405 18173 16439 18207
rect 17325 18173 17359 18207
rect 18061 18173 18095 18207
rect 20637 18173 20671 18207
rect 19073 18105 19107 18139
rect 15761 18037 15795 18071
rect 16313 18037 16347 18071
rect 17417 18037 17451 18071
rect 18981 18037 19015 18071
rect 19625 18037 19659 18071
rect 19993 18037 20027 18071
rect 20085 18037 20119 18071
rect 1961 17833 1995 17867
rect 2513 17833 2547 17867
rect 4077 17833 4111 17867
rect 7021 17833 7055 17867
rect 9045 17833 9079 17867
rect 11069 17833 11103 17867
rect 11345 17833 11379 17867
rect 11713 17833 11747 17867
rect 13277 17833 13311 17867
rect 15301 17833 15335 17867
rect 15761 17833 15795 17867
rect 16129 17833 16163 17867
rect 16497 17833 16531 17867
rect 16865 17833 16899 17867
rect 18613 17833 18647 17867
rect 13369 17765 13403 17799
rect 14013 17765 14047 17799
rect 1777 17697 1811 17731
rect 2329 17697 2363 17731
rect 2881 17697 2915 17731
rect 4445 17697 4479 17731
rect 5908 17697 5942 17731
rect 7665 17697 7699 17731
rect 8493 17697 8527 17731
rect 8953 17697 8987 17731
rect 9956 17697 9990 17731
rect 12357 17697 12391 17731
rect 14473 17697 14507 17731
rect 14749 17697 14783 17731
rect 15669 17697 15703 17731
rect 17325 17765 17359 17799
rect 19226 17765 19260 17799
rect 16313 17697 16347 17731
rect 17233 17697 17267 17731
rect 17877 17697 17911 17731
rect 18429 17697 18463 17731
rect 4537 17629 4571 17663
rect 4721 17629 4755 17663
rect 5641 17629 5675 17663
rect 7757 17629 7791 17663
rect 7849 17629 7883 17663
rect 9229 17629 9263 17663
rect 9689 17629 9723 17663
rect 11805 17629 11839 17663
rect 11897 17629 11931 17663
rect 12725 17629 12759 17663
rect 13553 17629 13587 17663
rect 15853 17629 15887 17663
rect 16129 17629 16163 17663
rect 17509 17629 17543 17663
rect 18981 17629 19015 17663
rect 3065 17561 3099 17595
rect 7297 17493 7331 17527
rect 8309 17493 8343 17527
rect 8585 17493 8619 17527
rect 12541 17493 12575 17527
rect 12725 17493 12759 17527
rect 12909 17493 12943 17527
rect 18061 17493 18095 17527
rect 20361 17493 20395 17527
rect 1961 17289 1995 17323
rect 2513 17289 2547 17323
rect 3617 17289 3651 17323
rect 4537 17289 4571 17323
rect 6009 17289 6043 17323
rect 6837 17289 6871 17323
rect 11253 17289 11287 17323
rect 15853 17289 15887 17323
rect 19073 17289 19107 17323
rect 4077 17153 4111 17187
rect 4261 17153 4295 17187
rect 13921 17221 13955 17255
rect 16405 17221 16439 17255
rect 20729 17221 20763 17255
rect 7297 17153 7331 17187
rect 7481 17153 7515 17187
rect 8401 17153 8435 17187
rect 10333 17153 10367 17187
rect 11713 17153 11747 17187
rect 11897 17153 11931 17187
rect 13369 17153 13403 17187
rect 13553 17153 13587 17187
rect 14381 17153 14415 17187
rect 14565 17153 14599 17187
rect 17141 17153 17175 17187
rect 18613 17153 18647 17187
rect 19717 17153 19751 17187
rect 20085 17153 20119 17187
rect 1777 17085 1811 17119
rect 2329 17085 2363 17119
rect 4537 17085 4571 17119
rect 4629 17085 4663 17119
rect 8217 17085 8251 17119
rect 8861 17085 8895 17119
rect 14933 17085 14967 17119
rect 15209 17085 15243 17119
rect 15669 17085 15703 17119
rect 16221 17085 16255 17119
rect 16957 17085 16991 17119
rect 19533 17085 19567 17119
rect 20545 17085 20579 17119
rect 4896 17017 4930 17051
rect 8309 17017 8343 17051
rect 9137 17017 9171 17051
rect 10057 17017 10091 17051
rect 10793 17017 10827 17051
rect 14289 17017 14323 17051
rect 18429 17017 18463 17051
rect 3985 16949 4019 16983
rect 7205 16949 7239 16983
rect 7849 16949 7883 16983
rect 9689 16949 9723 16983
rect 10149 16949 10183 16983
rect 11621 16949 11655 16983
rect 12909 16949 12943 16983
rect 13277 16949 13311 16983
rect 18061 16949 18095 16983
rect 18521 16949 18555 16983
rect 19441 16949 19475 16983
rect 1961 16745 1995 16779
rect 2605 16745 2639 16779
rect 2973 16745 3007 16779
rect 5457 16745 5491 16779
rect 9137 16745 9171 16779
rect 13369 16745 13403 16779
rect 14105 16745 14139 16779
rect 17877 16745 17911 16779
rect 19625 16745 19659 16779
rect 4344 16677 4378 16711
rect 8002 16677 8036 16711
rect 14565 16677 14599 16711
rect 15669 16677 15703 16711
rect 16764 16677 16798 16711
rect 1777 16609 1811 16643
rect 4077 16609 4111 16643
rect 6101 16609 6135 16643
rect 6368 16609 6402 16643
rect 10057 16609 10091 16643
rect 11345 16609 11379 16643
rect 11612 16609 11646 16643
rect 13461 16609 13495 16643
rect 14473 16609 14507 16643
rect 18245 16609 18279 16643
rect 18512 16609 18546 16643
rect 19901 16609 19935 16643
rect 20177 16609 20211 16643
rect 3065 16541 3099 16575
rect 3249 16541 3283 16575
rect 7757 16541 7791 16575
rect 10149 16541 10183 16575
rect 10333 16541 10367 16575
rect 13645 16541 13679 16575
rect 14749 16541 14783 16575
rect 15761 16541 15795 16575
rect 15853 16541 15887 16575
rect 16497 16541 16531 16575
rect 20913 16541 20947 16575
rect 7481 16473 7515 16507
rect 13001 16473 13035 16507
rect 9689 16405 9723 16439
rect 12725 16405 12759 16439
rect 15301 16405 15335 16439
rect 1961 16201 1995 16235
rect 3985 16201 4019 16235
rect 4353 16201 4387 16235
rect 5365 16201 5399 16235
rect 6929 16201 6963 16235
rect 13921 16201 13955 16235
rect 15577 16201 15611 16235
rect 2605 16065 2639 16099
rect 4997 16065 5031 16099
rect 7481 16065 7515 16099
rect 8493 16065 8527 16099
rect 9597 16065 9631 16099
rect 18245 16065 18279 16099
rect 18889 16065 18923 16099
rect 1777 15997 1811 16031
rect 4813 15997 4847 16031
rect 5549 15997 5583 16031
rect 9413 15997 9447 16031
rect 10057 15997 10091 16031
rect 10313 15997 10347 16031
rect 12265 15997 12299 16031
rect 12541 15997 12575 16031
rect 14197 15997 14231 16031
rect 14453 15997 14487 16031
rect 15853 15997 15887 16031
rect 16109 15997 16143 16031
rect 18061 15997 18095 16031
rect 20545 15997 20579 16031
rect 2872 15929 2906 15963
rect 4721 15929 4755 15963
rect 7297 15929 7331 15963
rect 9505 15929 9539 15963
rect 12786 15929 12820 15963
rect 19156 15929 19190 15963
rect 20821 15929 20855 15963
rect 7389 15861 7423 15895
rect 7941 15861 7975 15895
rect 8309 15861 8343 15895
rect 8401 15861 8435 15895
rect 9045 15861 9079 15895
rect 11437 15861 11471 15895
rect 12081 15861 12115 15895
rect 17233 15861 17267 15895
rect 17509 15861 17543 15895
rect 20269 15861 20303 15895
rect 1961 15657 1995 15691
rect 2421 15657 2455 15691
rect 2881 15657 2915 15691
rect 4077 15657 4111 15691
rect 4445 15657 4479 15691
rect 5089 15657 5123 15691
rect 11069 15657 11103 15691
rect 11345 15657 11379 15691
rect 12725 15657 12759 15691
rect 14105 15657 14139 15691
rect 14473 15657 14507 15691
rect 16773 15657 16807 15691
rect 18153 15657 18187 15691
rect 18613 15657 18647 15691
rect 18797 15657 18831 15691
rect 19165 15657 19199 15691
rect 7113 15589 7147 15623
rect 11805 15589 11839 15623
rect 16129 15589 16163 15623
rect 17141 15589 17175 15623
rect 1777 15521 1811 15555
rect 2789 15521 2823 15555
rect 3525 15521 3559 15555
rect 5457 15521 5491 15555
rect 7941 15521 7975 15555
rect 9689 15521 9723 15555
rect 9956 15521 9990 15555
rect 11713 15521 11747 15555
rect 13369 15521 13403 15555
rect 15301 15521 15335 15555
rect 18245 15521 18279 15555
rect 3065 15453 3099 15487
rect 4537 15453 4571 15487
rect 4721 15453 4755 15487
rect 5549 15453 5583 15487
rect 5641 15453 5675 15487
rect 8033 15453 8067 15487
rect 8217 15453 8251 15487
rect 11897 15453 11931 15487
rect 12817 15453 12851 15487
rect 13001 15453 13035 15487
rect 13553 15453 13587 15487
rect 14565 15453 14599 15487
rect 14657 15453 14691 15487
rect 16221 15453 16255 15487
rect 16405 15453 16439 15487
rect 17233 15453 17267 15487
rect 17417 15453 17451 15487
rect 18337 15453 18371 15487
rect 7573 15385 7607 15419
rect 12357 15385 12391 15419
rect 20177 15521 20211 15555
rect 19257 15453 19291 15487
rect 19349 15453 19383 15487
rect 20269 15453 20303 15487
rect 20361 15453 20395 15487
rect 19809 15385 19843 15419
rect 15761 15317 15795 15351
rect 17785 15317 17819 15351
rect 18613 15317 18647 15351
rect 4445 15113 4479 15147
rect 7849 15113 7883 15147
rect 10425 15113 10459 15147
rect 14289 15113 14323 15147
rect 14657 15113 14691 15147
rect 19441 15113 19475 15147
rect 19717 15113 19751 15147
rect 20913 15113 20947 15147
rect 3617 15045 3651 15079
rect 8401 15045 8435 15079
rect 11989 15045 12023 15079
rect 1777 14977 1811 15011
rect 2237 14977 2271 15011
rect 5089 14977 5123 15011
rect 7481 14977 7515 15011
rect 9045 14977 9079 15011
rect 10057 14977 10091 15011
rect 10977 14977 11011 15011
rect 13277 14977 13311 15011
rect 15209 14977 15243 15011
rect 16044 14977 16078 15011
rect 20269 14977 20303 15011
rect 1501 14909 1535 14943
rect 7205 14909 7239 14943
rect 8033 14909 8067 14943
rect 11805 14909 11839 14943
rect 14105 14909 14139 14943
rect 15945 14909 15979 14943
rect 18061 14909 18095 14943
rect 20729 14909 20763 14943
rect 2504 14841 2538 14875
rect 7297 14841 7331 14875
rect 8769 14841 8803 14875
rect 10793 14841 10827 14875
rect 13093 14841 13127 14875
rect 15025 14841 15059 14875
rect 16304 14841 16338 14875
rect 18328 14841 18362 14875
rect 20177 14841 20211 14875
rect 4813 14773 4847 14807
rect 4905 14773 4939 14807
rect 6837 14773 6871 14807
rect 8861 14773 8895 14807
rect 9413 14773 9447 14807
rect 9781 14773 9815 14807
rect 9873 14773 9907 14807
rect 10885 14773 10919 14807
rect 12633 14773 12667 14807
rect 13001 14773 13035 14807
rect 15117 14773 15151 14807
rect 15761 14773 15795 14807
rect 17417 14773 17451 14807
rect 20085 14773 20119 14807
rect 1961 14569 1995 14603
rect 2605 14569 2639 14603
rect 5825 14569 5859 14603
rect 8125 14569 8159 14603
rect 8217 14569 8251 14603
rect 10793 14569 10827 14603
rect 11253 14569 11287 14603
rect 14657 14569 14691 14603
rect 15577 14569 15611 14603
rect 16405 14569 16439 14603
rect 18337 14569 18371 14603
rect 18613 14569 18647 14603
rect 18981 14569 19015 14603
rect 19625 14569 19659 14603
rect 6346 14501 6380 14535
rect 10057 14501 10091 14535
rect 16313 14501 16347 14535
rect 16773 14501 16807 14535
rect 17224 14501 17258 14535
rect 1777 14433 1811 14467
rect 2973 14433 3007 14467
rect 3065 14433 3099 14467
rect 4445 14433 4479 14467
rect 4712 14433 4746 14467
rect 11621 14433 11655 14467
rect 12532 14433 12566 14467
rect 14105 14433 14139 14467
rect 14565 14433 14599 14467
rect 15393 14433 15427 14467
rect 19073 14433 19107 14467
rect 19993 14433 20027 14467
rect 3249 14365 3283 14399
rect 6101 14365 6135 14399
rect 8309 14365 8343 14399
rect 10149 14365 10183 14399
rect 10241 14365 10275 14399
rect 11713 14365 11747 14399
rect 11897 14365 11931 14399
rect 12265 14365 12299 14399
rect 14749 14365 14783 14399
rect 16589 14365 16623 14399
rect 16773 14365 16807 14399
rect 16957 14365 16991 14399
rect 19165 14365 19199 14399
rect 20085 14365 20119 14399
rect 20177 14365 20211 14399
rect 13921 14297 13955 14331
rect 15945 14297 15979 14331
rect 7481 14229 7515 14263
rect 7757 14229 7791 14263
rect 9689 14229 9723 14263
rect 13645 14229 13679 14263
rect 14197 14229 14231 14263
rect 2605 14025 2639 14059
rect 3157 14025 3191 14059
rect 5089 14025 5123 14059
rect 5365 14025 5399 14059
rect 8677 14025 8711 14059
rect 11345 14025 11379 14059
rect 13001 14025 13035 14059
rect 13277 14025 13311 14059
rect 15025 14025 15059 14059
rect 8861 13957 8895 13991
rect 10517 13957 10551 13991
rect 1869 13889 1903 13923
rect 5917 13889 5951 13923
rect 9321 13889 9355 13923
rect 9505 13889 9539 13923
rect 10149 13889 10183 13923
rect 10241 13889 10275 13923
rect 10977 13889 11011 13923
rect 11069 13889 11103 13923
rect 11897 13889 11931 13923
rect 14749 13957 14783 13991
rect 18245 13957 18279 13991
rect 13369 13889 13403 13923
rect 15577 13889 15611 13923
rect 16589 13889 16623 13923
rect 17509 13889 17543 13923
rect 20821 13889 20855 13923
rect 1685 13821 1719 13855
rect 2421 13821 2455 13855
rect 2973 13821 3007 13855
rect 3709 13821 3743 13855
rect 5825 13821 5859 13855
rect 7297 13821 7331 13855
rect 7564 13821 7598 13855
rect 12817 13821 12851 13855
rect 13277 13821 13311 13855
rect 13636 13821 13670 13855
rect 16497 13821 16531 13855
rect 17233 13821 17267 13855
rect 18061 13821 18095 13855
rect 18521 13821 18555 13855
rect 18613 13821 18647 13855
rect 18880 13821 18914 13855
rect 20729 13821 20763 13855
rect 3976 13753 4010 13787
rect 10885 13753 10919 13787
rect 11713 13753 11747 13787
rect 5733 13685 5767 13719
rect 9229 13685 9263 13719
rect 9689 13685 9723 13719
rect 10057 13685 10091 13719
rect 11805 13685 11839 13719
rect 15393 13685 15427 13719
rect 15485 13685 15519 13719
rect 16037 13685 16071 13719
rect 16405 13685 16439 13719
rect 18521 13685 18555 13719
rect 19993 13685 20027 13719
rect 20269 13685 20303 13719
rect 20637 13685 20671 13719
rect 1777 13481 1811 13515
rect 4445 13481 4479 13515
rect 5825 13481 5859 13515
rect 6929 13481 6963 13515
rect 11437 13481 11471 13515
rect 13001 13481 13035 13515
rect 13461 13481 13495 13515
rect 15301 13481 15335 13515
rect 15761 13481 15795 13515
rect 16221 13481 16255 13515
rect 17693 13481 17727 13515
rect 19625 13481 19659 13515
rect 2421 13413 2455 13447
rect 7748 13413 7782 13447
rect 14197 13413 14231 13447
rect 16580 13413 16614 13447
rect 1593 13345 1627 13379
rect 2145 13345 2179 13379
rect 4813 13345 4847 13379
rect 6837 13345 6871 13379
rect 10324 13345 10358 13379
rect 11785 13345 11819 13379
rect 13369 13345 13403 13379
rect 14289 13345 14323 13379
rect 14657 13345 14691 13379
rect 15669 13345 15703 13379
rect 16221 13345 16255 13379
rect 17969 13345 18003 13379
rect 18236 13345 18270 13379
rect 19533 13345 19567 13379
rect 19993 13345 20027 13379
rect 4905 13277 4939 13311
rect 5089 13277 5123 13311
rect 5917 13277 5951 13311
rect 6009 13277 6043 13311
rect 7113 13277 7147 13311
rect 7481 13277 7515 13311
rect 10057 13277 10091 13311
rect 11529 13277 11563 13311
rect 13645 13277 13679 13311
rect 14473 13277 14507 13311
rect 15945 13277 15979 13311
rect 16313 13277 16347 13311
rect 5457 13209 5491 13243
rect 8861 13209 8895 13243
rect 12909 13209 12943 13243
rect 20085 13277 20119 13311
rect 20177 13277 20211 13311
rect 6469 13141 6503 13175
rect 13829 13141 13863 13175
rect 14841 13141 14875 13175
rect 19349 13141 19383 13175
rect 19533 13141 19567 13175
rect 1501 12937 1535 12971
rect 3893 12937 3927 12971
rect 4721 12937 4755 12971
rect 7205 12937 7239 12971
rect 12725 12937 12759 12971
rect 18981 12937 19015 12971
rect 13277 12869 13311 12903
rect 15669 12869 15703 12903
rect 2145 12801 2179 12835
rect 4261 12801 4295 12835
rect 5365 12801 5399 12835
rect 6193 12801 6227 12835
rect 6377 12801 6411 12835
rect 7665 12801 7699 12835
rect 7849 12801 7883 12835
rect 8861 12801 8895 12835
rect 13737 12801 13771 12835
rect 13829 12801 13863 12835
rect 16497 12801 16531 12835
rect 17417 12801 17451 12835
rect 17509 12801 17543 12835
rect 18521 12801 18555 12835
rect 19625 12801 19659 12835
rect 20545 12801 20579 12835
rect 2513 12733 2547 12767
rect 2769 12733 2803 12767
rect 9873 12733 9907 12767
rect 11989 12733 12023 12767
rect 12909 12733 12943 12767
rect 14289 12733 14323 12767
rect 14556 12733 14590 12767
rect 16405 12733 16439 12767
rect 18245 12733 18279 12767
rect 19349 12733 19383 12767
rect 5181 12665 5215 12699
rect 7573 12665 7607 12699
rect 8585 12665 8619 12699
rect 9229 12665 9263 12699
rect 10425 12665 10459 12699
rect 16313 12665 16347 12699
rect 17325 12665 17359 12699
rect 19441 12665 19475 12699
rect 20361 12665 20395 12699
rect 1869 12597 1903 12631
rect 1961 12597 1995 12631
rect 5089 12597 5123 12631
rect 5733 12597 5767 12631
rect 6101 12597 6135 12631
rect 8217 12597 8251 12631
rect 8677 12597 8711 12631
rect 9689 12597 9723 12631
rect 13645 12597 13679 12631
rect 15945 12597 15979 12631
rect 16957 12597 16991 12631
rect 19993 12597 20027 12631
rect 20453 12597 20487 12631
rect 2973 12393 3007 12427
rect 6009 12393 6043 12427
rect 1860 12257 1894 12291
rect 4712 12257 4746 12291
rect 11069 12393 11103 12427
rect 14289 12393 14323 12427
rect 14749 12393 14783 12427
rect 15301 12393 15335 12427
rect 17877 12393 17911 12427
rect 19625 12393 19659 12427
rect 19993 12393 20027 12427
rect 20913 12393 20947 12427
rect 6357 12257 6391 12291
rect 8024 12257 8058 12291
rect 10609 12257 10643 12291
rect 1593 12189 1627 12223
rect 4445 12189 4479 12223
rect 6009 12189 6043 12223
rect 6101 12189 6135 12223
rect 7757 12189 7791 12223
rect 10701 12189 10735 12223
rect 10885 12189 10919 12223
rect 16764 12325 16798 12359
rect 11520 12257 11554 12291
rect 13176 12257 13210 12291
rect 15669 12257 15703 12291
rect 18981 12257 19015 12291
rect 11253 12189 11287 12223
rect 12909 12189 12943 12223
rect 15761 12189 15795 12223
rect 15853 12189 15887 12223
rect 16497 12189 16531 12223
rect 19073 12189 19107 12223
rect 19257 12189 19291 12223
rect 20085 12189 20119 12223
rect 20177 12189 20211 12223
rect 7481 12121 7515 12155
rect 11069 12121 11103 12155
rect 12633 12121 12667 12155
rect 18613 12121 18647 12155
rect 5825 12053 5859 12087
rect 9137 12053 9171 12087
rect 10241 12053 10275 12087
rect 2145 11849 2179 11883
rect 4169 11849 4203 11883
rect 14749 11849 14783 11883
rect 18613 11849 18647 11883
rect 7205 11781 7239 11815
rect 2697 11713 2731 11747
rect 3801 11713 3835 11747
rect 4813 11713 4847 11747
rect 5733 11713 5767 11747
rect 7849 11713 7883 11747
rect 8033 11713 8067 11747
rect 10609 11713 10643 11747
rect 11621 11713 11655 11747
rect 13093 11713 13127 11747
rect 15301 11713 15335 11747
rect 19533 11713 19567 11747
rect 20545 11713 20579 11747
rect 2605 11645 2639 11679
rect 3525 11645 3559 11679
rect 6653 11645 6687 11679
rect 7573 11645 7607 11679
rect 3617 11577 3651 11611
rect 7665 11577 7699 11611
rect 8217 11645 8251 11679
rect 8484 11645 8518 11679
rect 10425 11645 10459 11679
rect 11437 11645 11471 11679
rect 13360 11645 13394 11679
rect 15117 11645 15151 11679
rect 16044 11645 16078 11679
rect 18429 11645 18463 11679
rect 19349 11645 19383 11679
rect 11529 11577 11563 11611
rect 15209 11577 15243 11611
rect 16304 11577 16338 11611
rect 19441 11577 19475 11611
rect 20361 11577 20395 11611
rect 2513 11509 2547 11543
rect 3157 11509 3191 11543
rect 4537 11509 4571 11543
rect 4629 11509 4663 11543
rect 5181 11509 5215 11543
rect 5549 11509 5583 11543
rect 5641 11509 5675 11543
rect 6469 11509 6503 11543
rect 8033 11509 8067 11543
rect 9597 11509 9631 11543
rect 10057 11509 10091 11543
rect 10517 11509 10551 11543
rect 11069 11509 11103 11543
rect 14473 11509 14507 11543
rect 17417 11509 17451 11543
rect 18981 11509 19015 11543
rect 19993 11509 20027 11543
rect 20453 11509 20487 11543
rect 2881 11305 2915 11339
rect 5733 11305 5767 11339
rect 6193 11305 6227 11339
rect 6745 11305 6779 11339
rect 8953 11305 8987 11339
rect 10425 11305 10459 11339
rect 12633 11305 12667 11339
rect 13277 11305 13311 11339
rect 13645 11305 13679 11339
rect 14749 11305 14783 11339
rect 16681 11305 16715 11339
rect 17325 11305 17359 11339
rect 18521 11305 18555 11339
rect 18889 11305 18923 11339
rect 20913 11305 20947 11339
rect 7113 11237 7147 11271
rect 12725 11237 12759 11271
rect 17417 11237 17451 11271
rect 18705 11237 18739 11271
rect 19257 11237 19291 11271
rect 20269 11237 20303 11271
rect 1768 11169 1802 11203
rect 4077 11169 4111 11203
rect 4344 11169 4378 11203
rect 6101 11169 6135 11203
rect 7205 11169 7239 11203
rect 10793 11169 10827 11203
rect 12173 11169 12207 11203
rect 14473 11169 14507 11203
rect 14657 11169 14691 11203
rect 15557 11169 15591 11203
rect 18325 11169 18359 11203
rect 1501 11101 1535 11135
rect 6285 11101 6319 11135
rect 7297 11101 7331 11135
rect 9045 11101 9079 11135
rect 9137 11101 9171 11135
rect 10885 11101 10919 11135
rect 11069 11101 11103 11135
rect 12817 11101 12851 11135
rect 13737 11101 13771 11135
rect 13829 11101 13863 11135
rect 11989 11033 12023 11067
rect 12265 11033 12299 11067
rect 14289 11033 14323 11067
rect 15301 11101 15335 11135
rect 17509 11101 17543 11135
rect 19349 11169 19383 11203
rect 19993 11169 20027 11203
rect 19533 11101 19567 11135
rect 5457 10965 5491 10999
rect 8585 10965 8619 10999
rect 14657 10965 14691 10999
rect 16957 10965 16991 10999
rect 18705 10965 18739 10999
rect 1685 10761 1719 10795
rect 3893 10761 3927 10795
rect 8677 10761 8711 10795
rect 12081 10761 12115 10795
rect 14565 10761 14599 10795
rect 14933 10761 14967 10795
rect 18429 10761 18463 10795
rect 19257 10761 19291 10795
rect 2329 10625 2363 10659
rect 3341 10625 3375 10659
rect 4537 10625 4571 10659
rect 5549 10625 5583 10659
rect 7849 10625 7883 10659
rect 9137 10625 9171 10659
rect 9229 10625 9263 10659
rect 10241 10625 10275 10659
rect 10701 10625 10735 10659
rect 12909 10625 12943 10659
rect 13001 10625 13035 10659
rect 14197 10625 14231 10659
rect 4353 10557 4387 10591
rect 8493 10557 8527 10591
rect 10057 10557 10091 10591
rect 10149 10557 10183 10591
rect 10968 10557 11002 10591
rect 14013 10557 14047 10591
rect 2053 10489 2087 10523
rect 3157 10489 3191 10523
rect 5365 10489 5399 10523
rect 9045 10489 9079 10523
rect 15485 10625 15519 10659
rect 16773 10625 16807 10659
rect 18981 10625 19015 10659
rect 14841 10557 14875 10591
rect 15301 10557 15335 10591
rect 16497 10557 16531 10591
rect 18797 10557 18831 10591
rect 16589 10489 16623 10523
rect 19993 10625 20027 10659
rect 20453 10557 20487 10591
rect 19809 10489 19843 10523
rect 20729 10489 20763 10523
rect 2145 10421 2179 10455
rect 2697 10421 2731 10455
rect 3065 10421 3099 10455
rect 4261 10421 4295 10455
rect 4905 10421 4939 10455
rect 5273 10421 5307 10455
rect 7297 10421 7331 10455
rect 7665 10421 7699 10455
rect 7757 10421 7791 10455
rect 8309 10421 8343 10455
rect 9689 10421 9723 10455
rect 12449 10421 12483 10455
rect 12817 10421 12851 10455
rect 13645 10421 13679 10455
rect 14105 10421 14139 10455
rect 14473 10421 14507 10455
rect 14657 10421 14691 10455
rect 15393 10421 15427 10455
rect 16129 10421 16163 10455
rect 18889 10421 18923 10455
rect 19257 10421 19291 10455
rect 19441 10421 19475 10455
rect 19901 10421 19935 10455
rect 1869 10217 1903 10251
rect 2237 10217 2271 10251
rect 3893 10217 3927 10251
rect 4077 10217 4111 10251
rect 5089 10217 5123 10251
rect 5365 10217 5399 10251
rect 6837 10217 6871 10251
rect 7481 10217 7515 10251
rect 9321 10217 9355 10251
rect 9689 10217 9723 10251
rect 10149 10217 10183 10251
rect 12909 10217 12943 10251
rect 13369 10217 13403 10251
rect 14657 10217 14691 10251
rect 16221 10217 16255 10251
rect 18153 10217 18187 10251
rect 20177 10217 20211 10251
rect 1409 10149 1443 10183
rect 2881 10081 2915 10115
rect 3525 10081 3559 10115
rect 2329 10013 2363 10047
rect 2513 10013 2547 10047
rect 3065 9945 3099 9979
rect 14565 10149 14599 10183
rect 4445 10081 4479 10115
rect 4537 10081 4571 10115
rect 5273 10081 5307 10115
rect 5365 10081 5399 10115
rect 5457 10081 5491 10115
rect 5724 10081 5758 10115
rect 8197 10081 8231 10115
rect 10057 10081 10091 10115
rect 11253 10081 11287 10115
rect 11509 10081 11543 10115
rect 13277 10081 13311 10115
rect 15669 10081 15703 10115
rect 4629 10013 4663 10047
rect 7941 10013 7975 10047
rect 10241 10013 10275 10047
rect 13553 10013 13587 10047
rect 14841 10013 14875 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 16569 10081 16603 10115
rect 17969 10081 18003 10115
rect 18889 10081 18923 10115
rect 18981 10081 19015 10115
rect 20085 10081 20119 10115
rect 16313 10013 16347 10047
rect 19165 10013 19199 10047
rect 20361 10013 20395 10047
rect 16221 9945 16255 9979
rect 17693 9945 17727 9979
rect 3893 9877 3927 9911
rect 12633 9877 12667 9911
rect 14197 9877 14231 9911
rect 15301 9877 15335 9911
rect 18521 9877 18555 9911
rect 19717 9877 19751 9911
rect 16221 9673 16255 9707
rect 4077 9605 4111 9639
rect 18153 9605 18187 9639
rect 1961 9537 1995 9571
rect 4997 9537 5031 9571
rect 6009 9537 6043 9571
rect 7573 9537 7607 9571
rect 9965 9537 9999 9571
rect 13093 9537 13127 9571
rect 13461 9537 13495 9571
rect 14841 9537 14875 9571
rect 17049 9537 17083 9571
rect 18613 9537 18647 9571
rect 18797 9537 18831 9571
rect 19809 9537 19843 9571
rect 20729 9537 20763 9571
rect 1777 9469 1811 9503
rect 2697 9469 2731 9503
rect 4721 9469 4755 9503
rect 5825 9469 5859 9503
rect 7829 9469 7863 9503
rect 10232 9469 10266 9503
rect 20637 9469 20671 9503
rect 2942 9401 2976 9435
rect 15086 9401 15120 9435
rect 16865 9401 16899 9435
rect 18521 9401 18555 9435
rect 4353 9333 4387 9367
rect 4813 9333 4847 9367
rect 5365 9333 5399 9367
rect 5733 9333 5767 9367
rect 8953 9333 8987 9367
rect 11345 9333 11379 9367
rect 12449 9333 12483 9367
rect 12817 9333 12851 9367
rect 12909 9333 12943 9367
rect 14381 9333 14415 9367
rect 16497 9333 16531 9367
rect 16957 9333 16991 9367
rect 19165 9333 19199 9367
rect 19533 9333 19567 9367
rect 19625 9333 19659 9367
rect 20177 9333 20211 9367
rect 20545 9333 20579 9367
rect 2237 9129 2271 9163
rect 4445 9129 4479 9163
rect 4813 9129 4847 9163
rect 5457 9129 5491 9163
rect 7113 9129 7147 9163
rect 8125 9129 8159 9163
rect 8493 9129 8527 9163
rect 10149 9129 10183 9163
rect 10793 9129 10827 9163
rect 13277 9129 13311 9163
rect 14933 9129 14967 9163
rect 15301 9129 15335 9163
rect 15669 9129 15703 9163
rect 16773 9129 16807 9163
rect 20913 9129 20947 9163
rect 1777 9061 1811 9095
rect 5917 9061 5951 9095
rect 7573 9061 7607 9095
rect 10057 9061 10091 9095
rect 11253 9061 11287 9095
rect 13820 9061 13854 9095
rect 18512 9061 18546 9095
rect 20177 9061 20211 9095
rect 1501 8993 1535 9027
rect 2605 8993 2639 9027
rect 5825 8993 5859 9027
rect 7481 8993 7515 9027
rect 8585 8993 8619 9027
rect 11161 8993 11195 9027
rect 12153 8993 12187 9027
rect 16681 8993 16715 9027
rect 19901 8993 19935 9027
rect 2697 8925 2731 8959
rect 2881 8925 2915 8959
rect 4905 8925 4939 8959
rect 5089 8925 5123 8959
rect 6101 8925 6135 8959
rect 7665 8925 7699 8959
rect 8769 8925 8803 8959
rect 10241 8925 10275 8959
rect 11437 8925 11471 8959
rect 11897 8925 11931 8959
rect 13553 8925 13587 8959
rect 15761 8925 15795 8959
rect 15853 8925 15887 8959
rect 16957 8925 16991 8959
rect 18245 8925 18279 8959
rect 9689 8857 9723 8891
rect 16313 8789 16347 8823
rect 19625 8789 19659 8823
rect 2881 8585 2915 8619
rect 3157 8585 3191 8619
rect 4353 8585 4387 8619
rect 5365 8585 5399 8619
rect 10241 8585 10275 8619
rect 14749 8585 14783 8619
rect 15761 8585 15795 8619
rect 16957 8585 16991 8619
rect 19441 8585 19475 8619
rect 19717 8585 19751 8619
rect 20913 8585 20947 8619
rect 7573 8517 7607 8551
rect 8401 8517 8435 8551
rect 9965 8517 9999 8551
rect 10057 8517 10091 8551
rect 11253 8517 11287 8551
rect 3709 8449 3743 8483
rect 4813 8449 4847 8483
rect 4997 8449 5031 8483
rect 5825 8449 5859 8483
rect 6009 8449 6043 8483
rect 8125 8449 8159 8483
rect 1501 8381 1535 8415
rect 1768 8381 1802 8415
rect 3617 8381 3651 8415
rect 4721 8313 4755 8347
rect 5733 8313 5767 8347
rect 7941 8313 7975 8347
rect 8033 8313 8067 8347
rect 10793 8449 10827 8483
rect 11713 8449 11747 8483
rect 11805 8449 11839 8483
rect 12449 8449 12483 8483
rect 15301 8449 15335 8483
rect 16405 8449 16439 8483
rect 17509 8449 17543 8483
rect 20177 8449 20211 8483
rect 20269 8449 20303 8483
rect 8585 8381 8619 8415
rect 10057 8381 10091 8415
rect 10609 8381 10643 8415
rect 16129 8381 16163 8415
rect 18061 8381 18095 8415
rect 20085 8381 20119 8415
rect 20729 8381 20763 8415
rect 8852 8313 8886 8347
rect 12716 8313 12750 8347
rect 15209 8313 15243 8347
rect 16221 8313 16255 8347
rect 17325 8313 17359 8347
rect 18328 8313 18362 8347
rect 3525 8245 3559 8279
rect 8401 8245 8435 8279
rect 10701 8245 10735 8279
rect 11621 8245 11655 8279
rect 13829 8245 13863 8279
rect 15117 8245 15151 8279
rect 17417 8245 17451 8279
rect 2605 8041 2639 8075
rect 4077 8041 4111 8075
rect 4537 8041 4571 8075
rect 7113 8041 7147 8075
rect 7757 8041 7791 8075
rect 9229 8041 9263 8075
rect 9965 8041 9999 8075
rect 12357 8041 12391 8075
rect 18245 8041 18279 8075
rect 19441 8041 19475 8075
rect 19809 8041 19843 8075
rect 3065 7973 3099 8007
rect 2973 7905 3007 7939
rect 4445 7905 4479 7939
rect 5989 7905 6023 7939
rect 8116 7905 8150 7939
rect 10333 7905 10367 7939
rect 10425 7905 10459 7939
rect 12725 7905 12759 7939
rect 16865 7905 16899 7939
rect 17132 7905 17166 7939
rect 3157 7837 3191 7871
rect 4629 7837 4663 7871
rect 5733 7837 5767 7871
rect 7757 7837 7791 7871
rect 7849 7837 7883 7871
rect 10517 7837 10551 7871
rect 12817 7837 12851 7871
rect 12909 7837 12943 7871
rect 19901 7837 19935 7871
rect 19993 7837 20027 7871
rect 1501 7497 1535 7531
rect 3893 7497 3927 7531
rect 6377 7497 6411 7531
rect 8309 7497 8343 7531
rect 8585 7497 8619 7531
rect 16405 7497 16439 7531
rect 18061 7497 18095 7531
rect 19901 7497 19935 7531
rect 2145 7361 2179 7395
rect 6929 7361 6963 7395
rect 9137 7361 9171 7395
rect 17049 7361 17083 7395
rect 18613 7361 18647 7395
rect 19349 7361 19383 7395
rect 20453 7361 20487 7395
rect 2513 7293 2547 7327
rect 2780 7293 2814 7327
rect 4997 7293 5031 7327
rect 5264 7293 5298 7327
rect 16865 7293 16899 7327
rect 19165 7293 19199 7327
rect 1961 7225 1995 7259
rect 7174 7225 7208 7259
rect 8953 7225 8987 7259
rect 16773 7225 16807 7259
rect 18429 7225 18463 7259
rect 20269 7225 20303 7259
rect 1869 7157 1903 7191
rect 4537 7157 4571 7191
rect 9045 7157 9079 7191
rect 18521 7157 18555 7191
rect 20361 7157 20395 7191
rect 18061 6953 18095 6987
rect 4537 6885 4571 6919
rect 1860 6817 1894 6851
rect 5549 6817 5583 6851
rect 6561 6817 6595 6851
rect 7573 6817 7607 6851
rect 7665 6817 7699 6851
rect 16681 6817 16715 6851
rect 16948 6817 16982 6851
rect 19432 6817 19466 6851
rect 1593 6749 1627 6783
rect 3341 6749 3375 6783
rect 4629 6749 4663 6783
rect 4813 6749 4847 6783
rect 5641 6749 5675 6783
rect 5733 6749 5767 6783
rect 6653 6749 6687 6783
rect 6837 6749 6871 6783
rect 7849 6749 7883 6783
rect 19165 6749 19199 6783
rect 20913 6749 20947 6783
rect 2973 6681 3007 6715
rect 4169 6681 4203 6715
rect 7205 6681 7239 6715
rect 5181 6613 5215 6647
rect 6193 6613 6227 6647
rect 20545 6613 20579 6647
rect 2973 6409 3007 6443
rect 4997 6409 5031 6443
rect 20729 6409 20763 6443
rect 3617 6273 3651 6307
rect 5549 6273 5583 6307
rect 19349 6273 19383 6307
rect 3341 6205 3375 6239
rect 5365 6205 5399 6239
rect 19616 6137 19650 6171
rect 3433 6069 3467 6103
rect 5457 6069 5491 6103
rect 19809 5865 19843 5899
rect 20177 5865 20211 5899
rect 20269 5661 20303 5695
rect 20361 5661 20395 5695
rect 20085 5321 20119 5355
rect 20637 5185 20671 5219
rect 19901 4981 19935 5015
rect 20453 4981 20487 5015
rect 20545 4981 20579 5015
rect 4997 3009 5031 3043
rect 5825 3009 5859 3043
rect 15485 3009 15519 3043
rect 4721 2941 4755 2975
rect 5641 2941 5675 2975
rect 15209 2941 15243 2975
<< metal1 >>
rect 3694 20952 3700 21004
rect 3752 20992 3758 21004
rect 6086 20992 6092 21004
rect 3752 20964 6092 20992
rect 3752 20952 3758 20964
rect 6086 20952 6092 20964
rect 6144 20952 6150 21004
rect 14366 20272 14372 20324
rect 14424 20312 14430 20324
rect 14918 20312 14924 20324
rect 14424 20284 14924 20312
rect 14424 20272 14430 20284
rect 14918 20272 14924 20284
rect 14976 20272 14982 20324
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 2041 20043 2099 20049
rect 2041 20009 2053 20043
rect 2087 20040 2099 20043
rect 2774 20040 2780 20052
rect 2087 20012 2780 20040
rect 2087 20009 2099 20012
rect 2041 20003 2099 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 11146 20000 11152 20052
rect 11204 20000 11210 20052
rect 11606 20000 11612 20052
rect 11664 20040 11670 20052
rect 12158 20040 12164 20052
rect 11664 20012 12164 20040
rect 11664 20000 11670 20012
rect 12158 20000 12164 20012
rect 12216 20000 12222 20052
rect 12710 20000 12716 20052
rect 12768 20040 12774 20052
rect 13262 20040 13268 20052
rect 12768 20012 13268 20040
rect 12768 20000 12774 20012
rect 13262 20000 13268 20012
rect 13320 20000 13326 20052
rect 14921 20043 14979 20049
rect 14921 20009 14933 20043
rect 14967 20009 14979 20043
rect 14921 20003 14979 20009
rect 16577 20043 16635 20049
rect 16577 20009 16589 20043
rect 16623 20040 16635 20043
rect 17034 20040 17040 20052
rect 16623 20012 17040 20040
rect 16623 20009 16635 20012
rect 16577 20003 16635 20009
rect 198 19932 204 19984
rect 256 19972 262 19984
rect 256 19944 2452 19972
rect 256 19932 262 19944
rect 2424 19913 2452 19944
rect 2498 19932 2504 19984
rect 2556 19972 2562 19984
rect 3234 19972 3240 19984
rect 2556 19944 3240 19972
rect 2556 19932 2562 19944
rect 3234 19932 3240 19944
rect 3292 19932 3298 19984
rect 11164 19972 11192 20000
rect 12434 19972 12440 19984
rect 11164 19944 12440 19972
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 14936 19972 14964 20003
rect 17034 20000 17040 20012
rect 17092 20000 17098 20052
rect 17129 20043 17187 20049
rect 17129 20009 17141 20043
rect 17175 20040 17187 20043
rect 17494 20040 17500 20052
rect 17175 20012 17500 20040
rect 17175 20009 17187 20012
rect 17129 20003 17187 20009
rect 17494 20000 17500 20012
rect 17552 20000 17558 20052
rect 17681 20043 17739 20049
rect 17681 20009 17693 20043
rect 17727 20040 17739 20043
rect 18322 20040 18328 20052
rect 17727 20012 18328 20040
rect 17727 20009 17739 20012
rect 17681 20003 17739 20009
rect 18322 20000 18328 20012
rect 18380 20000 18386 20052
rect 18509 20043 18567 20049
rect 18509 20009 18521 20043
rect 18555 20040 18567 20043
rect 18782 20040 18788 20052
rect 18555 20012 18788 20040
rect 18555 20009 18567 20012
rect 18509 20003 18567 20009
rect 18782 20000 18788 20012
rect 18840 20000 18846 20052
rect 19610 20040 19616 20052
rect 19571 20012 19616 20040
rect 19610 20000 19616 20012
rect 19668 20000 19674 20052
rect 20162 20040 20168 20052
rect 20123 20012 20168 20040
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 20717 20043 20775 20049
rect 20717 20040 20729 20043
rect 20680 20012 20729 20040
rect 20680 20000 20686 20012
rect 20717 20009 20729 20012
rect 20763 20009 20775 20043
rect 20717 20003 20775 20009
rect 17862 19972 17868 19984
rect 14936 19944 17868 19972
rect 17862 19932 17868 19944
rect 17920 19932 17926 19984
rect 1857 19907 1915 19913
rect 1857 19873 1869 19907
rect 1903 19873 1915 19907
rect 1857 19867 1915 19873
rect 2409 19907 2467 19913
rect 2409 19873 2421 19907
rect 2455 19873 2467 19907
rect 2409 19867 2467 19873
rect 2961 19907 3019 19913
rect 2961 19873 2973 19907
rect 3007 19904 3019 19907
rect 3326 19904 3332 19916
rect 3007 19876 3332 19904
rect 3007 19873 3019 19876
rect 2961 19867 3019 19873
rect 1872 19768 1900 19867
rect 3326 19864 3332 19876
rect 3384 19864 3390 19916
rect 8478 19864 8484 19916
rect 8536 19904 8542 19916
rect 8665 19907 8723 19913
rect 8665 19904 8677 19907
rect 8536 19876 8677 19904
rect 8536 19864 8542 19876
rect 8665 19873 8677 19876
rect 8711 19873 8723 19907
rect 8665 19867 8723 19873
rect 8757 19907 8815 19913
rect 8757 19873 8769 19907
rect 8803 19904 8815 19907
rect 9582 19904 9588 19916
rect 8803 19876 9588 19904
rect 8803 19873 8815 19876
rect 8757 19867 8815 19873
rect 9582 19864 9588 19876
rect 9640 19864 9646 19916
rect 10229 19907 10287 19913
rect 10229 19904 10241 19907
rect 9692 19876 10241 19904
rect 3142 19796 3148 19848
rect 3200 19836 3206 19848
rect 3694 19836 3700 19848
rect 3200 19808 3700 19836
rect 3200 19796 3206 19808
rect 3694 19796 3700 19808
rect 3752 19796 3758 19848
rect 8846 19836 8852 19848
rect 8807 19808 8852 19836
rect 8846 19796 8852 19808
rect 8904 19796 8910 19848
rect 4154 19768 4160 19780
rect 1872 19740 4160 19768
rect 4154 19728 4160 19740
rect 4212 19728 4218 19780
rect 7558 19728 7564 19780
rect 7616 19768 7622 19780
rect 9692 19768 9720 19876
rect 10229 19873 10241 19876
rect 10275 19904 10287 19907
rect 10410 19904 10416 19916
rect 10275 19876 10416 19904
rect 10275 19873 10287 19876
rect 10229 19867 10287 19873
rect 10410 19864 10416 19876
rect 10468 19864 10474 19916
rect 11146 19864 11152 19916
rect 11204 19904 11210 19916
rect 11333 19907 11391 19913
rect 11333 19904 11345 19907
rect 11204 19876 11345 19904
rect 11204 19864 11210 19876
rect 11333 19873 11345 19876
rect 11379 19873 11391 19907
rect 11333 19867 11391 19873
rect 11425 19907 11483 19913
rect 11425 19873 11437 19907
rect 11471 19904 11483 19907
rect 11606 19904 11612 19916
rect 11471 19876 11612 19904
rect 11471 19873 11483 19876
rect 11425 19867 11483 19873
rect 11606 19864 11612 19876
rect 11664 19864 11670 19916
rect 13262 19904 13268 19916
rect 13223 19876 13268 19904
rect 13262 19864 13268 19876
rect 13320 19864 13326 19916
rect 14182 19904 14188 19916
rect 14143 19876 14188 19904
rect 14182 19864 14188 19876
rect 14240 19864 14246 19916
rect 14734 19904 14740 19916
rect 14695 19876 14740 19904
rect 14734 19864 14740 19876
rect 14792 19864 14798 19916
rect 15010 19864 15016 19916
rect 15068 19904 15074 19916
rect 15841 19907 15899 19913
rect 15841 19904 15853 19907
rect 15068 19876 15853 19904
rect 15068 19864 15074 19876
rect 15841 19873 15853 19876
rect 15887 19873 15899 19907
rect 15841 19867 15899 19873
rect 16022 19864 16028 19916
rect 16080 19904 16086 19916
rect 16393 19907 16451 19913
rect 16393 19904 16405 19907
rect 16080 19876 16405 19904
rect 16080 19864 16086 19876
rect 16393 19873 16405 19876
rect 16439 19873 16451 19907
rect 16393 19867 16451 19873
rect 16758 19864 16764 19916
rect 16816 19904 16822 19916
rect 16945 19907 17003 19913
rect 16945 19904 16957 19907
rect 16816 19876 16957 19904
rect 16816 19864 16822 19876
rect 16945 19873 16957 19876
rect 16991 19873 17003 19907
rect 16945 19867 17003 19873
rect 17497 19907 17555 19913
rect 17497 19873 17509 19907
rect 17543 19873 17555 19907
rect 17497 19867 17555 19873
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18506 19904 18512 19916
rect 18371 19876 18512 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 9950 19796 9956 19848
rect 10008 19836 10014 19848
rect 10321 19839 10379 19845
rect 10321 19836 10333 19839
rect 10008 19808 10333 19836
rect 10008 19796 10014 19808
rect 10321 19805 10333 19808
rect 10367 19805 10379 19839
rect 10502 19836 10508 19848
rect 10463 19808 10508 19836
rect 10321 19799 10379 19805
rect 10502 19796 10508 19808
rect 10560 19796 10566 19848
rect 11517 19839 11575 19845
rect 11517 19805 11529 19839
rect 11563 19836 11575 19839
rect 11790 19836 11796 19848
rect 11563 19808 11796 19836
rect 11563 19805 11575 19808
rect 11517 19799 11575 19805
rect 11790 19796 11796 19808
rect 11848 19796 11854 19848
rect 13354 19836 13360 19848
rect 13315 19808 13360 19836
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 13538 19836 13544 19848
rect 13499 19808 13544 19836
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 16574 19796 16580 19848
rect 16632 19836 16638 19848
rect 17512 19836 17540 19867
rect 18506 19864 18512 19876
rect 18564 19864 18570 19916
rect 18877 19907 18935 19913
rect 18877 19873 18889 19907
rect 18923 19873 18935 19907
rect 19426 19904 19432 19916
rect 19387 19876 19432 19904
rect 18877 19867 18935 19873
rect 16632 19808 17540 19836
rect 16632 19796 16638 19808
rect 17954 19796 17960 19848
rect 18012 19836 18018 19848
rect 18892 19836 18920 19867
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 19536 19876 19993 19904
rect 18012 19808 18920 19836
rect 18012 19796 18018 19808
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 19536 19836 19564 19876
rect 19981 19873 19993 19876
rect 20027 19873 20039 19907
rect 19981 19867 20039 19873
rect 20533 19907 20591 19913
rect 20533 19873 20545 19907
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 19392 19808 19564 19836
rect 19392 19796 19398 19808
rect 19610 19796 19616 19848
rect 19668 19836 19674 19848
rect 20548 19836 20576 19867
rect 19668 19808 20576 19836
rect 19668 19796 19674 19808
rect 7616 19740 9720 19768
rect 16025 19771 16083 19777
rect 7616 19728 7622 19740
rect 16025 19737 16037 19771
rect 16071 19768 16083 19771
rect 16666 19768 16672 19780
rect 16071 19740 16672 19768
rect 16071 19737 16083 19740
rect 16025 19731 16083 19737
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 19058 19768 19064 19780
rect 19019 19740 19064 19768
rect 19058 19728 19064 19740
rect 19116 19728 19122 19780
rect 2590 19700 2596 19712
rect 2551 19672 2596 19700
rect 2590 19660 2596 19672
rect 2648 19660 2654 19712
rect 3142 19700 3148 19712
rect 3103 19672 3148 19700
rect 3142 19660 3148 19672
rect 3200 19660 3206 19712
rect 8294 19700 8300 19712
rect 8255 19672 8300 19700
rect 8294 19660 8300 19672
rect 8352 19660 8358 19712
rect 9490 19660 9496 19712
rect 9548 19700 9554 19712
rect 9861 19703 9919 19709
rect 9861 19700 9873 19703
rect 9548 19672 9873 19700
rect 9548 19660 9554 19672
rect 9861 19669 9873 19672
rect 9907 19669 9919 19703
rect 9861 19663 9919 19669
rect 10965 19703 11023 19709
rect 10965 19669 10977 19703
rect 11011 19700 11023 19703
rect 11054 19700 11060 19712
rect 11011 19672 11060 19700
rect 11011 19669 11023 19672
rect 10965 19663 11023 19669
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 12897 19703 12955 19709
rect 12897 19669 12909 19703
rect 12943 19700 12955 19703
rect 14090 19700 14096 19712
rect 12943 19672 14096 19700
rect 12943 19669 12955 19672
rect 12897 19663 12955 19669
rect 14090 19660 14096 19672
rect 14148 19660 14154 19712
rect 14369 19703 14427 19709
rect 14369 19669 14381 19703
rect 14415 19700 14427 19703
rect 18598 19700 18604 19712
rect 14415 19672 18604 19700
rect 14415 19669 14427 19672
rect 14369 19663 14427 19669
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 3418 19496 3424 19508
rect 3379 19468 3424 19496
rect 3418 19456 3424 19468
rect 3476 19456 3482 19508
rect 6086 19496 6092 19508
rect 6047 19468 6092 19496
rect 6086 19456 6092 19468
rect 6144 19456 6150 19508
rect 8573 19499 8631 19505
rect 8573 19465 8585 19499
rect 8619 19496 8631 19499
rect 8846 19496 8852 19508
rect 8619 19468 8852 19496
rect 8619 19465 8631 19468
rect 8573 19459 8631 19465
rect 8846 19456 8852 19468
rect 8904 19456 8910 19508
rect 9950 19496 9956 19508
rect 8956 19468 9956 19496
rect 8956 19428 8984 19468
rect 9950 19456 9956 19468
rect 10008 19456 10014 19508
rect 8220 19400 8984 19428
rect 3804 19332 4108 19360
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 2130 19292 2136 19304
rect 1811 19264 2136 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 2130 19252 2136 19264
rect 2188 19252 2194 19304
rect 2314 19292 2320 19304
rect 2275 19264 2320 19292
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 3237 19295 3295 19301
rect 3237 19261 3249 19295
rect 3283 19292 3295 19295
rect 3804 19292 3832 19332
rect 3970 19292 3976 19304
rect 3283 19264 3832 19292
rect 3931 19264 3976 19292
rect 3283 19261 3295 19264
rect 3237 19255 3295 19261
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 4080 19292 4108 19332
rect 5534 19292 5540 19304
rect 4080 19264 5540 19292
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 5902 19292 5908 19304
rect 5863 19264 5908 19292
rect 5902 19252 5908 19264
rect 5960 19252 5966 19304
rect 7193 19295 7251 19301
rect 7193 19261 7205 19295
rect 7239 19261 7251 19295
rect 7193 19255 7251 19261
rect 1026 19184 1032 19236
rect 1084 19224 1090 19236
rect 4617 19227 4675 19233
rect 1084 19196 4200 19224
rect 1084 19184 1090 19196
rect 4172 19168 4200 19196
rect 4617 19193 4629 19227
rect 4663 19224 4675 19227
rect 6638 19224 6644 19236
rect 4663 19196 6644 19224
rect 4663 19193 4675 19196
rect 4617 19187 4675 19193
rect 6638 19184 6644 19196
rect 6696 19184 6702 19236
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2866 19156 2872 19168
rect 2547 19128 2872 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2866 19116 2872 19128
rect 2924 19116 2930 19168
rect 4154 19116 4160 19168
rect 4212 19116 4218 19168
rect 4246 19116 4252 19168
rect 4304 19156 4310 19168
rect 4982 19156 4988 19168
rect 4304 19128 4988 19156
rect 4304 19116 4310 19128
rect 4982 19116 4988 19128
rect 5040 19116 5046 19168
rect 7208 19156 7236 19255
rect 7282 19252 7288 19304
rect 7340 19292 7346 19304
rect 8220 19292 8248 19400
rect 9398 19388 9404 19440
rect 9456 19428 9462 19440
rect 16945 19431 17003 19437
rect 9456 19400 9536 19428
rect 9456 19388 9462 19400
rect 8294 19320 8300 19372
rect 8352 19360 8358 19372
rect 9508 19369 9536 19400
rect 16945 19397 16957 19431
rect 16991 19397 17003 19431
rect 16945 19391 17003 19397
rect 9309 19363 9367 19369
rect 9309 19360 9321 19363
rect 8352 19332 9321 19360
rect 8352 19320 8358 19332
rect 9309 19329 9321 19332
rect 9355 19329 9367 19363
rect 9309 19323 9367 19329
rect 9493 19363 9551 19369
rect 9493 19329 9505 19363
rect 9539 19329 9551 19363
rect 9493 19323 9551 19329
rect 14369 19363 14427 19369
rect 14369 19329 14381 19363
rect 14415 19360 14427 19363
rect 14734 19360 14740 19372
rect 14415 19332 14740 19360
rect 14415 19329 14427 19332
rect 14369 19323 14427 19329
rect 14734 19320 14740 19332
rect 14792 19320 14798 19372
rect 15470 19360 15476 19372
rect 15431 19332 15476 19360
rect 15470 19320 15476 19332
rect 15528 19320 15534 19372
rect 7340 19264 8248 19292
rect 7340 19252 7346 19264
rect 8662 19252 8668 19304
rect 8720 19292 8726 19304
rect 10042 19292 10048 19304
rect 8720 19264 10048 19292
rect 8720 19252 8726 19264
rect 10042 19252 10048 19264
rect 10100 19252 10106 19304
rect 10413 19295 10471 19301
rect 10413 19261 10425 19295
rect 10459 19292 10471 19295
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 10459 19264 12449 19292
rect 10459 19261 10471 19264
rect 10413 19255 10471 19261
rect 12437 19261 12449 19264
rect 12483 19292 12495 19295
rect 13170 19292 13176 19304
rect 12483 19264 13176 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 13170 19252 13176 19264
rect 13228 19252 13234 19304
rect 14090 19292 14096 19304
rect 14051 19264 14096 19292
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 15841 19295 15899 19301
rect 15841 19292 15853 19295
rect 14844 19264 15853 19292
rect 7460 19227 7518 19233
rect 7460 19193 7472 19227
rect 7506 19224 7518 19227
rect 10680 19227 10738 19233
rect 7506 19196 10272 19224
rect 7506 19193 7518 19196
rect 7460 19187 7518 19193
rect 7650 19156 7656 19168
rect 7208 19128 7656 19156
rect 7650 19116 7656 19128
rect 7708 19116 7714 19168
rect 8849 19159 8907 19165
rect 8849 19125 8861 19159
rect 8895 19156 8907 19159
rect 8938 19156 8944 19168
rect 8895 19128 8944 19156
rect 8895 19125 8907 19128
rect 8849 19119 8907 19125
rect 8938 19116 8944 19128
rect 8996 19116 9002 19168
rect 9214 19156 9220 19168
rect 9175 19128 9220 19156
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 9306 19116 9312 19168
rect 9364 19156 9370 19168
rect 9861 19159 9919 19165
rect 9861 19156 9873 19159
rect 9364 19128 9873 19156
rect 9364 19116 9370 19128
rect 9861 19125 9873 19128
rect 9907 19125 9919 19159
rect 10244 19156 10272 19196
rect 10680 19193 10692 19227
rect 10726 19224 10738 19227
rect 11698 19224 11704 19236
rect 10726 19196 11704 19224
rect 10726 19193 10738 19196
rect 10680 19187 10738 19193
rect 11698 19184 11704 19196
rect 11756 19184 11762 19236
rect 12704 19227 12762 19233
rect 12704 19193 12716 19227
rect 12750 19224 12762 19227
rect 12802 19224 12808 19236
rect 12750 19196 12808 19224
rect 12750 19193 12762 19196
rect 12704 19187 12762 19193
rect 12802 19184 12808 19196
rect 12860 19184 12866 19236
rect 14550 19224 14556 19236
rect 12912 19196 14556 19224
rect 11790 19156 11796 19168
rect 10244 19128 11796 19156
rect 9861 19119 9919 19125
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 12912 19156 12940 19196
rect 14550 19184 14556 19196
rect 14608 19184 14614 19236
rect 12492 19128 12940 19156
rect 12492 19116 12498 19128
rect 13538 19116 13544 19168
rect 13596 19156 13602 19168
rect 14844 19165 14872 19264
rect 15841 19261 15853 19264
rect 15887 19261 15899 19295
rect 15841 19255 15899 19261
rect 16117 19295 16175 19301
rect 16117 19261 16129 19295
rect 16163 19292 16175 19295
rect 16574 19292 16580 19304
rect 16163 19264 16580 19292
rect 16163 19261 16175 19264
rect 16117 19255 16175 19261
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 16960 19292 16988 19391
rect 17589 19363 17647 19369
rect 17589 19329 17601 19363
rect 17635 19360 17647 19363
rect 18230 19360 18236 19372
rect 17635 19332 18236 19360
rect 17635 19329 17647 19332
rect 17589 19323 17647 19329
rect 18230 19320 18236 19332
rect 18288 19320 18294 19372
rect 18325 19363 18383 19369
rect 18325 19329 18337 19363
rect 18371 19360 18383 19363
rect 18506 19360 18512 19372
rect 18371 19332 18512 19360
rect 18371 19329 18383 19332
rect 18325 19323 18383 19329
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 18598 19320 18604 19372
rect 18656 19360 18662 19372
rect 18656 19332 19380 19360
rect 18656 19320 18662 19332
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 16960 19264 18061 19292
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 19242 19292 19248 19304
rect 19203 19264 19248 19292
rect 18049 19255 18107 19261
rect 19242 19252 19248 19264
rect 19300 19252 19306 19304
rect 19352 19292 19380 19332
rect 19981 19295 20039 19301
rect 19352 19264 19656 19292
rect 15562 19184 15568 19236
rect 15620 19224 15626 19236
rect 19334 19224 19340 19236
rect 15620 19196 19340 19224
rect 15620 19184 15626 19196
rect 19334 19184 19340 19196
rect 19392 19184 19398 19236
rect 19518 19224 19524 19236
rect 19479 19196 19524 19224
rect 19518 19184 19524 19196
rect 19576 19184 19582 19236
rect 19628 19224 19656 19264
rect 19981 19261 19993 19295
rect 20027 19292 20039 19295
rect 20070 19292 20076 19304
rect 20027 19264 20076 19292
rect 20027 19261 20039 19264
rect 19981 19255 20039 19261
rect 20070 19252 20076 19264
rect 20128 19252 20134 19304
rect 20530 19292 20536 19304
rect 20491 19264 20536 19292
rect 20530 19252 20536 19264
rect 20588 19252 20594 19304
rect 22094 19224 22100 19236
rect 19628 19196 22100 19224
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 13817 19159 13875 19165
rect 13817 19156 13829 19159
rect 13596 19128 13829 19156
rect 13596 19116 13602 19128
rect 13817 19125 13829 19128
rect 13863 19125 13875 19159
rect 13817 19119 13875 19125
rect 14829 19159 14887 19165
rect 14829 19125 14841 19159
rect 14875 19125 14887 19159
rect 15194 19156 15200 19168
rect 15155 19128 15200 19156
rect 14829 19119 14887 19125
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 15289 19159 15347 19165
rect 15289 19125 15301 19159
rect 15335 19156 15347 19159
rect 15930 19156 15936 19168
rect 15335 19128 15936 19156
rect 15335 19125 15347 19128
rect 15289 19119 15347 19125
rect 15930 19116 15936 19128
rect 15988 19116 15994 19168
rect 17310 19156 17316 19168
rect 17271 19128 17316 19156
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 17402 19116 17408 19168
rect 17460 19156 17466 19168
rect 17460 19128 17505 19156
rect 17460 19116 17466 19128
rect 17586 19116 17592 19168
rect 17644 19156 17650 19168
rect 18785 19159 18843 19165
rect 18785 19156 18797 19159
rect 17644 19128 18797 19156
rect 17644 19116 17650 19128
rect 18785 19125 18797 19128
rect 18831 19125 18843 19159
rect 18785 19119 18843 19125
rect 19150 19116 19156 19168
rect 19208 19156 19214 19168
rect 20165 19159 20223 19165
rect 20165 19156 20177 19159
rect 19208 19128 20177 19156
rect 19208 19116 19214 19128
rect 20165 19125 20177 19128
rect 20211 19125 20223 19159
rect 20714 19156 20720 19168
rect 20675 19128 20720 19156
rect 20165 19119 20223 19125
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 2685 18955 2743 18961
rect 2685 18921 2697 18955
rect 2731 18952 2743 18955
rect 2774 18952 2780 18964
rect 2731 18924 2780 18952
rect 2731 18921 2743 18924
rect 2685 18915 2743 18921
rect 2774 18912 2780 18924
rect 2832 18912 2838 18964
rect 3786 18952 3792 18964
rect 2884 18924 3792 18952
rect 2884 18884 2912 18924
rect 3786 18912 3792 18924
rect 3844 18912 3850 18964
rect 4246 18952 4252 18964
rect 4207 18924 4252 18952
rect 4246 18912 4252 18924
rect 4304 18912 4310 18964
rect 7377 18955 7435 18961
rect 7377 18921 7389 18955
rect 7423 18921 7435 18955
rect 7377 18915 7435 18921
rect 7653 18955 7711 18961
rect 7653 18921 7665 18955
rect 7699 18952 7711 18955
rect 8754 18952 8760 18964
rect 7699 18924 8760 18952
rect 7699 18921 7711 18924
rect 7653 18915 7711 18921
rect 1780 18856 2912 18884
rect 1780 18825 1808 18856
rect 5902 18844 5908 18896
rect 5960 18884 5966 18896
rect 6549 18887 6607 18893
rect 6549 18884 6561 18887
rect 5960 18856 6561 18884
rect 5960 18844 5966 18856
rect 6549 18853 6561 18856
rect 6595 18853 6607 18887
rect 7392 18884 7420 18915
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 9125 18955 9183 18961
rect 9125 18921 9137 18955
rect 9171 18952 9183 18955
rect 9398 18952 9404 18964
rect 9171 18924 9404 18952
rect 9171 18921 9183 18924
rect 9125 18915 9183 18921
rect 9398 18912 9404 18924
rect 9456 18912 9462 18964
rect 12161 18955 12219 18961
rect 12161 18921 12173 18955
rect 12207 18952 12219 18955
rect 13354 18952 13360 18964
rect 12207 18924 13360 18952
rect 12207 18921 12219 18924
rect 12161 18915 12219 18921
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 15286 18912 15292 18964
rect 15344 18952 15350 18964
rect 16853 18955 16911 18961
rect 15344 18924 16804 18952
rect 15344 18912 15350 18924
rect 12529 18887 12587 18893
rect 7392 18856 10732 18884
rect 6549 18847 6607 18853
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18785 1823 18819
rect 2498 18816 2504 18828
rect 2459 18788 2504 18816
rect 1765 18779 1823 18785
rect 2498 18776 2504 18788
rect 2556 18776 2562 18828
rect 3053 18819 3111 18825
rect 3053 18785 3065 18819
rect 3099 18785 3111 18819
rect 3053 18779 3111 18785
rect 3068 18748 3096 18779
rect 3602 18776 3608 18828
rect 3660 18816 3666 18828
rect 4065 18819 4123 18825
rect 4065 18816 4077 18819
rect 3660 18788 4077 18816
rect 3660 18776 3666 18788
rect 4065 18785 4077 18788
rect 4111 18785 4123 18819
rect 4065 18779 4123 18785
rect 4890 18776 4896 18828
rect 4948 18816 4954 18828
rect 5445 18819 5503 18825
rect 5445 18816 5457 18819
rect 4948 18788 5457 18816
rect 4948 18776 4954 18788
rect 5445 18785 5457 18788
rect 5491 18785 5503 18819
rect 6270 18816 6276 18828
rect 6231 18788 6276 18816
rect 5445 18779 5503 18785
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 7193 18819 7251 18825
rect 7193 18785 7205 18819
rect 7239 18816 7251 18819
rect 7653 18819 7711 18825
rect 7653 18816 7665 18819
rect 7239 18788 7665 18816
rect 7239 18785 7251 18788
rect 7193 18779 7251 18785
rect 7653 18785 7665 18788
rect 7699 18785 7711 18819
rect 7653 18779 7711 18785
rect 8012 18819 8070 18825
rect 8012 18785 8024 18819
rect 8058 18816 8070 18819
rect 8846 18816 8852 18828
rect 8058 18788 8852 18816
rect 8058 18785 8070 18788
rect 8012 18779 8070 18785
rect 8846 18776 8852 18788
rect 8904 18776 8910 18828
rect 9398 18776 9404 18828
rect 9456 18816 9462 18828
rect 9933 18819 9991 18825
rect 9933 18816 9945 18819
rect 9456 18788 9945 18816
rect 9456 18776 9462 18788
rect 9933 18785 9945 18788
rect 9979 18785 9991 18819
rect 9933 18779 9991 18785
rect 3878 18748 3884 18760
rect 3068 18720 3884 18748
rect 3878 18708 3884 18720
rect 3936 18708 3942 18760
rect 3970 18708 3976 18760
rect 4028 18748 4034 18760
rect 7558 18748 7564 18760
rect 4028 18720 7564 18748
rect 4028 18708 4034 18720
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 7745 18751 7803 18757
rect 7745 18717 7757 18751
rect 7791 18717 7803 18751
rect 9674 18748 9680 18760
rect 9635 18720 9680 18748
rect 7745 18711 7803 18717
rect 1949 18683 2007 18689
rect 1949 18649 1961 18683
rect 1995 18680 2007 18683
rect 2958 18680 2964 18692
rect 1995 18652 2964 18680
rect 1995 18649 2007 18652
rect 1949 18643 2007 18649
rect 2958 18640 2964 18652
rect 3016 18640 3022 18692
rect 3234 18680 3240 18692
rect 3195 18652 3240 18680
rect 3234 18640 3240 18652
rect 3292 18640 3298 18692
rect 3694 18640 3700 18692
rect 3752 18680 3758 18692
rect 5074 18680 5080 18692
rect 3752 18652 5080 18680
rect 3752 18640 3758 18652
rect 5074 18640 5080 18652
rect 5132 18640 5138 18692
rect 7650 18640 7656 18692
rect 7708 18680 7714 18692
rect 7760 18680 7788 18711
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 7708 18652 7788 18680
rect 10704 18680 10732 18856
rect 12529 18853 12541 18887
rect 12575 18884 12587 18887
rect 13078 18884 13084 18896
rect 12575 18856 13084 18884
rect 12575 18853 12587 18856
rect 12529 18847 12587 18853
rect 13078 18844 13084 18856
rect 13136 18844 13142 18896
rect 13440 18887 13498 18893
rect 13440 18853 13452 18887
rect 13486 18884 13498 18887
rect 13538 18884 13544 18896
rect 13486 18856 13544 18884
rect 13486 18853 13498 18856
rect 13440 18847 13498 18853
rect 13538 18844 13544 18856
rect 13596 18844 13602 18896
rect 15470 18844 15476 18896
rect 15528 18884 15534 18896
rect 15718 18887 15776 18893
rect 15718 18884 15730 18887
rect 15528 18856 15730 18884
rect 15528 18844 15534 18856
rect 15718 18853 15730 18856
rect 15764 18853 15776 18887
rect 15718 18847 15776 18853
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11425 18819 11483 18825
rect 11425 18816 11437 18819
rect 11112 18788 11437 18816
rect 11112 18776 11118 18788
rect 11425 18785 11437 18788
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 11701 18819 11759 18825
rect 11701 18785 11713 18819
rect 11747 18816 11759 18819
rect 16022 18816 16028 18828
rect 11747 18788 16028 18816
rect 11747 18785 11759 18788
rect 11701 18779 11759 18785
rect 16022 18776 16028 18788
rect 16080 18776 16086 18828
rect 16776 18816 16804 18924
rect 16853 18921 16865 18955
rect 16899 18921 16911 18955
rect 16853 18915 16911 18921
rect 16868 18884 16896 18915
rect 18230 18912 18236 18964
rect 18288 18952 18294 18964
rect 18509 18955 18567 18961
rect 18509 18952 18521 18955
rect 18288 18924 18521 18952
rect 18288 18912 18294 18924
rect 18509 18921 18521 18924
rect 18555 18921 18567 18955
rect 18509 18915 18567 18921
rect 17374 18887 17432 18893
rect 17374 18884 17386 18887
rect 16868 18856 17386 18884
rect 17374 18853 17386 18856
rect 17420 18884 17432 18887
rect 17494 18884 17500 18896
rect 17420 18856 17500 18884
rect 17420 18853 17432 18856
rect 17374 18847 17432 18853
rect 17494 18844 17500 18856
rect 17552 18844 17558 18896
rect 18524 18884 18552 18915
rect 19030 18887 19088 18893
rect 19030 18884 19042 18887
rect 18524 18856 19042 18884
rect 19030 18853 19042 18856
rect 19076 18853 19088 18887
rect 19030 18847 19088 18853
rect 17129 18819 17187 18825
rect 17129 18816 17141 18819
rect 16776 18788 17141 18816
rect 17129 18785 17141 18788
rect 17175 18816 17187 18819
rect 18785 18819 18843 18825
rect 18785 18816 18797 18819
rect 17175 18788 18797 18816
rect 17175 18785 17187 18788
rect 17129 18779 17187 18785
rect 18785 18785 18797 18788
rect 18831 18785 18843 18819
rect 18785 18779 18843 18785
rect 12618 18748 12624 18760
rect 12579 18720 12624 18748
rect 12618 18708 12624 18720
rect 12676 18708 12682 18760
rect 12802 18748 12808 18760
rect 12763 18720 12808 18748
rect 12802 18708 12808 18720
rect 12860 18708 12866 18760
rect 13170 18748 13176 18760
rect 13131 18720 13176 18748
rect 13170 18708 13176 18720
rect 13228 18708 13234 18760
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 15473 18751 15531 18757
rect 15473 18748 15485 18751
rect 15344 18720 15485 18748
rect 15344 18708 15350 18720
rect 15473 18717 15485 18720
rect 15519 18717 15531 18751
rect 15473 18711 15531 18717
rect 11057 18683 11115 18689
rect 10704 18652 10916 18680
rect 7708 18640 7714 18652
rect 5629 18615 5687 18621
rect 5629 18581 5641 18615
rect 5675 18612 5687 18615
rect 10778 18612 10784 18624
rect 5675 18584 10784 18612
rect 5675 18581 5687 18584
rect 5629 18575 5687 18581
rect 10778 18572 10784 18584
rect 10836 18572 10842 18624
rect 10888 18612 10916 18652
rect 11057 18649 11069 18683
rect 11103 18680 11115 18683
rect 12820 18680 12848 18708
rect 11103 18652 12848 18680
rect 11103 18649 11115 18652
rect 11057 18643 11115 18649
rect 14274 18640 14280 18692
rect 14332 18680 14338 18692
rect 14332 18652 14688 18680
rect 14332 18640 14338 18652
rect 12434 18612 12440 18624
rect 10888 18584 12440 18612
rect 12434 18572 12440 18584
rect 12492 18572 12498 18624
rect 12526 18572 12532 18624
rect 12584 18612 12590 18624
rect 13906 18612 13912 18624
rect 12584 18584 13912 18612
rect 12584 18572 12590 18584
rect 13906 18572 13912 18584
rect 13964 18572 13970 18624
rect 14550 18612 14556 18624
rect 14511 18584 14556 18612
rect 14550 18572 14556 18584
rect 14608 18572 14614 18624
rect 14660 18612 14688 18652
rect 19426 18612 19432 18624
rect 14660 18584 19432 18612
rect 19426 18572 19432 18584
rect 19484 18572 19490 18624
rect 20162 18612 20168 18624
rect 20123 18584 20168 18612
rect 20162 18572 20168 18584
rect 20220 18572 20226 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 2501 18411 2559 18417
rect 2501 18377 2513 18411
rect 2547 18408 2559 18411
rect 3050 18408 3056 18420
rect 2547 18380 3056 18408
rect 2547 18377 2559 18380
rect 2501 18371 2559 18377
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 3970 18408 3976 18420
rect 3436 18380 3976 18408
rect 3436 18340 3464 18380
rect 3970 18368 3976 18380
rect 4028 18368 4034 18420
rect 4154 18368 4160 18420
rect 4212 18408 4218 18420
rect 8205 18411 8263 18417
rect 4212 18380 7420 18408
rect 4212 18368 4218 18380
rect 1780 18312 3464 18340
rect 1780 18213 1808 18312
rect 3510 18300 3516 18352
rect 3568 18340 3574 18352
rect 6730 18340 6736 18352
rect 3568 18312 6736 18340
rect 3568 18300 3574 18312
rect 6730 18300 6736 18312
rect 6788 18300 6794 18352
rect 2498 18232 2504 18284
rect 2556 18272 2562 18284
rect 3053 18275 3111 18281
rect 3053 18272 3065 18275
rect 2556 18244 3065 18272
rect 2556 18232 2562 18244
rect 3053 18241 3065 18244
rect 3099 18241 3111 18275
rect 3053 18235 3111 18241
rect 3786 18232 3792 18284
rect 3844 18272 3850 18284
rect 4890 18272 4896 18284
rect 3844 18244 4752 18272
rect 4851 18244 4896 18272
rect 3844 18232 3850 18244
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18173 1823 18207
rect 1765 18167 1823 18173
rect 2317 18207 2375 18213
rect 2317 18173 2329 18207
rect 2363 18173 2375 18207
rect 2317 18167 2375 18173
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18204 2927 18207
rect 3510 18204 3516 18216
rect 2915 18176 3516 18204
rect 2915 18173 2927 18176
rect 2869 18167 2927 18173
rect 2332 18136 2360 18167
rect 3510 18164 3516 18176
rect 3568 18164 3574 18216
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 4617 18207 4675 18213
rect 4617 18204 4629 18207
rect 4212 18176 4629 18204
rect 4212 18164 4218 18176
rect 4617 18173 4629 18176
rect 4663 18173 4675 18207
rect 4724 18204 4752 18244
rect 4890 18232 4896 18244
rect 4948 18232 4954 18284
rect 5626 18232 5632 18284
rect 5684 18272 5690 18284
rect 6362 18272 6368 18284
rect 5684 18244 6368 18272
rect 5684 18232 5690 18244
rect 6362 18232 6368 18244
rect 6420 18232 6426 18284
rect 6454 18232 6460 18284
rect 6512 18272 6518 18284
rect 7282 18272 7288 18284
rect 6512 18244 7288 18272
rect 6512 18232 6518 18244
rect 7282 18232 7288 18244
rect 7340 18232 7346 18284
rect 4798 18204 4804 18216
rect 4724 18176 4804 18204
rect 4617 18167 4675 18173
rect 4798 18164 4804 18176
rect 4856 18164 4862 18216
rect 6822 18164 6828 18216
rect 6880 18204 6886 18216
rect 6880 18176 7052 18204
rect 6880 18164 6886 18176
rect 6086 18136 6092 18148
rect 2332 18108 6092 18136
rect 6086 18096 6092 18108
rect 6144 18096 6150 18148
rect 6178 18096 6184 18148
rect 6236 18136 6242 18148
rect 6914 18136 6920 18148
rect 6236 18108 6920 18136
rect 6236 18096 6242 18108
rect 6914 18096 6920 18108
rect 6972 18096 6978 18148
rect 7024 18136 7052 18176
rect 7392 18136 7420 18380
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 9214 18408 9220 18420
rect 8251 18380 9220 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 9214 18368 9220 18380
rect 9272 18368 9278 18420
rect 12805 18411 12863 18417
rect 12805 18408 12817 18411
rect 9508 18380 12817 18408
rect 7466 18232 7472 18284
rect 7524 18272 7530 18284
rect 7561 18275 7619 18281
rect 7561 18272 7573 18275
rect 7524 18244 7573 18272
rect 7524 18232 7530 18244
rect 7561 18241 7573 18244
rect 7607 18272 7619 18275
rect 7742 18272 7748 18284
rect 7607 18244 7748 18272
rect 7607 18241 7619 18244
rect 7561 18235 7619 18241
rect 7742 18232 7748 18244
rect 7800 18232 7806 18284
rect 8846 18232 8852 18284
rect 8904 18272 8910 18284
rect 9508 18281 9536 18380
rect 12805 18377 12817 18380
rect 12851 18377 12863 18411
rect 12805 18371 12863 18377
rect 12897 18411 12955 18417
rect 12897 18377 12909 18411
rect 12943 18408 12955 18411
rect 13262 18408 13268 18420
rect 12943 18380 13268 18408
rect 12943 18377 12955 18380
rect 12897 18371 12955 18377
rect 13262 18368 13268 18380
rect 13320 18368 13326 18420
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 15657 18411 15715 18417
rect 15657 18408 15669 18411
rect 15528 18380 15669 18408
rect 15528 18368 15534 18380
rect 15657 18377 15669 18380
rect 15703 18377 15715 18411
rect 15930 18408 15936 18420
rect 15891 18380 15936 18408
rect 15657 18371 15715 18377
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 16945 18411 17003 18417
rect 16945 18377 16957 18411
rect 16991 18408 17003 18411
rect 17310 18408 17316 18420
rect 16991 18380 17316 18408
rect 16991 18377 17003 18380
rect 16945 18371 17003 18377
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 18233 18411 18291 18417
rect 18233 18377 18245 18411
rect 18279 18408 18291 18411
rect 18874 18408 18880 18420
rect 18279 18380 18880 18408
rect 18279 18377 18291 18380
rect 18233 18371 18291 18377
rect 18874 18368 18880 18380
rect 18932 18368 18938 18420
rect 20806 18408 20812 18420
rect 20767 18380 20812 18408
rect 20806 18368 20812 18380
rect 20864 18368 20870 18420
rect 11517 18343 11575 18349
rect 11517 18309 11529 18343
rect 11563 18340 11575 18343
rect 11698 18340 11704 18352
rect 11563 18312 11704 18340
rect 11563 18309 11575 18312
rect 11517 18303 11575 18309
rect 11698 18300 11704 18312
rect 11756 18300 11762 18352
rect 12250 18300 12256 18352
rect 12308 18340 12314 18352
rect 13170 18340 13176 18352
rect 12308 18312 13176 18340
rect 12308 18300 12314 18312
rect 13170 18300 13176 18312
rect 13228 18340 13234 18352
rect 15749 18343 15807 18349
rect 13228 18312 14320 18340
rect 13228 18300 13234 18312
rect 9493 18275 9551 18281
rect 8904 18244 8949 18272
rect 8904 18232 8910 18244
rect 9493 18241 9505 18275
rect 9539 18241 9551 18275
rect 9493 18235 9551 18241
rect 9600 18244 10272 18272
rect 8570 18204 8576 18216
rect 8531 18176 8576 18204
rect 8570 18164 8576 18176
rect 8628 18164 8634 18216
rect 8938 18164 8944 18216
rect 8996 18204 9002 18216
rect 9217 18207 9275 18213
rect 9217 18204 9229 18207
rect 8996 18176 9229 18204
rect 8996 18164 9002 18176
rect 9217 18173 9229 18176
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 7469 18139 7527 18145
rect 7469 18136 7481 18139
rect 7024 18108 7144 18136
rect 7392 18108 7481 18136
rect 7006 18068 7012 18080
rect 6967 18040 7012 18068
rect 7006 18028 7012 18040
rect 7064 18028 7070 18080
rect 7116 18068 7144 18108
rect 7469 18105 7481 18108
rect 7515 18105 7527 18139
rect 8662 18136 8668 18148
rect 8623 18108 8668 18136
rect 7469 18099 7527 18105
rect 7377 18071 7435 18077
rect 7377 18068 7389 18071
rect 7116 18040 7389 18068
rect 7377 18037 7389 18040
rect 7423 18037 7435 18071
rect 7484 18068 7512 18099
rect 8662 18096 8668 18108
rect 8720 18096 8726 18148
rect 9600 18136 9628 18244
rect 10244 18216 10272 18244
rect 11238 18232 11244 18284
rect 11296 18272 11302 18284
rect 11974 18272 11980 18284
rect 11296 18244 11980 18272
rect 11296 18232 11302 18244
rect 11974 18232 11980 18244
rect 12032 18232 12038 18284
rect 12802 18232 12808 18284
rect 12860 18272 12866 18284
rect 14292 18281 14320 18312
rect 15749 18309 15761 18343
rect 15795 18340 15807 18343
rect 16758 18340 16764 18352
rect 15795 18312 16764 18340
rect 15795 18309 15807 18312
rect 15749 18303 15807 18309
rect 16758 18300 16764 18312
rect 16816 18300 16822 18352
rect 18601 18343 18659 18349
rect 18601 18309 18613 18343
rect 18647 18340 18659 18343
rect 19334 18340 19340 18352
rect 18647 18312 19340 18340
rect 18647 18309 18659 18312
rect 18601 18303 18659 18309
rect 19334 18300 19340 18312
rect 19392 18300 19398 18352
rect 13449 18275 13507 18281
rect 13449 18272 13461 18275
rect 12860 18244 13461 18272
rect 12860 18232 12866 18244
rect 13449 18241 13461 18244
rect 13495 18241 13507 18275
rect 13449 18235 13507 18241
rect 14277 18275 14335 18281
rect 14277 18241 14289 18275
rect 14323 18241 14335 18275
rect 14277 18235 14335 18241
rect 16485 18275 16543 18281
rect 16485 18241 16497 18275
rect 16531 18241 16543 18275
rect 17494 18272 17500 18284
rect 17455 18244 17500 18272
rect 16485 18235 16543 18241
rect 9674 18164 9680 18216
rect 9732 18204 9738 18216
rect 10137 18207 10195 18213
rect 10137 18204 10149 18207
rect 9732 18176 10149 18204
rect 9732 18164 9738 18176
rect 10137 18173 10149 18176
rect 10183 18173 10195 18207
rect 10137 18167 10195 18173
rect 10226 18164 10232 18216
rect 10284 18164 10290 18216
rect 10778 18164 10784 18216
rect 10836 18204 10842 18216
rect 12526 18204 12532 18216
rect 10836 18176 12532 18204
rect 10836 18164 10842 18176
rect 12526 18164 12532 18176
rect 12584 18164 12590 18216
rect 13357 18207 13415 18213
rect 13357 18173 13369 18207
rect 13403 18204 13415 18207
rect 13538 18204 13544 18216
rect 13403 18176 13544 18204
rect 13403 18173 13415 18176
rect 13357 18167 13415 18173
rect 13538 18164 13544 18176
rect 13596 18164 13602 18216
rect 16393 18207 16451 18213
rect 16393 18204 16405 18207
rect 13924 18176 16405 18204
rect 9140 18108 9628 18136
rect 9140 18068 9168 18108
rect 9766 18096 9772 18148
rect 9824 18136 9830 18148
rect 10382 18139 10440 18145
rect 10382 18136 10394 18139
rect 9824 18108 10394 18136
rect 9824 18096 9830 18108
rect 10382 18105 10394 18108
rect 10428 18105 10440 18139
rect 10382 18099 10440 18105
rect 10594 18096 10600 18148
rect 10652 18136 10658 18148
rect 12066 18136 12072 18148
rect 10652 18108 12072 18136
rect 10652 18096 10658 18108
rect 12066 18096 12072 18108
rect 12124 18096 12130 18148
rect 12437 18139 12495 18145
rect 12437 18105 12449 18139
rect 12483 18136 12495 18139
rect 13265 18139 13323 18145
rect 13265 18136 13277 18139
rect 12483 18108 13277 18136
rect 12483 18105 12495 18108
rect 12437 18099 12495 18105
rect 13265 18105 13277 18108
rect 13311 18105 13323 18139
rect 13265 18099 13323 18105
rect 13446 18096 13452 18148
rect 13504 18136 13510 18148
rect 13924 18136 13952 18176
rect 16393 18173 16405 18176
rect 16439 18173 16451 18207
rect 16393 18167 16451 18173
rect 14550 18145 14556 18148
rect 14544 18136 14556 18145
rect 13504 18108 13952 18136
rect 14511 18108 14556 18136
rect 13504 18096 13510 18108
rect 14544 18099 14556 18108
rect 14608 18136 14614 18148
rect 15838 18136 15844 18148
rect 14608 18108 15844 18136
rect 14550 18096 14556 18099
rect 14608 18096 14614 18108
rect 15838 18096 15844 18108
rect 15896 18136 15902 18148
rect 16500 18136 16528 18235
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 19150 18232 19156 18284
rect 19208 18272 19214 18284
rect 19245 18275 19303 18281
rect 19245 18272 19257 18275
rect 19208 18244 19257 18272
rect 19208 18232 19214 18244
rect 19245 18241 19257 18244
rect 19291 18272 19303 18275
rect 20162 18272 20168 18284
rect 19291 18244 20168 18272
rect 19291 18241 19303 18244
rect 19245 18235 19303 18241
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 17313 18207 17371 18213
rect 17313 18173 17325 18207
rect 17359 18204 17371 18207
rect 17586 18204 17592 18216
rect 17359 18176 17592 18204
rect 17359 18173 17371 18176
rect 17313 18167 17371 18173
rect 17586 18164 17592 18176
rect 17644 18164 17650 18216
rect 18049 18207 18107 18213
rect 18049 18173 18061 18207
rect 18095 18204 18107 18207
rect 19518 18204 19524 18216
rect 18095 18176 19524 18204
rect 18095 18173 18107 18176
rect 18049 18167 18107 18173
rect 19518 18164 19524 18176
rect 19576 18164 19582 18216
rect 20254 18164 20260 18216
rect 20312 18204 20318 18216
rect 20625 18207 20683 18213
rect 20625 18204 20637 18207
rect 20312 18176 20637 18204
rect 20312 18164 20318 18176
rect 20625 18173 20637 18176
rect 20671 18173 20683 18207
rect 20625 18167 20683 18173
rect 19061 18139 19119 18145
rect 19061 18136 19073 18139
rect 15896 18108 16528 18136
rect 16592 18108 19073 18136
rect 15896 18096 15902 18108
rect 7484 18040 9168 18068
rect 7377 18031 7435 18037
rect 9214 18028 9220 18080
rect 9272 18068 9278 18080
rect 10870 18068 10876 18080
rect 9272 18040 10876 18068
rect 9272 18028 9278 18040
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 11790 18068 11796 18080
rect 11751 18040 11796 18068
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 12805 18071 12863 18077
rect 12805 18037 12817 18071
rect 12851 18068 12863 18071
rect 15749 18071 15807 18077
rect 15749 18068 15761 18071
rect 12851 18040 15761 18068
rect 12851 18037 12863 18040
rect 12805 18031 12863 18037
rect 15749 18037 15761 18040
rect 15795 18037 15807 18071
rect 16298 18068 16304 18080
rect 16259 18040 16304 18068
rect 15749 18031 15807 18037
rect 16298 18028 16304 18040
rect 16356 18028 16362 18080
rect 16482 18028 16488 18080
rect 16540 18068 16546 18080
rect 16592 18068 16620 18108
rect 19061 18105 19073 18108
rect 19107 18105 19119 18139
rect 19061 18099 19119 18105
rect 16540 18040 16620 18068
rect 17405 18071 17463 18077
rect 16540 18028 16546 18040
rect 17405 18037 17417 18071
rect 17451 18068 17463 18071
rect 17586 18068 17592 18080
rect 17451 18040 17592 18068
rect 17451 18037 17463 18040
rect 17405 18031 17463 18037
rect 17586 18028 17592 18040
rect 17644 18028 17650 18080
rect 18874 18028 18880 18080
rect 18932 18068 18938 18080
rect 18969 18071 19027 18077
rect 18969 18068 18981 18071
rect 18932 18040 18981 18068
rect 18932 18028 18938 18040
rect 18969 18037 18981 18040
rect 19015 18037 19027 18071
rect 18969 18031 19027 18037
rect 19426 18028 19432 18080
rect 19484 18068 19490 18080
rect 19613 18071 19671 18077
rect 19613 18068 19625 18071
rect 19484 18040 19625 18068
rect 19484 18028 19490 18040
rect 19613 18037 19625 18040
rect 19659 18037 19671 18071
rect 19978 18068 19984 18080
rect 19939 18040 19984 18068
rect 19613 18031 19671 18037
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 20073 18071 20131 18077
rect 20073 18037 20085 18071
rect 20119 18068 20131 18071
rect 20162 18068 20168 18080
rect 20119 18040 20168 18068
rect 20119 18037 20131 18040
rect 20073 18031 20131 18037
rect 20162 18028 20168 18040
rect 20220 18068 20226 18080
rect 20530 18068 20536 18080
rect 20220 18040 20536 18068
rect 20220 18028 20226 18040
rect 20530 18028 20536 18040
rect 20588 18028 20594 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1946 17864 1952 17876
rect 1907 17836 1952 17864
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 2498 17864 2504 17876
rect 2459 17836 2504 17864
rect 2498 17824 2504 17836
rect 2556 17824 2562 17876
rect 3786 17824 3792 17876
rect 3844 17864 3850 17876
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 3844 17836 4077 17864
rect 3844 17824 3850 17836
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 7009 17867 7067 17873
rect 7009 17833 7021 17867
rect 7055 17864 7067 17867
rect 7558 17864 7564 17876
rect 7055 17836 7564 17864
rect 7055 17833 7067 17836
rect 7009 17827 7067 17833
rect 7558 17824 7564 17836
rect 7616 17824 7622 17876
rect 7650 17824 7656 17876
rect 7708 17864 7714 17876
rect 8294 17864 8300 17876
rect 7708 17836 8300 17864
rect 7708 17824 7714 17836
rect 8294 17824 8300 17836
rect 8352 17824 8358 17876
rect 9033 17867 9091 17873
rect 9033 17833 9045 17867
rect 9079 17864 9091 17867
rect 9490 17864 9496 17876
rect 9079 17836 9496 17864
rect 9079 17833 9091 17836
rect 9033 17827 9091 17833
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 11057 17867 11115 17873
rect 11057 17864 11069 17867
rect 9824 17836 11069 17864
rect 9824 17824 9830 17836
rect 11057 17833 11069 17836
rect 11103 17833 11115 17867
rect 11057 17827 11115 17833
rect 11146 17824 11152 17876
rect 11204 17864 11210 17876
rect 11333 17867 11391 17873
rect 11333 17864 11345 17867
rect 11204 17836 11345 17864
rect 11204 17824 11210 17836
rect 11333 17833 11345 17836
rect 11379 17833 11391 17867
rect 11333 17827 11391 17833
rect 11701 17867 11759 17873
rect 11701 17833 11713 17867
rect 11747 17864 11759 17867
rect 11790 17864 11796 17876
rect 11747 17836 11796 17864
rect 11747 17833 11759 17836
rect 11701 17827 11759 17833
rect 11790 17824 11796 17836
rect 11848 17824 11854 17876
rect 12802 17824 12808 17876
rect 12860 17864 12866 17876
rect 13265 17867 13323 17873
rect 13265 17864 13277 17867
rect 12860 17836 13277 17864
rect 12860 17824 12866 17836
rect 13265 17833 13277 17836
rect 13311 17864 13323 17867
rect 13311 17836 14780 17864
rect 13311 17833 13323 17836
rect 13265 17827 13323 17833
rect 5994 17796 6000 17808
rect 1780 17768 6000 17796
rect 1780 17737 1808 17768
rect 5994 17756 6000 17768
rect 6052 17756 6058 17808
rect 6822 17756 6828 17808
rect 6880 17796 6886 17808
rect 9214 17796 9220 17808
rect 6880 17768 9220 17796
rect 6880 17756 6886 17768
rect 9214 17756 9220 17768
rect 9272 17756 9278 17808
rect 9306 17756 9312 17808
rect 9364 17796 9370 17808
rect 12526 17796 12532 17808
rect 9364 17768 12532 17796
rect 9364 17756 9370 17768
rect 12526 17756 12532 17768
rect 12584 17756 12590 17808
rect 12618 17756 12624 17808
rect 12676 17796 12682 17808
rect 13357 17799 13415 17805
rect 13357 17796 13369 17799
rect 12676 17768 13369 17796
rect 12676 17756 12682 17768
rect 13357 17765 13369 17768
rect 13403 17765 13415 17799
rect 13357 17759 13415 17765
rect 14001 17799 14059 17805
rect 14001 17765 14013 17799
rect 14047 17796 14059 17799
rect 14752 17796 14780 17836
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 15289 17867 15347 17873
rect 15289 17864 15301 17867
rect 15252 17836 15301 17864
rect 15252 17824 15258 17836
rect 15289 17833 15301 17836
rect 15335 17833 15347 17867
rect 15289 17827 15347 17833
rect 15749 17867 15807 17873
rect 15749 17833 15761 17867
rect 15795 17864 15807 17867
rect 16117 17867 16175 17873
rect 16117 17864 16129 17867
rect 15795 17836 16129 17864
rect 15795 17833 15807 17836
rect 15749 17827 15807 17833
rect 16117 17833 16129 17836
rect 16163 17833 16175 17867
rect 16117 17827 16175 17833
rect 16206 17824 16212 17876
rect 16264 17864 16270 17876
rect 16485 17867 16543 17873
rect 16485 17864 16497 17867
rect 16264 17836 16497 17864
rect 16264 17824 16270 17836
rect 16485 17833 16497 17836
rect 16531 17833 16543 17867
rect 16485 17827 16543 17833
rect 16853 17867 16911 17873
rect 16853 17833 16865 17867
rect 16899 17864 16911 17867
rect 17402 17864 17408 17876
rect 16899 17836 17408 17864
rect 16899 17833 16911 17836
rect 16853 17827 16911 17833
rect 17402 17824 17408 17836
rect 17460 17824 17466 17876
rect 18598 17864 18604 17876
rect 18559 17836 18604 17864
rect 18598 17824 18604 17836
rect 18656 17824 18662 17876
rect 19610 17864 19616 17876
rect 18708 17836 19616 17864
rect 17313 17799 17371 17805
rect 17313 17796 17325 17799
rect 14047 17768 14688 17796
rect 14752 17768 17325 17796
rect 14047 17765 14059 17768
rect 14001 17759 14059 17765
rect 1765 17731 1823 17737
rect 1765 17697 1777 17731
rect 1811 17697 1823 17731
rect 2314 17728 2320 17740
rect 2275 17700 2320 17728
rect 1765 17691 1823 17697
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 2869 17731 2927 17737
rect 2869 17697 2881 17731
rect 2915 17728 2927 17731
rect 2958 17728 2964 17740
rect 2915 17700 2964 17728
rect 2915 17697 2927 17700
rect 2869 17691 2927 17697
rect 2958 17688 2964 17700
rect 3016 17688 3022 17740
rect 4246 17688 4252 17740
rect 4304 17728 4310 17740
rect 5902 17737 5908 17740
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 4304 17700 4445 17728
rect 4304 17688 4310 17700
rect 4433 17697 4445 17700
rect 4479 17697 4491 17731
rect 4433 17691 4491 17697
rect 5896 17691 5908 17737
rect 5960 17728 5966 17740
rect 7466 17728 7472 17740
rect 5960 17700 7472 17728
rect 5902 17688 5908 17691
rect 5960 17688 5966 17700
rect 7466 17688 7472 17700
rect 7524 17688 7530 17740
rect 7650 17728 7656 17740
rect 7611 17700 7656 17728
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 8481 17731 8539 17737
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 8570 17728 8576 17740
rect 8527 17700 8576 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 8570 17688 8576 17700
rect 8628 17688 8634 17740
rect 8938 17728 8944 17740
rect 8899 17700 8944 17728
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 9766 17728 9772 17740
rect 9232 17700 9772 17728
rect 2590 17620 2596 17672
rect 2648 17660 2654 17672
rect 4525 17663 4583 17669
rect 4525 17660 4537 17663
rect 2648 17632 4537 17660
rect 2648 17620 2654 17632
rect 4525 17629 4537 17632
rect 4571 17629 4583 17663
rect 4706 17660 4712 17672
rect 4667 17632 4712 17660
rect 4525 17623 4583 17629
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 4798 17620 4804 17672
rect 4856 17660 4862 17672
rect 5629 17663 5687 17669
rect 5629 17660 5641 17663
rect 4856 17632 5641 17660
rect 4856 17620 4862 17632
rect 5629 17629 5641 17632
rect 5675 17629 5687 17663
rect 5629 17623 5687 17629
rect 6822 17620 6828 17672
rect 6880 17660 6886 17672
rect 9232 17669 9260 17700
rect 9766 17688 9772 17700
rect 9824 17688 9830 17740
rect 9944 17731 10002 17737
rect 9944 17697 9956 17731
rect 9990 17728 10002 17731
rect 10502 17728 10508 17740
rect 9990 17700 10508 17728
rect 9990 17697 10002 17700
rect 9944 17691 10002 17697
rect 10502 17688 10508 17700
rect 10560 17728 10566 17740
rect 10962 17728 10968 17740
rect 10560 17700 10968 17728
rect 10560 17688 10566 17700
rect 10962 17688 10968 17700
rect 11020 17688 11026 17740
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 12345 17731 12403 17737
rect 11756 17700 11928 17728
rect 11756 17688 11762 17700
rect 11900 17672 11928 17700
rect 12345 17697 12357 17731
rect 12391 17728 12403 17731
rect 13262 17728 13268 17740
rect 12391 17700 13268 17728
rect 12391 17697 12403 17700
rect 12345 17691 12403 17697
rect 13262 17688 13268 17700
rect 13320 17688 13326 17740
rect 14366 17728 14372 17740
rect 13372 17700 14372 17728
rect 7745 17663 7803 17669
rect 7745 17660 7757 17663
rect 6880 17632 7757 17660
rect 6880 17620 6886 17632
rect 7745 17629 7757 17632
rect 7791 17629 7803 17663
rect 7745 17623 7803 17629
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17629 7895 17663
rect 7837 17623 7895 17629
rect 9217 17663 9275 17669
rect 9217 17629 9229 17663
rect 9263 17629 9275 17663
rect 9674 17660 9680 17672
rect 9635 17632 9680 17660
rect 9217 17623 9275 17629
rect 3053 17595 3111 17601
rect 3053 17561 3065 17595
rect 3099 17592 3111 17595
rect 3099 17564 5672 17592
rect 3099 17561 3111 17564
rect 3053 17555 3111 17561
rect 5644 17536 5672 17564
rect 7466 17552 7472 17604
rect 7524 17592 7530 17604
rect 7852 17592 7880 17623
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 11790 17660 11796 17672
rect 11751 17632 11796 17660
rect 11790 17620 11796 17632
rect 11848 17620 11854 17672
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 11940 17632 12033 17660
rect 11940 17620 11946 17632
rect 12066 17620 12072 17672
rect 12124 17660 12130 17672
rect 12618 17660 12624 17672
rect 12124 17632 12624 17660
rect 12124 17620 12130 17632
rect 12618 17620 12624 17632
rect 12676 17620 12682 17672
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17660 12771 17663
rect 13372 17660 13400 17700
rect 14366 17688 14372 17700
rect 14424 17688 14430 17740
rect 14461 17731 14519 17737
rect 14461 17697 14473 17731
rect 14507 17697 14519 17731
rect 14461 17691 14519 17697
rect 12759 17632 13400 17660
rect 13541 17663 13599 17669
rect 12759 17629 12771 17632
rect 12713 17623 12771 17629
rect 13541 17629 13553 17663
rect 13587 17660 13599 17663
rect 13722 17660 13728 17672
rect 13587 17632 13728 17660
rect 13587 17629 13599 17632
rect 13541 17623 13599 17629
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 8846 17592 8852 17604
rect 7524 17564 7880 17592
rect 8128 17564 8852 17592
rect 7524 17552 7530 17564
rect 5626 17484 5632 17536
rect 5684 17484 5690 17536
rect 7285 17527 7343 17533
rect 7285 17493 7297 17527
rect 7331 17524 7343 17527
rect 8128 17524 8156 17564
rect 8846 17552 8852 17564
rect 8904 17552 8910 17604
rect 14476 17592 14504 17691
rect 14660 17660 14688 17768
rect 17313 17765 17325 17768
rect 17359 17765 17371 17799
rect 18708 17796 18736 17836
rect 19610 17824 19616 17836
rect 19668 17824 19674 17876
rect 17313 17759 17371 17765
rect 17880 17768 18736 17796
rect 17880 17740 17908 17768
rect 19150 17756 19156 17808
rect 19208 17805 19214 17808
rect 19208 17799 19272 17805
rect 19208 17765 19226 17799
rect 19260 17765 19272 17799
rect 19208 17759 19272 17765
rect 19208 17756 19214 17759
rect 19886 17756 19892 17808
rect 19944 17756 19950 17808
rect 14737 17731 14795 17737
rect 14737 17697 14749 17731
rect 14783 17728 14795 17731
rect 15010 17728 15016 17740
rect 14783 17700 15016 17728
rect 14783 17697 14795 17700
rect 14737 17691 14795 17697
rect 15010 17688 15016 17700
rect 15068 17688 15074 17740
rect 15657 17731 15715 17737
rect 15657 17697 15669 17731
rect 15703 17697 15715 17731
rect 15657 17691 15715 17697
rect 16301 17731 16359 17737
rect 16301 17697 16313 17731
rect 16347 17728 16359 17731
rect 17126 17728 17132 17740
rect 16347 17700 17132 17728
rect 16347 17697 16359 17700
rect 16301 17691 16359 17697
rect 15672 17660 15700 17691
rect 17126 17688 17132 17700
rect 17184 17688 17190 17740
rect 17221 17731 17279 17737
rect 17221 17697 17233 17731
rect 17267 17728 17279 17731
rect 17678 17728 17684 17740
rect 17267 17700 17684 17728
rect 17267 17697 17279 17700
rect 17221 17691 17279 17697
rect 17678 17688 17684 17700
rect 17736 17688 17742 17740
rect 17862 17728 17868 17740
rect 17775 17700 17868 17728
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 18417 17731 18475 17737
rect 18417 17697 18429 17731
rect 18463 17728 18475 17731
rect 18690 17728 18696 17740
rect 18463 17700 18696 17728
rect 18463 17697 18475 17700
rect 18417 17691 18475 17697
rect 18690 17688 18696 17700
rect 18748 17688 18754 17740
rect 19904 17728 19932 17756
rect 18800 17700 19932 17728
rect 15838 17660 15844 17672
rect 14660 17632 15700 17660
rect 15799 17632 15844 17660
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 16117 17663 16175 17669
rect 16117 17629 16129 17663
rect 16163 17660 16175 17663
rect 17310 17660 17316 17672
rect 16163 17632 17316 17660
rect 16163 17629 16175 17632
rect 16117 17623 16175 17629
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 17494 17660 17500 17672
rect 17455 17632 17500 17660
rect 17494 17620 17500 17632
rect 17552 17620 17558 17672
rect 10612 17564 14504 17592
rect 8294 17524 8300 17536
rect 7331 17496 8156 17524
rect 8255 17496 8300 17524
rect 7331 17493 7343 17496
rect 7285 17487 7343 17493
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 8573 17527 8631 17533
rect 8573 17493 8585 17527
rect 8619 17524 8631 17527
rect 10612 17524 10640 17564
rect 14550 17552 14556 17604
rect 14608 17592 14614 17604
rect 18800 17592 18828 17700
rect 18874 17620 18880 17672
rect 18932 17660 18938 17672
rect 18969 17663 19027 17669
rect 18969 17660 18981 17663
rect 18932 17632 18981 17660
rect 18932 17620 18938 17632
rect 18969 17629 18981 17632
rect 19015 17629 19027 17663
rect 18969 17623 19027 17629
rect 14608 17564 18828 17592
rect 14608 17552 14614 17564
rect 8619 17496 10640 17524
rect 8619 17493 8631 17496
rect 8573 17487 8631 17493
rect 11790 17484 11796 17536
rect 11848 17524 11854 17536
rect 12066 17524 12072 17536
rect 11848 17496 12072 17524
rect 11848 17484 11854 17496
rect 12066 17484 12072 17496
rect 12124 17484 12130 17536
rect 12529 17527 12587 17533
rect 12529 17493 12541 17527
rect 12575 17524 12587 17527
rect 12713 17527 12771 17533
rect 12713 17524 12725 17527
rect 12575 17496 12725 17524
rect 12575 17493 12587 17496
rect 12529 17487 12587 17493
rect 12713 17493 12725 17496
rect 12759 17493 12771 17527
rect 12713 17487 12771 17493
rect 12897 17527 12955 17533
rect 12897 17493 12909 17527
rect 12943 17524 12955 17527
rect 13170 17524 13176 17536
rect 12943 17496 13176 17524
rect 12943 17493 12955 17496
rect 12897 17487 12955 17493
rect 13170 17484 13176 17496
rect 13228 17484 13234 17536
rect 13354 17484 13360 17536
rect 13412 17524 13418 17536
rect 17954 17524 17960 17536
rect 13412 17496 17960 17524
rect 13412 17484 13418 17496
rect 17954 17484 17960 17496
rect 18012 17484 18018 17536
rect 18049 17527 18107 17533
rect 18049 17493 18061 17527
rect 18095 17524 18107 17527
rect 19702 17524 19708 17536
rect 18095 17496 19708 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 19886 17484 19892 17536
rect 19944 17524 19950 17536
rect 20349 17527 20407 17533
rect 20349 17524 20361 17527
rect 19944 17496 20361 17524
rect 19944 17484 19950 17496
rect 20349 17493 20361 17496
rect 20395 17493 20407 17527
rect 20349 17487 20407 17493
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1946 17320 1952 17332
rect 1907 17292 1952 17320
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 2501 17323 2559 17329
rect 2501 17289 2513 17323
rect 2547 17320 2559 17323
rect 2774 17320 2780 17332
rect 2547 17292 2780 17320
rect 2547 17289 2559 17292
rect 2501 17283 2559 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 3605 17323 3663 17329
rect 3605 17289 3617 17323
rect 3651 17320 3663 17323
rect 4154 17320 4160 17332
rect 3651 17292 4160 17320
rect 3651 17289 3663 17292
rect 3605 17283 3663 17289
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 4525 17323 4583 17329
rect 4525 17289 4537 17323
rect 4571 17320 4583 17323
rect 4798 17320 4804 17332
rect 4571 17292 4804 17320
rect 4571 17289 4583 17292
rect 4525 17283 4583 17289
rect 4798 17280 4804 17292
rect 4856 17280 4862 17332
rect 5902 17280 5908 17332
rect 5960 17320 5966 17332
rect 5997 17323 6055 17329
rect 5997 17320 6009 17323
rect 5960 17292 6009 17320
rect 5960 17280 5966 17292
rect 5997 17289 6009 17292
rect 6043 17289 6055 17323
rect 6822 17320 6828 17332
rect 6783 17292 6828 17320
rect 5997 17283 6055 17289
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 9582 17280 9588 17332
rect 9640 17320 9646 17332
rect 11054 17320 11060 17332
rect 9640 17292 11060 17320
rect 9640 17280 9646 17292
rect 11054 17280 11060 17292
rect 11112 17280 11118 17332
rect 11241 17323 11299 17329
rect 11241 17289 11253 17323
rect 11287 17320 11299 17323
rect 11606 17320 11612 17332
rect 11287 17292 11612 17320
rect 11287 17289 11299 17292
rect 11241 17283 11299 17289
rect 11606 17280 11612 17292
rect 11664 17280 11670 17332
rect 11716 17292 12480 17320
rect 2682 17212 2688 17264
rect 2740 17252 2746 17264
rect 2740 17224 4660 17252
rect 2740 17212 2746 17224
rect 3786 17144 3792 17196
rect 3844 17184 3850 17196
rect 4065 17187 4123 17193
rect 4065 17184 4077 17187
rect 3844 17156 4077 17184
rect 3844 17144 3850 17156
rect 4065 17153 4077 17156
rect 4111 17153 4123 17187
rect 4065 17147 4123 17153
rect 4249 17187 4307 17193
rect 4249 17153 4261 17187
rect 4295 17184 4307 17187
rect 4632 17184 4660 17224
rect 5626 17212 5632 17264
rect 5684 17252 5690 17264
rect 5684 17224 8892 17252
rect 5684 17212 5690 17224
rect 4295 17156 4476 17184
rect 4632 17156 4752 17184
rect 4295 17153 4307 17156
rect 4249 17147 4307 17153
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 2317 17119 2375 17125
rect 2317 17085 2329 17119
rect 2363 17085 2375 17119
rect 2317 17079 2375 17085
rect 2332 17048 2360 17079
rect 4448 17048 4476 17156
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17116 4583 17119
rect 4617 17119 4675 17125
rect 4617 17116 4629 17119
rect 4571 17088 4629 17116
rect 4571 17085 4583 17088
rect 4525 17079 4583 17085
rect 4617 17085 4629 17088
rect 4663 17085 4675 17119
rect 4724 17116 4752 17156
rect 7006 17144 7012 17196
rect 7064 17184 7070 17196
rect 7285 17187 7343 17193
rect 7285 17184 7297 17187
rect 7064 17156 7297 17184
rect 7064 17144 7070 17156
rect 7285 17153 7297 17156
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17184 7527 17187
rect 7558 17184 7564 17196
rect 7515 17156 7564 17184
rect 7515 17153 7527 17156
rect 7469 17147 7527 17153
rect 7558 17144 7564 17156
rect 7616 17144 7622 17196
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 8389 17187 8447 17193
rect 8389 17184 8401 17187
rect 7800 17156 8401 17184
rect 7800 17144 7806 17156
rect 8389 17153 8401 17156
rect 8435 17153 8447 17187
rect 8864 17184 8892 17224
rect 9490 17212 9496 17264
rect 9548 17252 9554 17264
rect 11716 17252 11744 17292
rect 9548 17224 11744 17252
rect 9548 17212 9554 17224
rect 10318 17184 10324 17196
rect 8864 17156 8984 17184
rect 10279 17156 10324 17184
rect 8389 17147 8447 17153
rect 4724 17088 7788 17116
rect 4617 17079 4675 17085
rect 4884 17051 4942 17057
rect 4884 17048 4896 17051
rect 2332 17020 4200 17048
rect 4448 17020 4896 17048
rect 2130 16940 2136 16992
rect 2188 16980 2194 16992
rect 3694 16980 3700 16992
rect 2188 16952 3700 16980
rect 2188 16940 2194 16952
rect 3694 16940 3700 16952
rect 3752 16940 3758 16992
rect 3970 16980 3976 16992
rect 3931 16952 3976 16980
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 4172 16980 4200 17020
rect 4884 17017 4896 17020
rect 4930 17048 4942 17051
rect 5442 17048 5448 17060
rect 4930 17020 5448 17048
rect 4930 17017 4942 17020
rect 4884 17011 4942 17017
rect 5442 17008 5448 17020
rect 5500 17008 5506 17060
rect 7098 17048 7104 17060
rect 6932 17020 7104 17048
rect 6932 16980 6960 17020
rect 7098 17008 7104 17020
rect 7156 17008 7162 17060
rect 7760 17048 7788 17088
rect 8202 17076 8208 17128
rect 8260 17116 8266 17128
rect 8846 17116 8852 17128
rect 8260 17088 8305 17116
rect 8807 17088 8852 17116
rect 8260 17076 8266 17088
rect 8846 17076 8852 17088
rect 8904 17076 8910 17128
rect 8956 17116 8984 17156
rect 10318 17144 10324 17156
rect 10376 17144 10382 17196
rect 10870 17144 10876 17196
rect 10928 17184 10934 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 10928 17156 11713 17184
rect 10928 17144 10934 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 11882 17184 11888 17196
rect 11843 17156 11888 17184
rect 11701 17147 11759 17153
rect 11882 17144 11888 17156
rect 11940 17144 11946 17196
rect 12452 17184 12480 17292
rect 12912 17292 14596 17320
rect 12526 17212 12532 17264
rect 12584 17252 12590 17264
rect 12912 17252 12940 17292
rect 13909 17255 13967 17261
rect 13909 17252 13921 17255
rect 12584 17224 12940 17252
rect 13004 17224 13921 17252
rect 12584 17212 12590 17224
rect 13004 17184 13032 17224
rect 13909 17221 13921 17224
rect 13955 17221 13967 17255
rect 13909 17215 13967 17221
rect 13354 17184 13360 17196
rect 12452 17156 13032 17184
rect 13315 17156 13360 17184
rect 13354 17144 13360 17156
rect 13412 17144 13418 17196
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17184 13599 17187
rect 13814 17184 13820 17196
rect 13587 17156 13820 17184
rect 13587 17153 13599 17156
rect 13541 17147 13599 17153
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 13998 17144 14004 17196
rect 14056 17184 14062 17196
rect 14366 17184 14372 17196
rect 14056 17156 14372 17184
rect 14056 17144 14062 17156
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 14568 17193 14596 17292
rect 15378 17280 15384 17332
rect 15436 17320 15442 17332
rect 15841 17323 15899 17329
rect 15841 17320 15853 17323
rect 15436 17292 15853 17320
rect 15436 17280 15442 17292
rect 15841 17289 15853 17292
rect 15887 17289 15899 17323
rect 15841 17283 15899 17289
rect 16574 17280 16580 17332
rect 16632 17320 16638 17332
rect 17586 17320 17592 17332
rect 16632 17292 17592 17320
rect 16632 17280 16638 17292
rect 17586 17280 17592 17292
rect 17644 17320 17650 17332
rect 19061 17323 19119 17329
rect 17644 17292 19012 17320
rect 17644 17280 17650 17292
rect 15746 17212 15752 17264
rect 15804 17252 15810 17264
rect 16393 17255 16451 17261
rect 16393 17252 16405 17255
rect 15804 17224 16405 17252
rect 15804 17212 15810 17224
rect 16393 17221 16405 17224
rect 16439 17221 16451 17255
rect 16393 17215 16451 17221
rect 16500 17224 18920 17252
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17184 14611 17187
rect 15010 17184 15016 17196
rect 14599 17156 15016 17184
rect 14599 17153 14611 17156
rect 14553 17147 14611 17153
rect 15010 17144 15016 17156
rect 15068 17144 15074 17196
rect 16500 17184 16528 17224
rect 17126 17184 17132 17196
rect 15120 17156 16528 17184
rect 17087 17156 17132 17184
rect 8956 17088 14412 17116
rect 8297 17051 8355 17057
rect 8297 17048 8309 17051
rect 7760 17020 8309 17048
rect 8297 17017 8309 17020
rect 8343 17048 8355 17051
rect 8662 17048 8668 17060
rect 8343 17020 8668 17048
rect 8343 17017 8355 17020
rect 8297 17011 8355 17017
rect 8662 17008 8668 17020
rect 8720 17008 8726 17060
rect 8754 17008 8760 17060
rect 8812 17048 8818 17060
rect 9125 17051 9183 17057
rect 9125 17048 9137 17051
rect 8812 17020 9137 17048
rect 8812 17008 8818 17020
rect 9125 17017 9137 17020
rect 9171 17017 9183 17051
rect 9125 17011 9183 17017
rect 9214 17008 9220 17060
rect 9272 17048 9278 17060
rect 9272 17020 9904 17048
rect 9272 17008 9278 17020
rect 4172 16952 6960 16980
rect 7193 16983 7251 16989
rect 7193 16949 7205 16983
rect 7239 16980 7251 16983
rect 7837 16983 7895 16989
rect 7837 16980 7849 16983
rect 7239 16952 7849 16980
rect 7239 16949 7251 16952
rect 7193 16943 7251 16949
rect 7837 16949 7849 16952
rect 7883 16949 7895 16983
rect 7837 16943 7895 16949
rect 8938 16940 8944 16992
rect 8996 16980 9002 16992
rect 9490 16980 9496 16992
rect 8996 16952 9496 16980
rect 8996 16940 9002 16952
rect 9490 16940 9496 16952
rect 9548 16940 9554 16992
rect 9677 16983 9735 16989
rect 9677 16949 9689 16983
rect 9723 16980 9735 16983
rect 9766 16980 9772 16992
rect 9723 16952 9772 16980
rect 9723 16949 9735 16952
rect 9677 16943 9735 16949
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 9876 16980 9904 17020
rect 9950 17008 9956 17060
rect 10008 17048 10014 17060
rect 10045 17051 10103 17057
rect 10045 17048 10057 17051
rect 10008 17020 10057 17048
rect 10008 17008 10014 17020
rect 10045 17017 10057 17020
rect 10091 17017 10103 17051
rect 10045 17011 10103 17017
rect 10781 17051 10839 17057
rect 10781 17017 10793 17051
rect 10827 17048 10839 17051
rect 14277 17051 14335 17057
rect 14277 17048 14289 17051
rect 10827 17020 14289 17048
rect 10827 17017 10839 17020
rect 10781 17011 10839 17017
rect 14277 17017 14289 17020
rect 14323 17017 14335 17051
rect 14384 17048 14412 17088
rect 14642 17076 14648 17128
rect 14700 17116 14706 17128
rect 14921 17119 14979 17125
rect 14921 17116 14933 17119
rect 14700 17088 14933 17116
rect 14700 17076 14706 17088
rect 14921 17085 14933 17088
rect 14967 17085 14979 17119
rect 15120 17116 15148 17156
rect 17126 17144 17132 17156
rect 17184 17144 17190 17196
rect 17770 17144 17776 17196
rect 17828 17184 17834 17196
rect 18601 17187 18659 17193
rect 18601 17184 18613 17187
rect 17828 17156 18613 17184
rect 17828 17144 17834 17156
rect 18601 17153 18613 17156
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 14921 17079 14979 17085
rect 15028 17088 15148 17116
rect 15197 17119 15255 17125
rect 15028 17048 15056 17088
rect 15197 17085 15209 17119
rect 15243 17116 15255 17119
rect 15657 17119 15715 17125
rect 15657 17116 15669 17119
rect 15243 17088 15669 17116
rect 15243 17085 15255 17088
rect 15197 17079 15255 17085
rect 15657 17085 15669 17088
rect 15703 17085 15715 17119
rect 15657 17079 15715 17085
rect 16209 17119 16267 17125
rect 16209 17085 16221 17119
rect 16255 17116 16267 17119
rect 16850 17116 16856 17128
rect 16255 17088 16856 17116
rect 16255 17085 16267 17088
rect 16209 17079 16267 17085
rect 16850 17076 16856 17088
rect 16908 17076 16914 17128
rect 16945 17119 17003 17125
rect 16945 17085 16957 17119
rect 16991 17116 17003 17119
rect 16991 17088 18092 17116
rect 16991 17085 17003 17088
rect 16945 17079 17003 17085
rect 14384 17020 15056 17048
rect 14277 17011 14335 17017
rect 15102 17008 15108 17060
rect 15160 17048 15166 17060
rect 17862 17048 17868 17060
rect 15160 17020 17868 17048
rect 15160 17008 15166 17020
rect 17862 17008 17868 17020
rect 17920 17008 17926 17060
rect 10137 16983 10195 16989
rect 10137 16980 10149 16983
rect 9876 16952 10149 16980
rect 10137 16949 10149 16952
rect 10183 16980 10195 16983
rect 11514 16980 11520 16992
rect 10183 16952 11520 16980
rect 10183 16949 10195 16952
rect 10137 16943 10195 16949
rect 11514 16940 11520 16952
rect 11572 16940 11578 16992
rect 11609 16983 11667 16989
rect 11609 16949 11621 16983
rect 11655 16980 11667 16983
rect 11882 16980 11888 16992
rect 11655 16952 11888 16980
rect 11655 16949 11667 16952
rect 11609 16943 11667 16949
rect 11882 16940 11888 16952
rect 11940 16980 11946 16992
rect 12066 16980 12072 16992
rect 11940 16952 12072 16980
rect 11940 16940 11946 16952
rect 12066 16940 12072 16952
rect 12124 16940 12130 16992
rect 12894 16980 12900 16992
rect 12855 16952 12900 16980
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 13170 16940 13176 16992
rect 13228 16980 13234 16992
rect 13265 16983 13323 16989
rect 13265 16980 13277 16983
rect 13228 16952 13277 16980
rect 13228 16940 13234 16952
rect 13265 16949 13277 16952
rect 13311 16949 13323 16983
rect 13265 16943 13323 16949
rect 13538 16940 13544 16992
rect 13596 16980 13602 16992
rect 16482 16980 16488 16992
rect 13596 16952 16488 16980
rect 13596 16940 13602 16952
rect 16482 16940 16488 16952
rect 16540 16940 16546 16992
rect 18064 16989 18092 17088
rect 18417 17051 18475 17057
rect 18417 17017 18429 17051
rect 18463 17048 18475 17051
rect 18782 17048 18788 17060
rect 18463 17020 18788 17048
rect 18463 17017 18475 17020
rect 18417 17011 18475 17017
rect 18782 17008 18788 17020
rect 18840 17008 18846 17060
rect 18892 17048 18920 17224
rect 18984 17116 19012 17292
rect 19061 17289 19073 17323
rect 19107 17320 19119 17323
rect 19242 17320 19248 17332
rect 19107 17292 19248 17320
rect 19107 17289 19119 17292
rect 19061 17283 19119 17289
rect 19242 17280 19248 17292
rect 19300 17280 19306 17332
rect 19886 17280 19892 17332
rect 19944 17320 19950 17332
rect 20162 17320 20168 17332
rect 19944 17292 20168 17320
rect 19944 17280 19950 17292
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 19150 17212 19156 17264
rect 19208 17252 19214 17264
rect 20717 17255 20775 17261
rect 20717 17252 20729 17255
rect 19208 17224 20729 17252
rect 19208 17212 19214 17224
rect 20717 17221 20729 17224
rect 20763 17221 20775 17255
rect 20717 17215 20775 17221
rect 19334 17144 19340 17196
rect 19392 17144 19398 17196
rect 19705 17187 19763 17193
rect 19705 17153 19717 17187
rect 19751 17184 19763 17187
rect 19794 17184 19800 17196
rect 19751 17156 19800 17184
rect 19751 17153 19763 17156
rect 19705 17147 19763 17153
rect 19794 17144 19800 17156
rect 19852 17144 19858 17196
rect 19978 17144 19984 17196
rect 20036 17184 20042 17196
rect 20073 17187 20131 17193
rect 20073 17184 20085 17187
rect 20036 17156 20085 17184
rect 20036 17144 20042 17156
rect 20073 17153 20085 17156
rect 20119 17153 20131 17187
rect 20073 17147 20131 17153
rect 19352 17116 19380 17144
rect 19518 17116 19524 17128
rect 18984 17088 19380 17116
rect 19479 17088 19524 17116
rect 19518 17076 19524 17088
rect 19576 17076 19582 17128
rect 19610 17076 19616 17128
rect 19668 17076 19674 17128
rect 20530 17116 20536 17128
rect 20491 17088 20536 17116
rect 20530 17076 20536 17088
rect 20588 17076 20594 17128
rect 19628 17048 19656 17076
rect 18892 17020 19656 17048
rect 18049 16983 18107 16989
rect 18049 16949 18061 16983
rect 18095 16949 18107 16983
rect 18049 16943 18107 16949
rect 18509 16983 18567 16989
rect 18509 16949 18521 16983
rect 18555 16980 18567 16983
rect 19150 16980 19156 16992
rect 18555 16952 19156 16980
rect 18555 16949 18567 16952
rect 18509 16943 18567 16949
rect 19150 16940 19156 16952
rect 19208 16940 19214 16992
rect 19426 16980 19432 16992
rect 19387 16952 19432 16980
rect 19426 16940 19432 16952
rect 19484 16940 19490 16992
rect 19610 16940 19616 16992
rect 19668 16980 19674 16992
rect 20254 16980 20260 16992
rect 19668 16952 20260 16980
rect 19668 16940 19674 16952
rect 20254 16940 20260 16952
rect 20312 16940 20318 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1946 16776 1952 16788
rect 1907 16748 1952 16776
rect 1946 16736 1952 16748
rect 2004 16736 2010 16788
rect 2590 16776 2596 16788
rect 2551 16748 2596 16776
rect 2590 16736 2596 16748
rect 2648 16736 2654 16788
rect 2961 16779 3019 16785
rect 2961 16745 2973 16779
rect 3007 16776 3019 16779
rect 3142 16776 3148 16788
rect 3007 16748 3148 16776
rect 3007 16745 3019 16748
rect 2961 16739 3019 16745
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 5442 16776 5448 16788
rect 5403 16748 5448 16776
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 9125 16779 9183 16785
rect 9125 16745 9137 16779
rect 9171 16776 9183 16779
rect 10318 16776 10324 16788
rect 9171 16748 10324 16776
rect 9171 16745 9183 16748
rect 9125 16739 9183 16745
rect 10318 16736 10324 16748
rect 10376 16736 10382 16788
rect 10870 16736 10876 16788
rect 10928 16776 10934 16788
rect 13357 16779 13415 16785
rect 13357 16776 13369 16779
rect 10928 16748 13369 16776
rect 10928 16736 10934 16748
rect 13357 16745 13369 16748
rect 13403 16745 13415 16779
rect 13357 16739 13415 16745
rect 14093 16779 14151 16785
rect 14093 16745 14105 16779
rect 14139 16776 14151 16779
rect 14366 16776 14372 16788
rect 14139 16748 14372 16776
rect 14139 16745 14151 16748
rect 14093 16739 14151 16745
rect 14366 16736 14372 16748
rect 14424 16736 14430 16788
rect 15010 16736 15016 16788
rect 15068 16776 15074 16788
rect 17865 16779 17923 16785
rect 17865 16776 17877 16779
rect 15068 16748 17877 16776
rect 15068 16736 15074 16748
rect 17865 16745 17877 16748
rect 17911 16745 17923 16779
rect 17865 16739 17923 16745
rect 18046 16736 18052 16788
rect 18104 16776 18110 16788
rect 19518 16776 19524 16788
rect 18104 16748 19524 16776
rect 18104 16736 18110 16748
rect 19518 16736 19524 16748
rect 19576 16736 19582 16788
rect 19613 16779 19671 16785
rect 19613 16745 19625 16779
rect 19659 16745 19671 16779
rect 19613 16739 19671 16745
rect 4154 16668 4160 16720
rect 4212 16708 4218 16720
rect 4332 16711 4390 16717
rect 4332 16708 4344 16711
rect 4212 16680 4344 16708
rect 4212 16668 4218 16680
rect 4332 16677 4344 16680
rect 4378 16708 4390 16711
rect 4706 16708 4712 16720
rect 4378 16680 4712 16708
rect 4378 16677 4390 16680
rect 4332 16671 4390 16677
rect 4706 16668 4712 16680
rect 4764 16668 4770 16720
rect 7374 16708 7380 16720
rect 6104 16680 7380 16708
rect 1765 16643 1823 16649
rect 1765 16609 1777 16643
rect 1811 16640 1823 16643
rect 3786 16640 3792 16652
rect 1811 16612 2544 16640
rect 1811 16609 1823 16612
rect 1765 16603 1823 16609
rect 2516 16504 2544 16612
rect 2884 16612 3792 16640
rect 2884 16504 2912 16612
rect 3786 16600 3792 16612
rect 3844 16600 3850 16652
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16640 4123 16643
rect 4798 16640 4804 16652
rect 4111 16612 4804 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 6104 16649 6132 16680
rect 7374 16668 7380 16680
rect 7432 16668 7438 16720
rect 7466 16668 7472 16720
rect 7524 16708 7530 16720
rect 7990 16711 8048 16717
rect 7990 16708 8002 16711
rect 7524 16680 8002 16708
rect 7524 16668 7530 16680
rect 7990 16677 8002 16680
rect 8036 16677 8048 16711
rect 10502 16708 10508 16720
rect 7990 16671 8048 16677
rect 10060 16680 10508 16708
rect 6089 16643 6147 16649
rect 6089 16609 6101 16643
rect 6135 16609 6147 16643
rect 6089 16603 6147 16609
rect 6356 16643 6414 16649
rect 6356 16609 6368 16643
rect 6402 16640 6414 16643
rect 7558 16640 7564 16652
rect 6402 16612 7564 16640
rect 6402 16609 6414 16612
rect 6356 16603 6414 16609
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 8294 16640 8300 16652
rect 7760 16612 8300 16640
rect 3050 16572 3056 16584
rect 3011 16544 3056 16572
rect 3050 16532 3056 16544
rect 3108 16532 3114 16584
rect 3234 16572 3240 16584
rect 3195 16544 3240 16572
rect 3234 16532 3240 16544
rect 3292 16532 3298 16584
rect 7374 16532 7380 16584
rect 7432 16572 7438 16584
rect 7760 16581 7788 16612
rect 8294 16600 8300 16612
rect 8352 16640 8358 16652
rect 9674 16640 9680 16652
rect 8352 16612 9680 16640
rect 8352 16600 8358 16612
rect 9674 16600 9680 16612
rect 9732 16640 9738 16652
rect 9858 16640 9864 16652
rect 9732 16612 9864 16640
rect 9732 16600 9738 16612
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 10060 16649 10088 16680
rect 10502 16668 10508 16680
rect 10560 16668 10566 16720
rect 12250 16708 12256 16720
rect 11348 16680 12256 16708
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 9968 16612 10057 16640
rect 7745 16575 7803 16581
rect 7745 16572 7757 16575
rect 7432 16544 7757 16572
rect 7432 16532 7438 16544
rect 7745 16541 7757 16544
rect 7791 16541 7803 16575
rect 9968 16572 9996 16612
rect 10045 16609 10057 16612
rect 10091 16609 10103 16643
rect 10045 16603 10103 16609
rect 10226 16600 10232 16652
rect 10284 16640 10290 16652
rect 11348 16649 11376 16680
rect 12250 16668 12256 16680
rect 12308 16668 12314 16720
rect 12894 16668 12900 16720
rect 12952 16708 12958 16720
rect 14553 16711 14611 16717
rect 14553 16708 14565 16711
rect 12952 16680 14565 16708
rect 12952 16668 12958 16680
rect 14553 16677 14565 16680
rect 14599 16677 14611 16711
rect 14553 16671 14611 16677
rect 15657 16711 15715 16717
rect 15657 16677 15669 16711
rect 15703 16708 15715 16711
rect 16022 16708 16028 16720
rect 15703 16680 16028 16708
rect 15703 16677 15715 16680
rect 15657 16671 15715 16677
rect 16022 16668 16028 16680
rect 16080 16668 16086 16720
rect 16752 16711 16810 16717
rect 16752 16677 16764 16711
rect 16798 16708 16810 16711
rect 17770 16708 17776 16720
rect 16798 16680 17776 16708
rect 16798 16677 16810 16680
rect 16752 16671 16810 16677
rect 17770 16668 17776 16680
rect 17828 16708 17834 16720
rect 19628 16708 19656 16739
rect 17828 16680 19656 16708
rect 17828 16668 17834 16680
rect 11333 16643 11391 16649
rect 10284 16612 11284 16640
rect 10284 16600 10290 16612
rect 7745 16535 7803 16541
rect 9508 16544 9996 16572
rect 10137 16575 10195 16581
rect 2516 16476 2912 16504
rect 5258 16464 5264 16516
rect 5316 16504 5322 16516
rect 5718 16504 5724 16516
rect 5316 16476 5724 16504
rect 5316 16464 5322 16476
rect 5718 16464 5724 16476
rect 5776 16464 5782 16516
rect 7466 16504 7472 16516
rect 7427 16476 7472 16504
rect 7466 16464 7472 16476
rect 7524 16464 7530 16516
rect 5074 16396 5080 16448
rect 5132 16436 5138 16448
rect 9508 16436 9536 16544
rect 10137 16541 10149 16575
rect 10183 16541 10195 16575
rect 10318 16572 10324 16584
rect 10279 16544 10324 16572
rect 10137 16535 10195 16541
rect 9582 16464 9588 16516
rect 9640 16504 9646 16516
rect 10152 16504 10180 16535
rect 10318 16532 10324 16544
rect 10376 16532 10382 16584
rect 11256 16572 11284 16612
rect 11333 16609 11345 16643
rect 11379 16609 11391 16643
rect 11333 16603 11391 16609
rect 11600 16643 11658 16649
rect 11600 16609 11612 16643
rect 11646 16640 11658 16643
rect 11882 16640 11888 16652
rect 11646 16612 11888 16640
rect 11646 16609 11658 16612
rect 11600 16603 11658 16609
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 13449 16643 13507 16649
rect 13449 16640 13461 16643
rect 12360 16612 13461 16640
rect 11256 16544 11376 16572
rect 9640 16476 10180 16504
rect 9640 16464 9646 16476
rect 9674 16436 9680 16448
rect 5132 16408 9536 16436
rect 9635 16408 9680 16436
rect 5132 16396 5138 16408
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 11348 16436 11376 16544
rect 12360 16436 12388 16612
rect 13449 16609 13461 16612
rect 13495 16640 13507 16643
rect 13495 16612 14044 16640
rect 13495 16609 13507 16612
rect 13449 16603 13507 16609
rect 13633 16575 13691 16581
rect 13633 16541 13645 16575
rect 13679 16541 13691 16575
rect 14016 16572 14044 16612
rect 14090 16600 14096 16652
rect 14148 16640 14154 16652
rect 14461 16643 14519 16649
rect 14461 16640 14473 16643
rect 14148 16612 14473 16640
rect 14148 16600 14154 16612
rect 14461 16609 14473 16612
rect 14507 16609 14519 16643
rect 15102 16640 15108 16652
rect 14461 16603 14519 16609
rect 14568 16612 15108 16640
rect 14568 16572 14596 16612
rect 15102 16600 15108 16612
rect 15160 16600 15166 16652
rect 15286 16600 15292 16652
rect 15344 16640 15350 16652
rect 18233 16643 18291 16649
rect 18233 16640 18245 16643
rect 15344 16612 15976 16640
rect 15344 16600 15350 16612
rect 15948 16584 15976 16612
rect 16500 16612 18245 16640
rect 14016 16544 14596 16572
rect 14737 16575 14795 16581
rect 13633 16535 13691 16541
rect 14737 16541 14749 16575
rect 14783 16572 14795 16575
rect 15562 16572 15568 16584
rect 14783 16544 15568 16572
rect 14783 16541 14795 16544
rect 14737 16535 14795 16541
rect 12989 16507 13047 16513
rect 12989 16473 13001 16507
rect 13035 16504 13047 16507
rect 13354 16504 13360 16516
rect 13035 16476 13360 16504
rect 13035 16473 13047 16476
rect 12989 16467 13047 16473
rect 13354 16464 13360 16476
rect 13412 16464 13418 16516
rect 13648 16504 13676 16535
rect 15562 16532 15568 16544
rect 15620 16532 15626 16584
rect 15654 16532 15660 16584
rect 15712 16572 15718 16584
rect 15749 16575 15807 16581
rect 15749 16572 15761 16575
rect 15712 16544 15761 16572
rect 15712 16532 15718 16544
rect 15749 16541 15761 16544
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 13722 16504 13728 16516
rect 13635 16476 13728 16504
rect 12710 16436 12716 16448
rect 11348 16408 12388 16436
rect 12623 16408 12716 16436
rect 12710 16396 12716 16408
rect 12768 16436 12774 16448
rect 13648 16436 13676 16476
rect 13722 16464 13728 16476
rect 13780 16504 13786 16516
rect 15194 16504 15200 16516
rect 13780 16476 15200 16504
rect 13780 16464 13786 16476
rect 15194 16464 15200 16476
rect 15252 16504 15258 16516
rect 15856 16504 15884 16535
rect 15930 16532 15936 16584
rect 15988 16572 15994 16584
rect 16500 16581 16528 16612
rect 18233 16609 18245 16612
rect 18279 16609 18291 16643
rect 18233 16603 18291 16609
rect 18500 16643 18558 16649
rect 18500 16609 18512 16643
rect 18546 16640 18558 16643
rect 19058 16640 19064 16652
rect 18546 16612 19064 16640
rect 18546 16609 18558 16612
rect 18500 16603 18558 16609
rect 16485 16575 16543 16581
rect 16485 16572 16497 16575
rect 15988 16544 16497 16572
rect 15988 16532 15994 16544
rect 16485 16541 16497 16544
rect 16531 16541 16543 16575
rect 16485 16535 16543 16541
rect 15252 16476 15884 16504
rect 15252 16464 15258 16476
rect 15286 16436 15292 16448
rect 12768 16408 13676 16436
rect 15247 16408 15292 16436
rect 12768 16396 12774 16408
rect 15286 16396 15292 16408
rect 15344 16396 15350 16448
rect 18248 16436 18276 16603
rect 19058 16600 19064 16612
rect 19116 16600 19122 16652
rect 19242 16600 19248 16652
rect 19300 16640 19306 16652
rect 19889 16643 19947 16649
rect 19889 16640 19901 16643
rect 19300 16612 19901 16640
rect 19300 16600 19306 16612
rect 19889 16609 19901 16612
rect 19935 16609 19947 16643
rect 19889 16603 19947 16609
rect 19978 16600 19984 16652
rect 20036 16640 20042 16652
rect 20165 16643 20223 16649
rect 20165 16640 20177 16643
rect 20036 16612 20177 16640
rect 20036 16600 20042 16612
rect 20165 16609 20177 16612
rect 20211 16609 20223 16643
rect 20165 16603 20223 16609
rect 20898 16572 20904 16584
rect 20859 16544 20904 16572
rect 20898 16532 20904 16544
rect 20956 16532 20962 16584
rect 18598 16436 18604 16448
rect 18248 16408 18604 16436
rect 18598 16396 18604 16408
rect 18656 16436 18662 16448
rect 18966 16436 18972 16448
rect 18656 16408 18972 16436
rect 18656 16396 18662 16408
rect 18966 16396 18972 16408
rect 19024 16396 19030 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 3973 16235 4031 16241
rect 2608 16204 3556 16232
rect 2222 16056 2228 16108
rect 2280 16096 2286 16108
rect 2608 16105 2636 16204
rect 3528 16164 3556 16204
rect 3973 16201 3985 16235
rect 4019 16232 4031 16235
rect 4154 16232 4160 16244
rect 4019 16204 4160 16232
rect 4019 16201 4031 16204
rect 3973 16195 4031 16201
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 4246 16192 4252 16244
rect 4304 16232 4310 16244
rect 4341 16235 4399 16241
rect 4341 16232 4353 16235
rect 4304 16204 4353 16232
rect 4304 16192 4310 16204
rect 4341 16201 4353 16204
rect 4387 16201 4399 16235
rect 4798 16232 4804 16244
rect 4341 16195 4399 16201
rect 4448 16204 4804 16232
rect 4448 16164 4476 16204
rect 4798 16192 4804 16204
rect 4856 16232 4862 16244
rect 5353 16235 5411 16241
rect 5353 16232 5365 16235
rect 4856 16204 5365 16232
rect 4856 16192 4862 16204
rect 5353 16201 5365 16204
rect 5399 16201 5411 16235
rect 5353 16195 5411 16201
rect 6917 16235 6975 16241
rect 6917 16201 6929 16235
rect 6963 16232 6975 16235
rect 7650 16232 7656 16244
rect 6963 16204 7656 16232
rect 6963 16201 6975 16204
rect 6917 16195 6975 16201
rect 7650 16192 7656 16204
rect 7708 16192 7714 16244
rect 11790 16232 11796 16244
rect 10060 16204 11796 16232
rect 10060 16164 10088 16204
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 13909 16235 13967 16241
rect 13909 16232 13921 16235
rect 13872 16204 13921 16232
rect 13872 16192 13878 16204
rect 13909 16201 13921 16204
rect 13955 16201 13967 16235
rect 15562 16232 15568 16244
rect 15523 16204 15568 16232
rect 13909 16195 13967 16201
rect 3528 16136 4476 16164
rect 4724 16136 7144 16164
rect 4264 16108 4292 16136
rect 2593 16099 2651 16105
rect 2593 16096 2605 16099
rect 2280 16068 2605 16096
rect 2280 16056 2286 16068
rect 2593 16065 2605 16068
rect 2639 16065 2651 16099
rect 2593 16059 2651 16065
rect 4246 16056 4252 16108
rect 4304 16056 4310 16108
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 15997 1823 16031
rect 4724 16028 4752 16136
rect 4985 16099 5043 16105
rect 4985 16065 4997 16099
rect 5031 16096 5043 16099
rect 5258 16096 5264 16108
rect 5031 16068 5264 16096
rect 5031 16065 5043 16068
rect 4985 16059 5043 16065
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 7116 16096 7144 16136
rect 7392 16136 10088 16164
rect 7392 16096 7420 16136
rect 7116 16068 7420 16096
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16096 7527 16099
rect 7650 16096 7656 16108
rect 7515 16068 7656 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 7650 16056 7656 16068
rect 7708 16056 7714 16108
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 8202 16096 8208 16108
rect 7800 16068 8208 16096
rect 7800 16056 7806 16068
rect 8202 16056 8208 16068
rect 8260 16096 8266 16108
rect 8481 16099 8539 16105
rect 8481 16096 8493 16099
rect 8260 16068 8493 16096
rect 8260 16056 8266 16068
rect 8481 16065 8493 16068
rect 8527 16065 8539 16099
rect 8481 16059 8539 16065
rect 9585 16099 9643 16105
rect 9585 16065 9597 16099
rect 9631 16096 9643 16099
rect 13924 16096 13952 16195
rect 15562 16192 15568 16204
rect 15620 16192 15626 16244
rect 15580 16096 15608 16192
rect 9631 16068 10180 16096
rect 13924 16068 14320 16096
rect 15580 16068 15976 16096
rect 9631 16065 9643 16068
rect 9585 16059 9643 16065
rect 1765 15991 1823 15997
rect 2792 16000 4752 16028
rect 4801 16031 4859 16037
rect 1780 15960 1808 15991
rect 2792 15960 2820 16000
rect 4801 15997 4813 16031
rect 4847 16028 4859 16031
rect 5074 16028 5080 16040
rect 4847 16000 5080 16028
rect 4847 15997 4859 16000
rect 4801 15991 4859 15997
rect 5074 15988 5080 16000
rect 5132 15988 5138 16040
rect 5537 16031 5595 16037
rect 5537 15997 5549 16031
rect 5583 16028 5595 16031
rect 8570 16028 8576 16040
rect 5583 16000 8576 16028
rect 5583 15997 5595 16000
rect 5537 15991 5595 15997
rect 8570 15988 8576 16000
rect 8628 15988 8634 16040
rect 9401 16031 9459 16037
rect 9401 15997 9413 16031
rect 9447 16028 9459 16031
rect 9674 16028 9680 16040
rect 9447 16000 9680 16028
rect 9447 15997 9459 16000
rect 9401 15991 9459 15997
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 9858 15988 9864 16040
rect 9916 16028 9922 16040
rect 10045 16031 10103 16037
rect 10045 16028 10057 16031
rect 9916 16000 10057 16028
rect 9916 15988 9922 16000
rect 10045 15997 10057 16000
rect 10091 15997 10103 16031
rect 10152 16028 10180 16068
rect 10301 16031 10359 16037
rect 10301 16028 10313 16031
rect 10152 16000 10313 16028
rect 10045 15991 10103 15997
rect 10301 15997 10313 16000
rect 10347 16028 10359 16031
rect 10870 16028 10876 16040
rect 10347 16000 10876 16028
rect 10347 15997 10359 16000
rect 10301 15991 10359 15997
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 15997 12311 16031
rect 12526 16028 12532 16040
rect 12487 16000 12532 16028
rect 12253 15991 12311 15997
rect 1780 15932 2820 15960
rect 2860 15963 2918 15969
rect 2860 15929 2872 15963
rect 2906 15960 2918 15963
rect 3234 15960 3240 15972
rect 2906 15932 3240 15960
rect 2906 15929 2918 15932
rect 2860 15923 2918 15929
rect 3234 15920 3240 15932
rect 3292 15960 3298 15972
rect 3694 15960 3700 15972
rect 3292 15932 3700 15960
rect 3292 15920 3298 15932
rect 3694 15920 3700 15932
rect 3752 15920 3758 15972
rect 4709 15963 4767 15969
rect 4709 15929 4721 15963
rect 4755 15960 4767 15963
rect 5442 15960 5448 15972
rect 4755 15932 5448 15960
rect 4755 15929 4767 15932
rect 4709 15923 4767 15929
rect 5442 15920 5448 15932
rect 5500 15920 5506 15972
rect 7285 15963 7343 15969
rect 7285 15929 7297 15963
rect 7331 15960 7343 15963
rect 9493 15963 9551 15969
rect 7331 15932 7972 15960
rect 7331 15929 7343 15932
rect 7285 15923 7343 15929
rect 566 15852 572 15904
rect 624 15892 630 15904
rect 2774 15892 2780 15904
rect 624 15864 2780 15892
rect 624 15852 630 15864
rect 2774 15852 2780 15864
rect 2832 15852 2838 15904
rect 4890 15852 4896 15904
rect 4948 15892 4954 15904
rect 7190 15892 7196 15904
rect 4948 15864 7196 15892
rect 4948 15852 4954 15864
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 7377 15895 7435 15901
rect 7377 15861 7389 15895
rect 7423 15892 7435 15895
rect 7650 15892 7656 15904
rect 7423 15864 7656 15892
rect 7423 15861 7435 15864
rect 7377 15855 7435 15861
rect 7650 15852 7656 15864
rect 7708 15852 7714 15904
rect 7944 15901 7972 15932
rect 9493 15929 9505 15963
rect 9539 15960 9551 15963
rect 9766 15960 9772 15972
rect 9539 15932 9772 15960
rect 9539 15929 9551 15932
rect 9493 15923 9551 15929
rect 9766 15920 9772 15932
rect 9824 15920 9830 15972
rect 12268 15960 12296 15991
rect 12526 15988 12532 16000
rect 12584 16028 12590 16040
rect 14185 16031 14243 16037
rect 14185 16028 14197 16031
rect 12584 16000 14197 16028
rect 12584 15988 12590 16000
rect 14185 15997 14197 16000
rect 14231 15997 14243 16031
rect 14292 16028 14320 16068
rect 14458 16037 14464 16040
rect 14441 16031 14464 16037
rect 14441 16028 14453 16031
rect 14292 16000 14453 16028
rect 14185 15991 14243 15997
rect 14441 15997 14453 16000
rect 14516 16028 14522 16040
rect 15838 16028 15844 16040
rect 14516 16000 14589 16028
rect 15799 16000 15844 16028
rect 14441 15991 14464 15997
rect 14458 15988 14464 15991
rect 14516 15988 14522 16000
rect 15838 15988 15844 16000
rect 15896 15988 15902 16040
rect 15948 16028 15976 16068
rect 16850 16056 16856 16108
rect 16908 16096 16914 16108
rect 18233 16099 18291 16105
rect 18233 16096 18245 16099
rect 16908 16068 18245 16096
rect 16908 16056 16914 16068
rect 18233 16065 18245 16068
rect 18279 16065 18291 16099
rect 18233 16059 18291 16065
rect 18598 16056 18604 16108
rect 18656 16096 18662 16108
rect 18877 16099 18935 16105
rect 18877 16096 18889 16099
rect 18656 16068 18889 16096
rect 18656 16056 18662 16068
rect 18877 16065 18889 16068
rect 18923 16065 18935 16099
rect 18877 16059 18935 16065
rect 16097 16031 16155 16037
rect 16097 16028 16109 16031
rect 15948 16000 16109 16028
rect 16097 15997 16109 16000
rect 16143 15997 16155 16031
rect 18046 16028 18052 16040
rect 18007 16000 18052 16028
rect 16097 15991 16155 15997
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 19518 16028 19524 16040
rect 18984 16000 19524 16028
rect 12268 15932 12664 15960
rect 7929 15895 7987 15901
rect 7929 15861 7941 15895
rect 7975 15861 7987 15895
rect 8294 15892 8300 15904
rect 8255 15864 8300 15892
rect 7929 15855 7987 15861
rect 8294 15852 8300 15864
rect 8352 15852 8358 15904
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 9033 15895 9091 15901
rect 8444 15864 8489 15892
rect 8444 15852 8450 15864
rect 9033 15861 9045 15895
rect 9079 15892 9091 15895
rect 11238 15892 11244 15904
rect 9079 15864 11244 15892
rect 9079 15861 9091 15864
rect 9033 15855 9091 15861
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 11425 15895 11483 15901
rect 11425 15861 11437 15895
rect 11471 15892 11483 15895
rect 11882 15892 11888 15904
rect 11471 15864 11888 15892
rect 11471 15861 11483 15864
rect 11425 15855 11483 15861
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 12069 15895 12127 15901
rect 12069 15861 12081 15895
rect 12115 15892 12127 15895
rect 12250 15892 12256 15904
rect 12115 15864 12256 15892
rect 12115 15861 12127 15864
rect 12069 15855 12127 15861
rect 12250 15852 12256 15864
rect 12308 15892 12314 15904
rect 12526 15892 12532 15904
rect 12308 15864 12532 15892
rect 12308 15852 12314 15864
rect 12526 15852 12532 15864
rect 12584 15852 12590 15904
rect 12636 15892 12664 15932
rect 12710 15920 12716 15972
rect 12768 15969 12774 15972
rect 12768 15963 12832 15969
rect 12768 15929 12786 15963
rect 12820 15929 12832 15963
rect 12768 15923 12832 15929
rect 12768 15920 12774 15923
rect 15470 15920 15476 15972
rect 15528 15960 15534 15972
rect 18984 15960 19012 16000
rect 19518 15988 19524 16000
rect 19576 15988 19582 16040
rect 20530 16028 20536 16040
rect 20491 16000 20536 16028
rect 20530 15988 20536 16000
rect 20588 15988 20594 16040
rect 15528 15932 19012 15960
rect 19144 15963 19202 15969
rect 15528 15920 15534 15932
rect 19144 15929 19156 15963
rect 19190 15960 19202 15963
rect 19426 15960 19432 15972
rect 19190 15932 19432 15960
rect 19190 15929 19202 15932
rect 19144 15923 19202 15929
rect 19426 15920 19432 15932
rect 19484 15920 19490 15972
rect 20806 15960 20812 15972
rect 20767 15932 20812 15960
rect 20806 15920 20812 15932
rect 20864 15920 20870 15972
rect 13722 15892 13728 15904
rect 12636 15864 13728 15892
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 16390 15852 16396 15904
rect 16448 15892 16454 15904
rect 17221 15895 17279 15901
rect 17221 15892 17233 15895
rect 16448 15864 17233 15892
rect 16448 15852 16454 15864
rect 17221 15861 17233 15864
rect 17267 15861 17279 15895
rect 17221 15855 17279 15861
rect 17497 15895 17555 15901
rect 17497 15861 17509 15895
rect 17543 15892 17555 15895
rect 18966 15892 18972 15904
rect 17543 15864 18972 15892
rect 17543 15861 17555 15864
rect 17497 15855 17555 15861
rect 18966 15852 18972 15864
rect 19024 15852 19030 15904
rect 19058 15852 19064 15904
rect 19116 15892 19122 15904
rect 20257 15895 20315 15901
rect 20257 15892 20269 15895
rect 19116 15864 20269 15892
rect 19116 15852 19122 15864
rect 20257 15861 20269 15864
rect 20303 15861 20315 15895
rect 20257 15855 20315 15861
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 2409 15691 2467 15697
rect 2409 15657 2421 15691
rect 2455 15657 2467 15691
rect 2409 15651 2467 15657
rect 2424 15620 2452 15651
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 2869 15691 2927 15697
rect 2869 15688 2881 15691
rect 2832 15660 2881 15688
rect 2832 15648 2838 15660
rect 2869 15657 2881 15660
rect 2915 15657 2927 15691
rect 2869 15651 2927 15657
rect 3970 15648 3976 15700
rect 4028 15688 4034 15700
rect 4065 15691 4123 15697
rect 4065 15688 4077 15691
rect 4028 15660 4077 15688
rect 4028 15648 4034 15660
rect 4065 15657 4077 15660
rect 4111 15657 4123 15691
rect 4065 15651 4123 15657
rect 4433 15691 4491 15697
rect 4433 15657 4445 15691
rect 4479 15688 4491 15691
rect 5077 15691 5135 15697
rect 5077 15688 5089 15691
rect 4479 15660 5089 15688
rect 4479 15657 4491 15660
rect 4433 15651 4491 15657
rect 5077 15657 5089 15660
rect 5123 15657 5135 15691
rect 5077 15651 5135 15657
rect 5350 15648 5356 15700
rect 5408 15688 5414 15700
rect 5408 15660 5755 15688
rect 5408 15648 5414 15660
rect 3050 15620 3056 15632
rect 2424 15592 3056 15620
rect 3050 15580 3056 15592
rect 3108 15580 3114 15632
rect 3694 15580 3700 15632
rect 3752 15620 3758 15632
rect 5258 15620 5264 15632
rect 3752 15592 5264 15620
rect 3752 15580 3758 15592
rect 5258 15580 5264 15592
rect 5316 15620 5322 15632
rect 5316 15592 5672 15620
rect 5316 15580 5322 15592
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15521 1823 15555
rect 1765 15515 1823 15521
rect 1780 15416 1808 15515
rect 2406 15512 2412 15564
rect 2464 15552 2470 15564
rect 2777 15555 2835 15561
rect 2777 15552 2789 15555
rect 2464 15524 2789 15552
rect 2464 15512 2470 15524
rect 2777 15521 2789 15524
rect 2823 15521 2835 15555
rect 2777 15515 2835 15521
rect 3513 15555 3571 15561
rect 3513 15521 3525 15555
rect 3559 15552 3571 15555
rect 5445 15555 5503 15561
rect 5445 15552 5457 15555
rect 3559 15524 5457 15552
rect 3559 15521 3571 15524
rect 3513 15515 3571 15521
rect 5445 15521 5457 15524
rect 5491 15521 5503 15555
rect 5445 15515 5503 15521
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 3234 15484 3240 15496
rect 3099 15456 3240 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 4525 15487 4583 15493
rect 4525 15484 4537 15487
rect 4212 15456 4537 15484
rect 4212 15444 4218 15456
rect 4525 15453 4537 15456
rect 4571 15453 4583 15487
rect 4706 15484 4712 15496
rect 4667 15456 4712 15484
rect 4525 15447 4583 15453
rect 4706 15444 4712 15456
rect 4764 15444 4770 15496
rect 5534 15484 5540 15496
rect 5495 15456 5540 15484
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 5644 15493 5672 15592
rect 5727 15552 5755 15660
rect 6178 15648 6184 15700
rect 6236 15688 6242 15700
rect 10410 15688 10416 15700
rect 6236 15660 10416 15688
rect 6236 15648 6242 15660
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 10870 15648 10876 15700
rect 10928 15688 10934 15700
rect 11057 15691 11115 15697
rect 11057 15688 11069 15691
rect 10928 15660 11069 15688
rect 10928 15648 10934 15660
rect 11057 15657 11069 15660
rect 11103 15657 11115 15691
rect 11057 15651 11115 15657
rect 11333 15691 11391 15697
rect 11333 15657 11345 15691
rect 11379 15688 11391 15691
rect 12713 15691 12771 15697
rect 11379 15660 12388 15688
rect 11379 15657 11391 15660
rect 11333 15651 11391 15657
rect 7101 15623 7159 15629
rect 7101 15589 7113 15623
rect 7147 15620 7159 15623
rect 8294 15620 8300 15632
rect 7147 15592 8300 15620
rect 7147 15589 7159 15592
rect 7101 15583 7159 15589
rect 8294 15580 8300 15592
rect 8352 15580 8358 15632
rect 9600 15592 11100 15620
rect 7190 15552 7196 15564
rect 5727 15524 7196 15552
rect 7190 15512 7196 15524
rect 7248 15552 7254 15564
rect 7929 15555 7987 15561
rect 7929 15552 7941 15555
rect 7248 15524 7941 15552
rect 7248 15512 7254 15524
rect 7929 15521 7941 15524
rect 7975 15521 7987 15555
rect 7929 15515 7987 15521
rect 8110 15512 8116 15564
rect 8168 15552 8174 15564
rect 9600 15552 9628 15592
rect 8168 15524 9628 15552
rect 9677 15555 9735 15561
rect 8168 15512 8174 15524
rect 9677 15521 9689 15555
rect 9723 15552 9735 15555
rect 9766 15552 9772 15564
rect 9723 15524 9772 15552
rect 9723 15521 9735 15524
rect 9677 15515 9735 15521
rect 9766 15512 9772 15524
rect 9824 15512 9830 15564
rect 9944 15555 10002 15561
rect 9944 15521 9956 15555
rect 9990 15552 10002 15555
rect 10318 15552 10324 15564
rect 9990 15524 10324 15552
rect 9990 15521 10002 15524
rect 9944 15515 10002 15521
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 5629 15487 5687 15493
rect 5629 15453 5641 15487
rect 5675 15453 5687 15487
rect 5629 15447 5687 15453
rect 7466 15444 7472 15496
rect 7524 15484 7530 15496
rect 8021 15487 8079 15493
rect 8021 15484 8033 15487
rect 7524 15456 8033 15484
rect 7524 15444 7530 15456
rect 8021 15453 8033 15456
rect 8067 15453 8079 15487
rect 8202 15484 8208 15496
rect 8163 15456 8208 15484
rect 8021 15447 8079 15453
rect 8202 15444 8208 15456
rect 8260 15444 8266 15496
rect 5350 15416 5356 15428
rect 1780 15388 5356 15416
rect 5350 15376 5356 15388
rect 5408 15376 5414 15428
rect 7561 15419 7619 15425
rect 7561 15385 7573 15419
rect 7607 15416 7619 15419
rect 7650 15416 7656 15428
rect 7607 15388 7656 15416
rect 7607 15385 7619 15388
rect 7561 15379 7619 15385
rect 7650 15376 7656 15388
rect 7708 15376 7714 15428
rect 7834 15376 7840 15428
rect 7892 15416 7898 15428
rect 8570 15416 8576 15428
rect 7892 15388 8576 15416
rect 7892 15376 7898 15388
rect 8570 15376 8576 15388
rect 8628 15376 8634 15428
rect 11072 15416 11100 15592
rect 11238 15580 11244 15632
rect 11296 15620 11302 15632
rect 11793 15623 11851 15629
rect 11793 15620 11805 15623
rect 11296 15592 11805 15620
rect 11296 15580 11302 15592
rect 11793 15589 11805 15592
rect 11839 15589 11851 15623
rect 11793 15583 11851 15589
rect 11698 15552 11704 15564
rect 11659 15524 11704 15552
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 12360 15552 12388 15660
rect 12713 15657 12725 15691
rect 12759 15688 12771 15691
rect 12802 15688 12808 15700
rect 12759 15660 12808 15688
rect 12759 15657 12771 15660
rect 12713 15651 12771 15657
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 14090 15688 14096 15700
rect 14051 15660 14096 15688
rect 14090 15648 14096 15660
rect 14148 15648 14154 15700
rect 14461 15691 14519 15697
rect 14461 15657 14473 15691
rect 14507 15688 14519 15691
rect 15286 15688 15292 15700
rect 14507 15660 15292 15688
rect 14507 15657 14519 15660
rect 14461 15651 14519 15657
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 16761 15691 16819 15697
rect 16761 15657 16773 15691
rect 16807 15688 16819 15691
rect 18046 15688 18052 15700
rect 16807 15660 18052 15688
rect 16807 15657 16819 15660
rect 16761 15651 16819 15657
rect 18046 15648 18052 15660
rect 18104 15648 18110 15700
rect 18141 15691 18199 15697
rect 18141 15657 18153 15691
rect 18187 15688 18199 15691
rect 18601 15691 18659 15697
rect 18601 15688 18613 15691
rect 18187 15660 18613 15688
rect 18187 15657 18199 15660
rect 18141 15651 18199 15657
rect 18601 15657 18613 15660
rect 18647 15657 18659 15691
rect 18782 15688 18788 15700
rect 18743 15660 18788 15688
rect 18601 15651 18659 15657
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 19153 15691 19211 15697
rect 19153 15657 19165 15691
rect 19199 15688 19211 15691
rect 20898 15688 20904 15700
rect 19199 15660 20904 15688
rect 19199 15657 19211 15660
rect 19153 15651 19211 15657
rect 20898 15648 20904 15660
rect 20956 15648 20962 15700
rect 16117 15623 16175 15629
rect 16117 15589 16129 15623
rect 16163 15620 16175 15623
rect 16206 15620 16212 15632
rect 16163 15592 16212 15620
rect 16163 15589 16175 15592
rect 16117 15583 16175 15589
rect 16206 15580 16212 15592
rect 16264 15580 16270 15632
rect 17129 15623 17187 15629
rect 17129 15589 17141 15623
rect 17175 15620 17187 15623
rect 17175 15592 18736 15620
rect 17175 15589 17187 15592
rect 17129 15583 17187 15589
rect 13357 15555 13415 15561
rect 13357 15552 13369 15555
rect 12360 15524 13369 15552
rect 13357 15521 13369 15524
rect 13403 15521 13415 15555
rect 13357 15515 13415 15521
rect 14458 15512 14464 15564
rect 14516 15552 14522 15564
rect 15289 15555 15347 15561
rect 14516 15524 14688 15552
rect 14516 15512 14522 15524
rect 11882 15444 11888 15496
rect 11940 15484 11946 15496
rect 12802 15484 12808 15496
rect 11940 15456 11985 15484
rect 12763 15456 12808 15484
rect 11940 15444 11946 15456
rect 12802 15444 12808 15456
rect 12860 15444 12866 15496
rect 12986 15484 12992 15496
rect 12947 15456 12992 15484
rect 12986 15444 12992 15456
rect 13044 15444 13050 15496
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 13541 15487 13599 15493
rect 13541 15484 13553 15487
rect 13320 15456 13553 15484
rect 13320 15444 13326 15456
rect 13541 15453 13553 15456
rect 13587 15453 13599 15487
rect 14550 15484 14556 15496
rect 14511 15456 14556 15484
rect 13541 15447 13599 15453
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 14660 15493 14688 15524
rect 15289 15521 15301 15555
rect 15335 15552 15347 15555
rect 16022 15552 16028 15564
rect 15335 15524 16028 15552
rect 15335 15521 15347 15524
rect 15289 15515 15347 15521
rect 16022 15512 16028 15524
rect 16080 15512 16086 15564
rect 16482 15552 16488 15564
rect 16224 15524 16488 15552
rect 16224 15493 16252 15524
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 17494 15552 17500 15564
rect 16592 15524 17500 15552
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 16209 15487 16267 15493
rect 16209 15453 16221 15487
rect 16255 15453 16267 15487
rect 16390 15484 16396 15496
rect 16351 15456 16396 15484
rect 16209 15447 16267 15453
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 12345 15419 12403 15425
rect 11072 15388 11744 15416
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 4890 15348 4896 15360
rect 4764 15320 4896 15348
rect 4764 15308 4770 15320
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 5534 15308 5540 15360
rect 5592 15348 5598 15360
rect 11606 15348 11612 15360
rect 5592 15320 11612 15348
rect 5592 15308 5598 15320
rect 11606 15308 11612 15320
rect 11664 15308 11670 15360
rect 11716 15348 11744 15388
rect 12345 15385 12357 15419
rect 12391 15416 12403 15419
rect 15470 15416 15476 15428
rect 12391 15388 15476 15416
rect 12391 15385 12403 15388
rect 12345 15379 12403 15385
rect 15470 15376 15476 15388
rect 15528 15376 15534 15428
rect 16592 15416 16620 15524
rect 17494 15512 17500 15524
rect 17552 15512 17558 15564
rect 18233 15555 18291 15561
rect 18233 15521 18245 15555
rect 18279 15552 18291 15555
rect 18598 15552 18604 15564
rect 18279 15524 18604 15552
rect 18279 15521 18291 15524
rect 18233 15515 18291 15521
rect 18598 15512 18604 15524
rect 18656 15512 18662 15564
rect 18708 15496 18736 15592
rect 19058 15512 19064 15564
rect 19116 15552 19122 15564
rect 20162 15552 20168 15564
rect 19116 15524 19380 15552
rect 20123 15524 20168 15552
rect 19116 15512 19122 15524
rect 16666 15444 16672 15496
rect 16724 15484 16730 15496
rect 17221 15487 17279 15493
rect 17221 15484 17233 15487
rect 16724 15456 17233 15484
rect 16724 15444 16730 15456
rect 17221 15453 17233 15456
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 17405 15487 17463 15493
rect 17405 15453 17417 15487
rect 17451 15453 17463 15487
rect 17405 15447 17463 15453
rect 15580 15388 16620 15416
rect 17420 15416 17448 15447
rect 17586 15444 17592 15496
rect 17644 15484 17650 15496
rect 18325 15487 18383 15493
rect 18325 15484 18337 15487
rect 17644 15456 18337 15484
rect 17644 15444 17650 15456
rect 18325 15453 18337 15456
rect 18371 15453 18383 15487
rect 18325 15447 18383 15453
rect 18690 15444 18696 15496
rect 18748 15444 18754 15496
rect 19242 15484 19248 15496
rect 19203 15456 19248 15484
rect 19242 15444 19248 15456
rect 19300 15444 19306 15496
rect 19352 15493 19380 15524
rect 20162 15512 20168 15524
rect 20220 15512 20226 15564
rect 19337 15487 19395 15493
rect 19337 15453 19349 15487
rect 19383 15484 19395 15487
rect 20254 15484 20260 15496
rect 19383 15456 20116 15484
rect 20215 15456 20260 15484
rect 19383 15453 19395 15456
rect 19337 15447 19395 15453
rect 18506 15416 18512 15428
rect 17420 15388 18512 15416
rect 15580 15348 15608 15388
rect 18506 15376 18512 15388
rect 18564 15376 18570 15428
rect 19150 15376 19156 15428
rect 19208 15416 19214 15428
rect 19797 15419 19855 15425
rect 19797 15416 19809 15419
rect 19208 15388 19809 15416
rect 19208 15376 19214 15388
rect 19797 15385 19809 15388
rect 19843 15385 19855 15419
rect 20088 15416 20116 15456
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15453 20407 15487
rect 20349 15447 20407 15453
rect 20364 15416 20392 15447
rect 20088 15388 20392 15416
rect 19797 15379 19855 15385
rect 11716 15320 15608 15348
rect 15749 15351 15807 15357
rect 15749 15317 15761 15351
rect 15795 15348 15807 15351
rect 16298 15348 16304 15360
rect 15795 15320 16304 15348
rect 15795 15317 15807 15320
rect 15749 15311 15807 15317
rect 16298 15308 16304 15320
rect 16356 15308 16362 15360
rect 17310 15308 17316 15360
rect 17368 15348 17374 15360
rect 17773 15351 17831 15357
rect 17773 15348 17785 15351
rect 17368 15320 17785 15348
rect 17368 15308 17374 15320
rect 17773 15317 17785 15320
rect 17819 15317 17831 15351
rect 17773 15311 17831 15317
rect 18601 15351 18659 15357
rect 18601 15317 18613 15351
rect 18647 15348 18659 15351
rect 19610 15348 19616 15360
rect 18647 15320 19616 15348
rect 18647 15317 18659 15320
rect 18601 15311 18659 15317
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 4433 15147 4491 15153
rect 4433 15144 4445 15147
rect 1504 15116 4445 15144
rect 1504 14949 1532 15116
rect 4433 15113 4445 15116
rect 4479 15113 4491 15147
rect 4433 15107 4491 15113
rect 7282 15104 7288 15156
rect 7340 15144 7346 15156
rect 7650 15144 7656 15156
rect 7340 15116 7656 15144
rect 7340 15104 7346 15116
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 7834 15144 7840 15156
rect 7795 15116 7840 15144
rect 7834 15104 7840 15116
rect 7892 15104 7898 15156
rect 9950 15144 9956 15156
rect 7944 15116 9956 15144
rect 3605 15079 3663 15085
rect 3605 15045 3617 15079
rect 3651 15076 3663 15079
rect 3694 15076 3700 15088
rect 3651 15048 3700 15076
rect 3651 15045 3663 15048
rect 3605 15039 3663 15045
rect 3694 15036 3700 15048
rect 3752 15036 3758 15088
rect 1762 15008 1768 15020
rect 1723 14980 1768 15008
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 2222 15008 2228 15020
rect 2183 14980 2228 15008
rect 2222 14968 2228 14980
rect 2280 14968 2286 15020
rect 5077 15011 5135 15017
rect 5077 14977 5089 15011
rect 5123 15008 5135 15011
rect 5810 15008 5816 15020
rect 5123 14980 5816 15008
rect 5123 14977 5135 14980
rect 5077 14971 5135 14977
rect 5810 14968 5816 14980
rect 5868 14968 5874 15020
rect 7469 15011 7527 15017
rect 7469 14977 7481 15011
rect 7515 15008 7527 15011
rect 7742 15008 7748 15020
rect 7515 14980 7748 15008
rect 7515 14977 7527 14980
rect 7469 14971 7527 14977
rect 7742 14968 7748 14980
rect 7800 14968 7806 15020
rect 1489 14943 1547 14949
rect 1489 14909 1501 14943
rect 1535 14909 1547 14943
rect 1489 14903 1547 14909
rect 7193 14943 7251 14949
rect 7193 14909 7205 14943
rect 7239 14940 7251 14943
rect 7944 14940 7972 15116
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 10413 15147 10471 15153
rect 10413 15113 10425 15147
rect 10459 15144 10471 15147
rect 11698 15144 11704 15156
rect 10459 15116 11704 15144
rect 10459 15113 10471 15116
rect 10413 15107 10471 15113
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 12802 15144 12808 15156
rect 11808 15116 12808 15144
rect 8389 15079 8447 15085
rect 8389 15045 8401 15079
rect 8435 15076 8447 15079
rect 11808 15076 11836 15116
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 14274 15144 14280 15156
rect 14235 15116 14280 15144
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 14550 15104 14556 15156
rect 14608 15144 14614 15156
rect 14645 15147 14703 15153
rect 14645 15144 14657 15147
rect 14608 15116 14657 15144
rect 14608 15104 14614 15116
rect 14645 15113 14657 15116
rect 14691 15113 14703 15147
rect 14645 15107 14703 15113
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 15562 15144 15568 15156
rect 14792 15116 15568 15144
rect 14792 15104 14798 15116
rect 15562 15104 15568 15116
rect 15620 15104 15626 15156
rect 17954 15144 17960 15156
rect 16040 15116 17960 15144
rect 8435 15048 11836 15076
rect 11977 15079 12035 15085
rect 8435 15045 8447 15048
rect 8389 15039 8447 15045
rect 11977 15045 11989 15079
rect 12023 15076 12035 15079
rect 16040 15076 16068 15116
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 19426 15144 19432 15156
rect 19387 15116 19432 15144
rect 19426 15104 19432 15116
rect 19484 15104 19490 15156
rect 19705 15147 19763 15153
rect 19705 15113 19717 15147
rect 19751 15144 19763 15147
rect 20254 15144 20260 15156
rect 19751 15116 20260 15144
rect 19751 15113 19763 15116
rect 19705 15107 19763 15113
rect 20254 15104 20260 15116
rect 20312 15104 20318 15156
rect 20622 15104 20628 15156
rect 20680 15144 20686 15156
rect 20901 15147 20959 15153
rect 20901 15144 20913 15147
rect 20680 15116 20913 15144
rect 20680 15104 20686 15116
rect 20901 15113 20913 15116
rect 20947 15113 20959 15147
rect 20901 15107 20959 15113
rect 12023 15048 16068 15076
rect 12023 15045 12035 15048
rect 11977 15039 12035 15045
rect 9033 15011 9091 15017
rect 9033 14977 9045 15011
rect 9079 15008 9091 15011
rect 9858 15008 9864 15020
rect 9079 14980 9864 15008
rect 9079 14977 9091 14980
rect 9033 14971 9091 14977
rect 9858 14968 9864 14980
rect 9916 14968 9922 15020
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 15008 10103 15011
rect 10318 15008 10324 15020
rect 10091 14980 10324 15008
rect 10091 14977 10103 14980
rect 10045 14971 10103 14977
rect 10318 14968 10324 14980
rect 10376 14968 10382 15020
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 10928 14980 10977 15008
rect 10928 14968 10934 14980
rect 10965 14977 10977 14980
rect 11011 14977 11023 15011
rect 12894 15008 12900 15020
rect 10965 14971 11023 14977
rect 11072 14980 12900 15008
rect 7239 14912 7972 14940
rect 8021 14943 8079 14949
rect 7239 14909 7251 14912
rect 7193 14903 7251 14909
rect 8021 14909 8033 14943
rect 8067 14940 8079 14943
rect 8202 14940 8208 14952
rect 8067 14912 8208 14940
rect 8067 14909 8079 14912
rect 8021 14903 8079 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 11072 14940 11100 14980
rect 12894 14968 12900 14980
rect 12952 15008 12958 15020
rect 13170 15008 13176 15020
rect 12952 14980 13176 15008
rect 12952 14968 12958 14980
rect 13170 14968 13176 14980
rect 13228 14968 13234 15020
rect 13265 15011 13323 15017
rect 13265 14977 13277 15011
rect 13311 15008 13323 15011
rect 13630 15008 13636 15020
rect 13311 14980 13636 15008
rect 13311 14977 13323 14980
rect 13265 14971 13323 14977
rect 13630 14968 13636 14980
rect 13688 14968 13694 15020
rect 14734 15008 14740 15020
rect 14108 14980 14740 15008
rect 8352 14912 11100 14940
rect 8352 14900 8358 14912
rect 11606 14900 11612 14952
rect 11664 14940 11670 14952
rect 11793 14943 11851 14949
rect 11793 14940 11805 14943
rect 11664 14912 11805 14940
rect 11664 14900 11670 14912
rect 11793 14909 11805 14912
rect 11839 14909 11851 14943
rect 11793 14903 11851 14909
rect 13814 14900 13820 14952
rect 13872 14940 13878 14952
rect 14108 14949 14136 14980
rect 14734 14968 14740 14980
rect 14792 14968 14798 15020
rect 15194 15008 15200 15020
rect 15155 14980 15200 15008
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 15838 14968 15844 15020
rect 15896 15008 15902 15020
rect 16032 15011 16090 15017
rect 16032 15008 16044 15011
rect 15896 14980 16044 15008
rect 15896 14968 15902 14980
rect 16032 14977 16044 14980
rect 16078 14977 16090 15011
rect 19444 15008 19472 15104
rect 20257 15011 20315 15017
rect 20257 15008 20269 15011
rect 19444 14980 20269 15008
rect 16032 14971 16090 14977
rect 20257 14977 20269 14980
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 13872 14912 14105 14940
rect 13872 14900 13878 14912
rect 14093 14909 14105 14912
rect 14139 14909 14151 14943
rect 15933 14943 15991 14949
rect 15933 14940 15945 14943
rect 14093 14903 14151 14909
rect 14384 14912 15945 14940
rect 2492 14875 2550 14881
rect 2492 14841 2504 14875
rect 2538 14872 2550 14875
rect 3234 14872 3240 14884
rect 2538 14844 3240 14872
rect 2538 14841 2550 14844
rect 2492 14835 2550 14841
rect 3234 14832 3240 14844
rect 3292 14832 3298 14884
rect 7285 14875 7343 14881
rect 7285 14841 7297 14875
rect 7331 14872 7343 14875
rect 7558 14872 7564 14884
rect 7331 14844 7564 14872
rect 7331 14841 7343 14844
rect 7285 14835 7343 14841
rect 7558 14832 7564 14844
rect 7616 14832 7622 14884
rect 8757 14875 8815 14881
rect 8757 14841 8769 14875
rect 8803 14872 8815 14875
rect 9122 14872 9128 14884
rect 8803 14844 9128 14872
rect 8803 14841 8815 14844
rect 8757 14835 8815 14841
rect 9122 14832 9128 14844
rect 9180 14832 9186 14884
rect 10781 14875 10839 14881
rect 10781 14872 10793 14875
rect 9416 14844 10793 14872
rect 4798 14804 4804 14816
rect 4759 14776 4804 14804
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 4893 14807 4951 14813
rect 4893 14773 4905 14807
rect 4939 14804 4951 14807
rect 5350 14804 5356 14816
rect 4939 14776 5356 14804
rect 4939 14773 4951 14776
rect 4893 14767 4951 14773
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7650 14764 7656 14816
rect 7708 14804 7714 14816
rect 8846 14804 8852 14816
rect 7708 14776 8852 14804
rect 7708 14764 7714 14776
rect 8846 14764 8852 14776
rect 8904 14764 8910 14816
rect 9416 14813 9444 14844
rect 10781 14841 10793 14844
rect 10827 14841 10839 14875
rect 10781 14835 10839 14841
rect 12526 14832 12532 14884
rect 12584 14872 12590 14884
rect 13081 14875 13139 14881
rect 13081 14872 13093 14875
rect 12584 14844 13093 14872
rect 12584 14832 12590 14844
rect 13081 14841 13093 14844
rect 13127 14841 13139 14875
rect 13081 14835 13139 14841
rect 13722 14832 13728 14884
rect 13780 14872 13786 14884
rect 14384 14872 14412 14912
rect 15933 14909 15945 14912
rect 15979 14909 15991 14943
rect 15933 14903 15991 14909
rect 17770 14900 17776 14952
rect 17828 14940 17834 14952
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 17828 14912 18061 14940
rect 17828 14900 17834 14912
rect 18049 14909 18061 14912
rect 18095 14909 18107 14943
rect 20717 14943 20775 14949
rect 20717 14940 20729 14943
rect 18049 14903 18107 14909
rect 18156 14912 20729 14940
rect 13780 14844 14412 14872
rect 15013 14875 15071 14881
rect 13780 14832 13786 14844
rect 15013 14841 15025 14875
rect 15059 14872 15071 14875
rect 16292 14875 16350 14881
rect 15059 14844 16252 14872
rect 15059 14841 15071 14844
rect 15013 14835 15071 14841
rect 9401 14807 9459 14813
rect 9401 14773 9413 14807
rect 9447 14773 9459 14807
rect 9766 14804 9772 14816
rect 9727 14776 9772 14804
rect 9401 14767 9459 14773
rect 9766 14764 9772 14776
rect 9824 14764 9830 14816
rect 9861 14807 9919 14813
rect 9861 14773 9873 14807
rect 9907 14804 9919 14807
rect 10410 14804 10416 14816
rect 9907 14776 10416 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 10870 14804 10876 14816
rect 10831 14776 10876 14804
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 12618 14804 12624 14816
rect 12579 14776 12624 14804
rect 12618 14764 12624 14776
rect 12676 14764 12682 14816
rect 12986 14804 12992 14816
rect 12947 14776 12992 14804
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 15105 14807 15163 14813
rect 15105 14773 15117 14807
rect 15151 14804 15163 14807
rect 15470 14804 15476 14816
rect 15151 14776 15476 14804
rect 15151 14773 15163 14776
rect 15105 14767 15163 14773
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 15749 14807 15807 14813
rect 15749 14773 15761 14807
rect 15795 14804 15807 14807
rect 15838 14804 15844 14816
rect 15795 14776 15844 14804
rect 15795 14773 15807 14776
rect 15749 14767 15807 14773
rect 15838 14764 15844 14776
rect 15896 14804 15902 14816
rect 16114 14804 16120 14816
rect 15896 14776 16120 14804
rect 15896 14764 15902 14776
rect 16114 14764 16120 14776
rect 16172 14764 16178 14816
rect 16224 14804 16252 14844
rect 16292 14841 16304 14875
rect 16338 14872 16350 14875
rect 16390 14872 16396 14884
rect 16338 14844 16396 14872
rect 16338 14841 16350 14844
rect 16292 14835 16350 14841
rect 16390 14832 16396 14844
rect 16448 14832 16454 14884
rect 17494 14832 17500 14884
rect 17552 14872 17558 14884
rect 18156 14872 18184 14912
rect 20717 14909 20729 14912
rect 20763 14909 20775 14943
rect 20717 14903 20775 14909
rect 17552 14844 18184 14872
rect 18316 14875 18374 14881
rect 17552 14832 17558 14844
rect 18316 14841 18328 14875
rect 18362 14872 18374 14875
rect 18506 14872 18512 14884
rect 18362 14844 18512 14872
rect 18362 14841 18374 14844
rect 18316 14835 18374 14841
rect 18506 14832 18512 14844
rect 18564 14832 18570 14884
rect 19702 14832 19708 14884
rect 19760 14872 19766 14884
rect 20165 14875 20223 14881
rect 20165 14872 20177 14875
rect 19760 14844 20177 14872
rect 19760 14832 19766 14844
rect 20165 14841 20177 14844
rect 20211 14841 20223 14875
rect 20165 14835 20223 14841
rect 16850 14804 16856 14816
rect 16224 14776 16856 14804
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 17402 14804 17408 14816
rect 17363 14776 17408 14804
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 19334 14804 19340 14816
rect 18012 14776 19340 14804
rect 18012 14764 18018 14776
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 20073 14807 20131 14813
rect 20073 14773 20085 14807
rect 20119 14804 20131 14807
rect 20346 14804 20352 14816
rect 20119 14776 20352 14804
rect 20119 14773 20131 14776
rect 20073 14767 20131 14773
rect 20346 14764 20352 14776
rect 20404 14764 20410 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 2593 14603 2651 14609
rect 2593 14569 2605 14603
rect 2639 14600 2651 14603
rect 4154 14600 4160 14612
rect 2639 14572 4160 14600
rect 2639 14569 2651 14572
rect 2593 14563 2651 14569
rect 4154 14560 4160 14572
rect 4212 14560 4218 14612
rect 5810 14600 5816 14612
rect 5771 14572 5816 14600
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 8113 14603 8171 14609
rect 8113 14600 8125 14603
rect 7156 14572 8125 14600
rect 7156 14560 7162 14572
rect 8113 14569 8125 14572
rect 8159 14569 8171 14603
rect 8113 14563 8171 14569
rect 8205 14603 8263 14609
rect 8205 14569 8217 14603
rect 8251 14600 8263 14603
rect 8294 14600 8300 14612
rect 8251 14572 8300 14600
rect 8251 14569 8263 14572
rect 8205 14563 8263 14569
rect 5828 14532 5856 14560
rect 6334 14535 6392 14541
rect 6334 14532 6346 14535
rect 2792 14504 3096 14532
rect 1765 14467 1823 14473
rect 1765 14433 1777 14467
rect 1811 14464 1823 14467
rect 1854 14464 1860 14476
rect 1811 14436 1860 14464
rect 1811 14433 1823 14436
rect 1765 14427 1823 14433
rect 1854 14424 1860 14436
rect 1912 14424 1918 14476
rect 2406 14424 2412 14476
rect 2464 14464 2470 14476
rect 2792 14464 2820 14504
rect 2464 14436 2820 14464
rect 2464 14424 2470 14436
rect 2866 14424 2872 14476
rect 2924 14464 2930 14476
rect 3068 14473 3096 14504
rect 4448 14504 5212 14532
rect 5828 14504 6346 14532
rect 2961 14467 3019 14473
rect 2961 14464 2973 14467
rect 2924 14436 2973 14464
rect 2924 14424 2930 14436
rect 2961 14433 2973 14436
rect 3007 14433 3019 14467
rect 2961 14427 3019 14433
rect 3053 14467 3111 14473
rect 3053 14433 3065 14467
rect 3099 14464 3111 14467
rect 3099 14436 3832 14464
rect 3099 14433 3111 14436
rect 3053 14427 3111 14433
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14396 3295 14399
rect 3694 14396 3700 14408
rect 3283 14368 3700 14396
rect 3283 14365 3295 14368
rect 3237 14359 3295 14365
rect 3694 14356 3700 14368
rect 3752 14356 3758 14408
rect 3804 14260 3832 14436
rect 4246 14424 4252 14476
rect 4304 14464 4310 14476
rect 4448 14473 4476 14504
rect 4433 14467 4491 14473
rect 4433 14464 4445 14467
rect 4304 14436 4445 14464
rect 4304 14424 4310 14436
rect 4433 14433 4445 14436
rect 4479 14433 4491 14467
rect 4433 14427 4491 14433
rect 4700 14467 4758 14473
rect 4700 14433 4712 14467
rect 4746 14464 4758 14467
rect 5074 14464 5080 14476
rect 4746 14436 5080 14464
rect 4746 14433 4758 14436
rect 4700 14427 4758 14433
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5184 14464 5212 14504
rect 6334 14501 6346 14504
rect 6380 14501 6392 14535
rect 6334 14495 6392 14501
rect 7558 14492 7564 14544
rect 7616 14532 7622 14544
rect 8128 14532 8156 14563
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 9674 14600 9680 14612
rect 9048 14572 9680 14600
rect 9048 14532 9076 14572
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 10781 14603 10839 14609
rect 10781 14600 10793 14603
rect 9824 14572 10793 14600
rect 9824 14560 9830 14572
rect 10781 14569 10793 14572
rect 10827 14569 10839 14603
rect 10781 14563 10839 14569
rect 11241 14603 11299 14609
rect 11241 14569 11253 14603
rect 11287 14600 11299 14603
rect 12526 14600 12532 14612
rect 11287 14572 12532 14600
rect 11287 14569 11299 14572
rect 11241 14563 11299 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 12676 14572 14657 14600
rect 12676 14560 12682 14572
rect 14645 14569 14657 14572
rect 14691 14569 14703 14603
rect 14645 14563 14703 14569
rect 15565 14603 15623 14609
rect 15565 14569 15577 14603
rect 15611 14600 15623 14603
rect 15654 14600 15660 14612
rect 15611 14572 15660 14600
rect 15611 14569 15623 14572
rect 15565 14563 15623 14569
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 16390 14600 16396 14612
rect 16351 14572 16396 14600
rect 16390 14560 16396 14572
rect 16448 14560 16454 14612
rect 18325 14603 18383 14609
rect 18325 14569 18337 14603
rect 18371 14600 18383 14603
rect 18506 14600 18512 14612
rect 18371 14572 18512 14600
rect 18371 14569 18383 14572
rect 18325 14563 18383 14569
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 18601 14603 18659 14609
rect 18601 14569 18613 14603
rect 18647 14600 18659 14603
rect 18690 14600 18696 14612
rect 18647 14572 18696 14600
rect 18647 14569 18659 14572
rect 18601 14563 18659 14569
rect 18690 14560 18696 14572
rect 18748 14560 18754 14612
rect 18966 14600 18972 14612
rect 18927 14572 18972 14600
rect 18966 14560 18972 14572
rect 19024 14560 19030 14612
rect 19610 14600 19616 14612
rect 19571 14572 19616 14600
rect 19610 14560 19616 14572
rect 19668 14560 19674 14612
rect 7616 14504 8064 14532
rect 8128 14504 9076 14532
rect 7616 14492 7622 14504
rect 5184 14436 5488 14464
rect 5460 14396 5488 14436
rect 5534 14424 5540 14476
rect 5592 14464 5598 14476
rect 8036 14464 8064 14504
rect 9122 14492 9128 14544
rect 9180 14532 9186 14544
rect 10045 14535 10103 14541
rect 10045 14532 10057 14535
rect 9180 14504 10057 14532
rect 9180 14492 9186 14504
rect 10045 14501 10057 14504
rect 10091 14501 10103 14535
rect 10045 14495 10103 14501
rect 10134 14492 10140 14544
rect 10192 14532 10198 14544
rect 12710 14532 12716 14544
rect 10192 14504 12716 14532
rect 10192 14492 10198 14504
rect 12710 14492 12716 14504
rect 12768 14492 12774 14544
rect 16298 14532 16304 14544
rect 16259 14504 16304 14532
rect 16298 14492 16304 14504
rect 16356 14492 16362 14544
rect 16761 14535 16819 14541
rect 16761 14501 16773 14535
rect 16807 14532 16819 14535
rect 17212 14535 17270 14541
rect 17212 14532 17224 14535
rect 16807 14504 17224 14532
rect 16807 14501 16819 14504
rect 16761 14495 16819 14501
rect 17212 14501 17224 14504
rect 17258 14532 17270 14535
rect 17402 14532 17408 14544
rect 17258 14504 17408 14532
rect 17258 14501 17270 14504
rect 17212 14495 17270 14501
rect 17402 14492 17408 14504
rect 17460 14532 17466 14544
rect 17460 14504 19196 14532
rect 17460 14492 17466 14504
rect 9766 14464 9772 14476
rect 5592 14436 7788 14464
rect 8036 14436 9772 14464
rect 5592 14424 5598 14436
rect 7760 14408 7788 14436
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 12526 14473 12532 14476
rect 11609 14467 11667 14473
rect 11609 14464 11621 14467
rect 10008 14436 11621 14464
rect 10008 14424 10014 14436
rect 11609 14433 11621 14436
rect 11655 14433 11667 14467
rect 12520 14464 12532 14473
rect 11609 14427 11667 14433
rect 11900 14436 12532 14464
rect 6089 14399 6147 14405
rect 6089 14396 6101 14399
rect 5460 14368 6101 14396
rect 6089 14365 6101 14368
rect 6135 14365 6147 14399
rect 6089 14359 6147 14365
rect 7742 14356 7748 14408
rect 7800 14396 7806 14408
rect 8297 14399 8355 14405
rect 8297 14396 8309 14399
rect 7800 14368 8309 14396
rect 7800 14356 7806 14368
rect 8297 14365 8309 14368
rect 8343 14365 8355 14399
rect 8297 14359 8355 14365
rect 8846 14356 8852 14408
rect 8904 14396 8910 14408
rect 10137 14399 10195 14405
rect 10137 14396 10149 14399
rect 8904 14368 10149 14396
rect 8904 14356 8910 14368
rect 10137 14365 10149 14368
rect 10183 14365 10195 14399
rect 10137 14359 10195 14365
rect 10226 14356 10232 14408
rect 10284 14396 10290 14408
rect 10284 14368 10329 14396
rect 10284 14356 10290 14368
rect 10502 14356 10508 14408
rect 10560 14396 10566 14408
rect 11900 14405 11928 14436
rect 12520 14427 12532 14436
rect 12526 14424 12532 14427
rect 12584 14424 12590 14476
rect 13998 14424 14004 14476
rect 14056 14464 14062 14476
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 14056 14436 14105 14464
rect 14056 14424 14062 14436
rect 14093 14433 14105 14436
rect 14139 14433 14151 14467
rect 14093 14427 14151 14433
rect 14553 14467 14611 14473
rect 14553 14433 14565 14467
rect 14599 14464 14611 14467
rect 15010 14464 15016 14476
rect 14599 14436 15016 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 15010 14424 15016 14436
rect 15068 14424 15074 14476
rect 15381 14467 15439 14473
rect 15381 14433 15393 14467
rect 15427 14464 15439 14467
rect 15427 14436 15884 14464
rect 15427 14433 15439 14436
rect 15381 14427 15439 14433
rect 11701 14399 11759 14405
rect 11701 14396 11713 14399
rect 10560 14368 11713 14396
rect 10560 14356 10566 14368
rect 11701 14365 11713 14368
rect 11747 14365 11759 14399
rect 11701 14359 11759 14365
rect 11885 14399 11943 14405
rect 11885 14365 11897 14399
rect 11931 14365 11943 14399
rect 12250 14396 12256 14408
rect 12211 14368 12256 14396
rect 11885 14359 11943 14365
rect 12250 14356 12256 14368
rect 12308 14356 12314 14408
rect 14737 14399 14795 14405
rect 14737 14365 14749 14399
rect 14783 14365 14795 14399
rect 14737 14359 14795 14365
rect 7024 14300 11744 14328
rect 7024 14260 7052 14300
rect 11716 14272 11744 14300
rect 13722 14288 13728 14340
rect 13780 14328 13786 14340
rect 13909 14331 13967 14337
rect 13909 14328 13921 14331
rect 13780 14300 13921 14328
rect 13780 14288 13786 14300
rect 13909 14297 13921 14300
rect 13955 14297 13967 14331
rect 13909 14291 13967 14297
rect 14550 14288 14556 14340
rect 14608 14328 14614 14340
rect 14752 14328 14780 14359
rect 14608 14300 14780 14328
rect 14608 14288 14614 14300
rect 3804 14232 7052 14260
rect 7469 14263 7527 14269
rect 7469 14229 7481 14263
rect 7515 14260 7527 14263
rect 7558 14260 7564 14272
rect 7515 14232 7564 14260
rect 7515 14229 7527 14232
rect 7469 14223 7527 14229
rect 7558 14220 7564 14232
rect 7616 14220 7622 14272
rect 7742 14260 7748 14272
rect 7703 14232 7748 14260
rect 7742 14220 7748 14232
rect 7800 14220 7806 14272
rect 9677 14263 9735 14269
rect 9677 14229 9689 14263
rect 9723 14260 9735 14263
rect 10962 14260 10968 14272
rect 9723 14232 10968 14260
rect 9723 14229 9735 14232
rect 9677 14223 9735 14229
rect 10962 14220 10968 14232
rect 11020 14220 11026 14272
rect 11698 14220 11704 14272
rect 11756 14220 11762 14272
rect 13630 14260 13636 14272
rect 13591 14232 13636 14260
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 14185 14263 14243 14269
rect 14185 14229 14197 14263
rect 14231 14260 14243 14263
rect 15102 14260 15108 14272
rect 14231 14232 15108 14260
rect 14231 14229 14243 14232
rect 14185 14223 14243 14229
rect 15102 14220 15108 14232
rect 15160 14220 15166 14272
rect 15856 14260 15884 14436
rect 16482 14424 16488 14476
rect 16540 14464 16546 14476
rect 18782 14464 18788 14476
rect 16540 14436 18788 14464
rect 16540 14424 16546 14436
rect 18782 14424 18788 14436
rect 18840 14464 18846 14476
rect 19061 14467 19119 14473
rect 19061 14464 19073 14467
rect 18840 14436 19073 14464
rect 18840 14424 18846 14436
rect 19061 14433 19073 14436
rect 19107 14433 19119 14467
rect 19061 14427 19119 14433
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14396 16635 14399
rect 16761 14399 16819 14405
rect 16761 14396 16773 14399
rect 16623 14368 16773 14396
rect 16623 14365 16635 14368
rect 16577 14359 16635 14365
rect 16761 14365 16773 14368
rect 16807 14365 16819 14399
rect 16942 14396 16948 14408
rect 16903 14368 16948 14396
rect 16761 14359 16819 14365
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 19168 14405 19196 14504
rect 19981 14467 20039 14473
rect 19981 14433 19993 14467
rect 20027 14464 20039 14467
rect 20622 14464 20628 14476
rect 20027 14436 20628 14464
rect 20027 14433 20039 14436
rect 19981 14427 20039 14433
rect 20622 14424 20628 14436
rect 20680 14424 20686 14476
rect 19153 14399 19211 14405
rect 19153 14365 19165 14399
rect 19199 14365 19211 14399
rect 19153 14359 19211 14365
rect 19334 14356 19340 14408
rect 19392 14396 19398 14408
rect 20073 14399 20131 14405
rect 20073 14396 20085 14399
rect 19392 14368 20085 14396
rect 19392 14356 19398 14368
rect 20073 14365 20085 14368
rect 20119 14365 20131 14399
rect 20073 14359 20131 14365
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14365 20223 14399
rect 20165 14359 20223 14365
rect 15933 14331 15991 14337
rect 15933 14297 15945 14331
rect 15979 14328 15991 14331
rect 16666 14328 16672 14340
rect 15979 14300 16672 14328
rect 15979 14297 15991 14300
rect 15933 14291 15991 14297
rect 16666 14288 16672 14300
rect 16724 14288 16730 14340
rect 18874 14288 18880 14340
rect 18932 14328 18938 14340
rect 20180 14328 20208 14359
rect 18932 14300 20208 14328
rect 18932 14288 18938 14300
rect 19978 14260 19984 14272
rect 15856 14232 19984 14260
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 2593 14059 2651 14065
rect 2593 14025 2605 14059
rect 2639 14056 2651 14059
rect 2774 14056 2780 14068
rect 2639 14028 2780 14056
rect 2639 14025 2651 14028
rect 2593 14019 2651 14025
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 3142 14056 3148 14068
rect 3103 14028 3148 14056
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 3510 14016 3516 14068
rect 3568 14056 3574 14068
rect 5074 14056 5080 14068
rect 3568 14028 4936 14056
rect 5035 14028 5080 14056
rect 3568 14016 3574 14028
rect 4908 13988 4936 14028
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 5350 14056 5356 14068
rect 5311 14028 5356 14056
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 8662 14056 8668 14068
rect 5920 14028 8248 14056
rect 8575 14028 8668 14056
rect 5920 13988 5948 14028
rect 4908 13960 5948 13988
rect 8220 13988 8248 14028
rect 8662 14016 8668 14028
rect 8720 14056 8726 14068
rect 8720 14028 10640 14056
rect 8720 14016 8726 14028
rect 8849 13991 8907 13997
rect 8849 13988 8861 13991
rect 8220 13960 8861 13988
rect 8849 13957 8861 13960
rect 8895 13957 8907 13991
rect 10505 13991 10563 13997
rect 10505 13988 10517 13991
rect 8849 13951 8907 13957
rect 9324 13960 10517 13988
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 5905 13923 5963 13929
rect 5905 13920 5917 13923
rect 5132 13892 5917 13920
rect 5132 13880 5138 13892
rect 5905 13889 5917 13892
rect 5951 13920 5963 13923
rect 5994 13920 6000 13932
rect 5951 13892 6000 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 5994 13880 6000 13892
rect 6052 13880 6058 13932
rect 9324 13929 9352 13960
rect 10505 13957 10517 13960
rect 10551 13957 10563 13991
rect 10612 13988 10640 14028
rect 10870 14016 10876 14068
rect 10928 14056 10934 14068
rect 11333 14059 11391 14065
rect 11333 14056 11345 14059
rect 10928 14028 11345 14056
rect 10928 14016 10934 14028
rect 11333 14025 11345 14028
rect 11379 14025 11391 14059
rect 11333 14019 11391 14025
rect 12989 14059 13047 14065
rect 12989 14025 13001 14059
rect 13035 14056 13047 14059
rect 13078 14056 13084 14068
rect 13035 14028 13084 14056
rect 13035 14025 13047 14028
rect 12989 14019 13047 14025
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 13265 14059 13323 14065
rect 13265 14025 13277 14059
rect 13311 14056 13323 14059
rect 15010 14056 15016 14068
rect 13311 14028 14872 14056
rect 14971 14028 15016 14056
rect 13311 14025 13323 14028
rect 13265 14019 13323 14025
rect 10612 13960 11100 13988
rect 10505 13951 10563 13957
rect 9309 13923 9367 13929
rect 9309 13889 9321 13923
rect 9355 13889 9367 13923
rect 9309 13883 9367 13889
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13920 9551 13923
rect 9582 13920 9588 13932
rect 9539 13892 9588 13920
rect 9539 13889 9551 13892
rect 9493 13883 9551 13889
rect 9582 13880 9588 13892
rect 9640 13880 9646 13932
rect 10134 13920 10140 13932
rect 10095 13892 10140 13920
rect 10134 13880 10140 13892
rect 10192 13880 10198 13932
rect 10226 13880 10232 13932
rect 10284 13920 10290 13932
rect 10962 13920 10968 13932
rect 10284 13892 10329 13920
rect 10923 13892 10968 13920
rect 10284 13880 10290 13892
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 11072 13929 11100 13960
rect 14550 13948 14556 14000
rect 14608 13988 14614 14000
rect 14737 13991 14795 13997
rect 14737 13988 14749 13991
rect 14608 13960 14749 13988
rect 14608 13948 14614 13960
rect 14737 13957 14749 13960
rect 14783 13957 14795 13991
rect 14844 13988 14872 14028
rect 15010 14016 15016 14028
rect 15068 14016 15074 14068
rect 15102 14016 15108 14068
rect 15160 14056 15166 14068
rect 17862 14056 17868 14068
rect 15160 14028 17868 14056
rect 15160 14016 15166 14028
rect 17862 14016 17868 14028
rect 17920 14016 17926 14068
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 19242 14056 19248 14068
rect 18012 14028 19248 14056
rect 18012 14016 18018 14028
rect 14844 13960 18000 13988
rect 14737 13951 14795 13957
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13889 11115 13923
rect 11057 13883 11115 13889
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13889 11943 13923
rect 11885 13883 11943 13889
rect 1670 13852 1676 13864
rect 1631 13824 1676 13852
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 2406 13852 2412 13864
rect 2367 13824 2412 13852
rect 2406 13812 2412 13824
rect 2464 13812 2470 13864
rect 2958 13852 2964 13864
rect 2919 13824 2964 13852
rect 2958 13812 2964 13824
rect 3016 13812 3022 13864
rect 3697 13855 3755 13861
rect 3697 13821 3709 13855
rect 3743 13852 3755 13855
rect 4246 13852 4252 13864
rect 3743 13824 4252 13852
rect 3743 13821 3755 13824
rect 3697 13815 3755 13821
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13852 5871 13855
rect 6822 13852 6828 13864
rect 5859 13824 6828 13852
rect 5859 13821 5871 13824
rect 5813 13815 5871 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7282 13852 7288 13864
rect 7243 13824 7288 13852
rect 7282 13812 7288 13824
rect 7340 13812 7346 13864
rect 7558 13861 7564 13864
rect 7552 13852 7564 13861
rect 7471 13824 7564 13852
rect 7552 13815 7564 13824
rect 7616 13852 7622 13864
rect 8938 13852 8944 13864
rect 7616 13824 8944 13852
rect 7558 13812 7564 13815
rect 7616 13812 7622 13824
rect 8938 13812 8944 13824
rect 8996 13852 9002 13864
rect 10244 13852 10272 13880
rect 8996 13824 10272 13852
rect 8996 13812 9002 13824
rect 10318 13812 10324 13864
rect 10376 13852 10382 13864
rect 11900 13852 11928 13883
rect 12250 13880 12256 13932
rect 12308 13920 12314 13932
rect 13357 13923 13415 13929
rect 13357 13920 13369 13923
rect 12308 13892 13369 13920
rect 12308 13880 12314 13892
rect 13357 13889 13369 13892
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 13630 13861 13636 13864
rect 10376 13824 11928 13852
rect 12805 13855 12863 13861
rect 10376 13812 10382 13824
rect 12805 13821 12817 13855
rect 12851 13852 12863 13855
rect 13265 13855 13323 13861
rect 13265 13852 13277 13855
rect 12851 13824 13277 13852
rect 12851 13821 12863 13824
rect 12805 13815 12863 13821
rect 13265 13821 13277 13824
rect 13311 13821 13323 13855
rect 13624 13852 13636 13861
rect 13543 13824 13636 13852
rect 13265 13815 13323 13821
rect 13624 13815 13636 13824
rect 13688 13852 13694 13864
rect 15580 13852 15608 13883
rect 16390 13880 16396 13932
rect 16448 13920 16454 13932
rect 16577 13923 16635 13929
rect 16577 13920 16589 13923
rect 16448 13892 16589 13920
rect 16448 13880 16454 13892
rect 16577 13889 16589 13892
rect 16623 13889 16635 13923
rect 17494 13920 17500 13932
rect 17455 13892 17500 13920
rect 16577 13883 16635 13889
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 13688 13824 15608 13852
rect 13630 13812 13636 13815
rect 13688 13812 13694 13824
rect 16298 13812 16304 13864
rect 16356 13812 16362 13864
rect 16485 13855 16543 13861
rect 16485 13821 16497 13855
rect 16531 13852 16543 13855
rect 17126 13852 17132 13864
rect 16531 13824 17132 13852
rect 16531 13821 16543 13824
rect 16485 13815 16543 13821
rect 17126 13812 17132 13824
rect 17184 13812 17190 13864
rect 17218 13812 17224 13864
rect 17276 13852 17282 13864
rect 17276 13824 17321 13852
rect 17276 13812 17282 13824
rect 3970 13793 3976 13796
rect 3964 13784 3976 13793
rect 3883 13756 3976 13784
rect 3964 13747 3976 13756
rect 4028 13784 4034 13796
rect 5534 13784 5540 13796
rect 4028 13756 5540 13784
rect 3970 13744 3976 13747
rect 4028 13744 4034 13756
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 8846 13744 8852 13796
rect 8904 13784 8910 13796
rect 9582 13784 9588 13796
rect 8904 13756 9588 13784
rect 8904 13744 8910 13756
rect 9582 13744 9588 13756
rect 9640 13744 9646 13796
rect 10873 13787 10931 13793
rect 10873 13784 10885 13787
rect 9692 13756 10885 13784
rect 5721 13719 5779 13725
rect 5721 13685 5733 13719
rect 5767 13716 5779 13719
rect 7742 13716 7748 13728
rect 5767 13688 7748 13716
rect 5767 13685 5779 13688
rect 5721 13679 5779 13685
rect 7742 13676 7748 13688
rect 7800 13676 7806 13728
rect 9214 13716 9220 13728
rect 9175 13688 9220 13716
rect 9214 13676 9220 13688
rect 9272 13676 9278 13728
rect 9692 13725 9720 13756
rect 10873 13753 10885 13756
rect 10919 13753 10931 13787
rect 10873 13747 10931 13753
rect 11701 13787 11759 13793
rect 11701 13753 11713 13787
rect 11747 13784 11759 13787
rect 14366 13784 14372 13796
rect 11747 13756 14372 13784
rect 11747 13753 11759 13756
rect 11701 13747 11759 13753
rect 14366 13744 14372 13756
rect 14424 13744 14430 13796
rect 15010 13744 15016 13796
rect 15068 13784 15074 13796
rect 15930 13784 15936 13796
rect 15068 13756 15936 13784
rect 15068 13744 15074 13756
rect 15930 13744 15936 13756
rect 15988 13744 15994 13796
rect 16316 13784 16344 13812
rect 17862 13784 17868 13796
rect 16316 13756 17868 13784
rect 17862 13744 17868 13756
rect 17920 13744 17926 13796
rect 17972 13784 18000 13960
rect 18064 13861 18092 14028
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 18230 13988 18236 14000
rect 18191 13960 18236 13988
rect 18230 13948 18236 13960
rect 18288 13948 18294 14000
rect 19702 13880 19708 13932
rect 19760 13920 19766 13932
rect 20809 13923 20867 13929
rect 20809 13920 20821 13923
rect 19760 13892 20821 13920
rect 19760 13880 19766 13892
rect 20809 13889 20821 13892
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18509 13855 18567 13861
rect 18509 13821 18521 13855
rect 18555 13852 18567 13855
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18555 13824 18613 13852
rect 18555 13821 18567 13824
rect 18509 13815 18567 13821
rect 18601 13821 18613 13824
rect 18647 13821 18659 13855
rect 18601 13815 18659 13821
rect 18868 13855 18926 13861
rect 18868 13821 18880 13855
rect 18914 13852 18926 13855
rect 19426 13852 19432 13864
rect 18914 13824 19432 13852
rect 18914 13821 18926 13824
rect 18868 13815 18926 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 20438 13812 20444 13864
rect 20496 13852 20502 13864
rect 20717 13855 20775 13861
rect 20717 13852 20729 13855
rect 20496 13824 20729 13852
rect 20496 13812 20502 13824
rect 20717 13821 20729 13824
rect 20763 13821 20775 13855
rect 20717 13815 20775 13821
rect 17972 13756 18644 13784
rect 18616 13728 18644 13756
rect 9677 13719 9735 13725
rect 9677 13685 9689 13719
rect 9723 13685 9735 13719
rect 9677 13679 9735 13685
rect 10045 13719 10103 13725
rect 10045 13685 10057 13719
rect 10091 13716 10103 13719
rect 10134 13716 10140 13728
rect 10091 13688 10140 13716
rect 10091 13685 10103 13688
rect 10045 13679 10103 13685
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 10502 13676 10508 13728
rect 10560 13716 10566 13728
rect 10778 13716 10784 13728
rect 10560 13688 10784 13716
rect 10560 13676 10566 13688
rect 10778 13676 10784 13688
rect 10836 13676 10842 13728
rect 11790 13716 11796 13728
rect 11751 13688 11796 13716
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 12894 13676 12900 13728
rect 12952 13716 12958 13728
rect 15194 13716 15200 13728
rect 12952 13688 15200 13716
rect 12952 13676 12958 13688
rect 15194 13676 15200 13688
rect 15252 13676 15258 13728
rect 15286 13676 15292 13728
rect 15344 13716 15350 13728
rect 15381 13719 15439 13725
rect 15381 13716 15393 13719
rect 15344 13688 15393 13716
rect 15344 13676 15350 13688
rect 15381 13685 15393 13688
rect 15427 13685 15439 13719
rect 15381 13679 15439 13685
rect 15473 13719 15531 13725
rect 15473 13685 15485 13719
rect 15519 13716 15531 13719
rect 16025 13719 16083 13725
rect 16025 13716 16037 13719
rect 15519 13688 16037 13716
rect 15519 13685 15531 13688
rect 15473 13679 15531 13685
rect 16025 13685 16037 13688
rect 16071 13685 16083 13719
rect 16025 13679 16083 13685
rect 16298 13676 16304 13728
rect 16356 13716 16362 13728
rect 16393 13719 16451 13725
rect 16393 13716 16405 13719
rect 16356 13688 16405 13716
rect 16356 13676 16362 13688
rect 16393 13685 16405 13688
rect 16439 13716 16451 13719
rect 16482 13716 16488 13728
rect 16439 13688 16488 13716
rect 16439 13685 16451 13688
rect 16393 13679 16451 13685
rect 16482 13676 16488 13688
rect 16540 13676 16546 13728
rect 17770 13676 17776 13728
rect 17828 13716 17834 13728
rect 18509 13719 18567 13725
rect 18509 13716 18521 13719
rect 17828 13688 18521 13716
rect 17828 13676 17834 13688
rect 18509 13685 18521 13688
rect 18555 13685 18567 13719
rect 18509 13679 18567 13685
rect 18598 13676 18604 13728
rect 18656 13676 18662 13728
rect 18966 13676 18972 13728
rect 19024 13716 19030 13728
rect 19242 13716 19248 13728
rect 19024 13688 19248 13716
rect 19024 13676 19030 13688
rect 19242 13676 19248 13688
rect 19300 13676 19306 13728
rect 19886 13676 19892 13728
rect 19944 13716 19950 13728
rect 19981 13719 20039 13725
rect 19981 13716 19993 13719
rect 19944 13688 19993 13716
rect 19944 13676 19950 13688
rect 19981 13685 19993 13688
rect 20027 13685 20039 13719
rect 20254 13716 20260 13728
rect 20215 13688 20260 13716
rect 19981 13679 20039 13685
rect 20254 13676 20260 13688
rect 20312 13676 20318 13728
rect 20625 13719 20683 13725
rect 20625 13685 20637 13719
rect 20671 13716 20683 13719
rect 20714 13716 20720 13728
rect 20671 13688 20720 13716
rect 20671 13685 20683 13688
rect 20625 13679 20683 13685
rect 20714 13676 20720 13688
rect 20772 13676 20778 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 1762 13512 1768 13524
rect 1723 13484 1768 13512
rect 1762 13472 1768 13484
rect 1820 13472 1826 13524
rect 4433 13515 4491 13521
rect 4433 13481 4445 13515
rect 4479 13512 4491 13515
rect 5813 13515 5871 13521
rect 5813 13512 5825 13515
rect 4479 13484 5825 13512
rect 4479 13481 4491 13484
rect 4433 13475 4491 13481
rect 5813 13481 5825 13484
rect 5859 13481 5871 13515
rect 5813 13475 5871 13481
rect 6086 13472 6092 13524
rect 6144 13512 6150 13524
rect 6917 13515 6975 13521
rect 6917 13512 6929 13515
rect 6144 13484 6929 13512
rect 6144 13472 6150 13484
rect 6917 13481 6929 13484
rect 6963 13512 6975 13515
rect 9398 13512 9404 13524
rect 6963 13484 9404 13512
rect 6963 13481 6975 13484
rect 6917 13475 6975 13481
rect 9398 13472 9404 13484
rect 9456 13472 9462 13524
rect 9858 13472 9864 13524
rect 9916 13512 9922 13524
rect 11425 13515 11483 13521
rect 11425 13512 11437 13515
rect 9916 13484 11437 13512
rect 9916 13472 9922 13484
rect 11425 13481 11437 13484
rect 11471 13481 11483 13515
rect 12986 13512 12992 13524
rect 12947 13484 12992 13512
rect 11425 13475 11483 13481
rect 2409 13447 2467 13453
rect 2409 13413 2421 13447
rect 2455 13444 2467 13447
rect 2958 13444 2964 13456
rect 2455 13416 2964 13444
rect 2455 13413 2467 13416
rect 2409 13407 2467 13413
rect 2958 13404 2964 13416
rect 3016 13404 3022 13456
rect 4706 13404 4712 13456
rect 4764 13444 4770 13456
rect 5350 13444 5356 13456
rect 4764 13416 5356 13444
rect 4764 13404 4770 13416
rect 5350 13404 5356 13416
rect 5408 13404 5414 13456
rect 6638 13404 6644 13456
rect 6696 13444 6702 13456
rect 7736 13447 7794 13453
rect 6696 13416 7696 13444
rect 6696 13404 6702 13416
rect 1578 13376 1584 13388
rect 1539 13348 1584 13376
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 2133 13379 2191 13385
rect 2133 13345 2145 13379
rect 2179 13376 2191 13379
rect 4154 13376 4160 13388
rect 2179 13348 4160 13376
rect 2179 13345 2191 13348
rect 2133 13339 2191 13345
rect 4154 13336 4160 13348
rect 4212 13336 4218 13388
rect 4246 13336 4252 13388
rect 4304 13376 4310 13388
rect 4801 13379 4859 13385
rect 4801 13376 4813 13379
rect 4304 13348 4813 13376
rect 4304 13336 4310 13348
rect 4801 13345 4813 13348
rect 4847 13345 4859 13379
rect 4801 13339 4859 13345
rect 6270 13336 6276 13388
rect 6328 13376 6334 13388
rect 6825 13379 6883 13385
rect 6825 13376 6837 13379
rect 6328 13348 6837 13376
rect 6328 13336 6334 13348
rect 6825 13345 6837 13348
rect 6871 13345 6883 13379
rect 7558 13376 7564 13388
rect 6825 13339 6883 13345
rect 7116 13348 7564 13376
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 4893 13311 4951 13317
rect 4893 13308 4905 13311
rect 4764 13280 4905 13308
rect 4764 13268 4770 13280
rect 4893 13277 4905 13280
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 5077 13311 5135 13317
rect 5077 13277 5089 13311
rect 5123 13308 5135 13311
rect 5534 13308 5540 13320
rect 5123 13280 5540 13308
rect 5123 13277 5135 13280
rect 5077 13271 5135 13277
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 5902 13308 5908 13320
rect 5863 13280 5908 13308
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 5994 13268 6000 13320
rect 6052 13308 6058 13320
rect 7116 13317 7144 13348
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 7668 13376 7696 13416
rect 7736 13413 7748 13447
rect 7782 13444 7794 13447
rect 8662 13444 8668 13456
rect 7782 13416 8668 13444
rect 7782 13413 7794 13416
rect 7736 13407 7794 13413
rect 8662 13404 8668 13416
rect 8720 13404 8726 13456
rect 10134 13376 10140 13388
rect 7668 13348 10140 13376
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 10312 13379 10370 13385
rect 10312 13345 10324 13379
rect 10358 13376 10370 13379
rect 11330 13376 11336 13388
rect 10358 13348 11336 13376
rect 10358 13345 10370 13348
rect 10312 13339 10370 13345
rect 11330 13336 11336 13348
rect 11388 13336 11394 13388
rect 11440 13376 11468 13475
rect 12986 13472 12992 13484
rect 13044 13472 13050 13524
rect 13170 13472 13176 13524
rect 13228 13512 13234 13524
rect 13449 13515 13507 13521
rect 13449 13512 13461 13515
rect 13228 13484 13461 13512
rect 13228 13472 13234 13484
rect 13449 13481 13461 13484
rect 13495 13481 13507 13515
rect 15286 13512 15292 13524
rect 15247 13484 15292 13512
rect 13449 13475 13507 13481
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 15746 13512 15752 13524
rect 15659 13484 15752 13512
rect 15746 13472 15752 13484
rect 15804 13512 15810 13524
rect 16022 13512 16028 13524
rect 15804 13484 16028 13512
rect 15804 13472 15810 13484
rect 16022 13472 16028 13484
rect 16080 13472 16086 13524
rect 16209 13515 16267 13521
rect 16209 13481 16221 13515
rect 16255 13512 16267 13515
rect 16390 13512 16396 13524
rect 16255 13484 16396 13512
rect 16255 13481 16267 13484
rect 16209 13475 16267 13481
rect 16390 13472 16396 13484
rect 16448 13512 16454 13524
rect 17681 13515 17739 13521
rect 17681 13512 17693 13515
rect 16448 13484 17693 13512
rect 16448 13472 16454 13484
rect 17681 13481 17693 13484
rect 17727 13481 17739 13515
rect 17681 13475 17739 13481
rect 19613 13515 19671 13521
rect 19613 13481 19625 13515
rect 19659 13512 19671 13515
rect 20530 13512 20536 13524
rect 19659 13484 20536 13512
rect 19659 13481 19671 13484
rect 19613 13475 19671 13481
rect 20530 13472 20536 13484
rect 20588 13472 20594 13524
rect 14185 13447 14243 13453
rect 14185 13413 14197 13447
rect 14231 13444 14243 13447
rect 15194 13444 15200 13456
rect 14231 13416 15200 13444
rect 14231 13413 14243 13416
rect 14185 13407 14243 13413
rect 15194 13404 15200 13416
rect 15252 13404 15258 13456
rect 16568 13447 16626 13453
rect 15856 13416 16344 13444
rect 11773 13379 11831 13385
rect 11773 13376 11785 13379
rect 11440 13348 11785 13376
rect 11773 13345 11785 13348
rect 11819 13345 11831 13379
rect 11773 13339 11831 13345
rect 12710 13336 12716 13388
rect 12768 13376 12774 13388
rect 13357 13379 13415 13385
rect 13357 13376 13369 13379
rect 12768 13348 13369 13376
rect 12768 13336 12774 13348
rect 13357 13345 13369 13348
rect 13403 13345 13415 13379
rect 13357 13339 13415 13345
rect 14277 13379 14335 13385
rect 14277 13345 14289 13379
rect 14323 13376 14335 13379
rect 14645 13379 14703 13385
rect 14323 13348 14596 13376
rect 14323 13345 14335 13348
rect 14277 13339 14335 13345
rect 14568 13320 14596 13348
rect 14645 13345 14657 13379
rect 14691 13345 14703 13379
rect 14645 13339 14703 13345
rect 7101 13311 7159 13317
rect 6052 13280 6097 13308
rect 6052 13268 6058 13280
rect 7101 13277 7113 13311
rect 7147 13277 7159 13311
rect 7101 13271 7159 13277
rect 7282 13268 7288 13320
rect 7340 13308 7346 13320
rect 7469 13311 7527 13317
rect 7469 13308 7481 13311
rect 7340 13280 7481 13308
rect 7340 13268 7346 13280
rect 7469 13277 7481 13280
rect 7515 13277 7527 13311
rect 7469 13271 7527 13277
rect 9122 13268 9128 13320
rect 9180 13308 9186 13320
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 9180 13280 10057 13308
rect 9180 13268 9186 13280
rect 10045 13277 10057 13280
rect 10091 13277 10103 13311
rect 10045 13271 10103 13277
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 4798 13200 4804 13252
rect 4856 13240 4862 13252
rect 5445 13243 5503 13249
rect 5445 13240 5457 13243
rect 4856 13212 5457 13240
rect 4856 13200 4862 13212
rect 5445 13209 5457 13212
rect 5491 13209 5503 13243
rect 8846 13240 8852 13252
rect 8807 13212 8852 13240
rect 5445 13203 5503 13209
rect 8846 13200 8852 13212
rect 8904 13200 8910 13252
rect 6457 13175 6515 13181
rect 6457 13141 6469 13175
rect 6503 13172 6515 13175
rect 7650 13172 7656 13184
rect 6503 13144 7656 13172
rect 6503 13141 6515 13144
rect 6457 13135 6515 13141
rect 7650 13132 7656 13144
rect 7708 13132 7714 13184
rect 11532 13172 11560 13271
rect 12526 13268 12532 13320
rect 12584 13308 12590 13320
rect 13633 13311 13691 13317
rect 13633 13308 13645 13311
rect 12584 13280 13645 13308
rect 12584 13268 12590 13280
rect 13633 13277 13645 13280
rect 13679 13277 13691 13311
rect 14458 13308 14464 13320
rect 14419 13280 14464 13308
rect 13633 13271 13691 13277
rect 12894 13240 12900 13252
rect 12855 13212 12900 13240
rect 12894 13200 12900 13212
rect 12952 13200 12958 13252
rect 13648 13240 13676 13271
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 14550 13268 14556 13320
rect 14608 13268 14614 13320
rect 14660 13308 14688 13339
rect 15010 13336 15016 13388
rect 15068 13376 15074 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 15068 13348 15669 13376
rect 15068 13336 15074 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 15856 13308 15884 13416
rect 16209 13379 16267 13385
rect 16209 13376 16221 13379
rect 15948 13348 16221 13376
rect 15948 13317 15976 13348
rect 16209 13345 16221 13348
rect 16255 13345 16267 13379
rect 16316 13376 16344 13416
rect 16568 13413 16580 13447
rect 16614 13444 16626 13447
rect 19886 13444 19892 13456
rect 16614 13416 19892 13444
rect 16614 13413 16626 13416
rect 16568 13407 16626 13413
rect 19886 13404 19892 13416
rect 19944 13444 19950 13456
rect 19944 13416 20208 13444
rect 19944 13404 19950 13416
rect 16316 13348 17724 13376
rect 16209 13339 16267 13345
rect 14660 13280 15884 13308
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13277 15991 13311
rect 15933 13271 15991 13277
rect 15948 13240 15976 13271
rect 16114 13268 16120 13320
rect 16172 13308 16178 13320
rect 16301 13311 16359 13317
rect 16301 13308 16313 13311
rect 16172 13280 16313 13308
rect 16172 13268 16178 13280
rect 16301 13277 16313 13280
rect 16347 13277 16359 13311
rect 16301 13271 16359 13277
rect 13648 13212 15976 13240
rect 12250 13172 12256 13184
rect 11532 13144 12256 13172
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 13817 13175 13875 13181
rect 13817 13172 13829 13175
rect 13780 13144 13829 13172
rect 13780 13132 13786 13144
rect 13817 13141 13829 13144
rect 13863 13141 13875 13175
rect 13817 13135 13875 13141
rect 13906 13132 13912 13184
rect 13964 13172 13970 13184
rect 14274 13172 14280 13184
rect 13964 13144 14280 13172
rect 13964 13132 13970 13144
rect 14274 13132 14280 13144
rect 14332 13132 14338 13184
rect 14829 13175 14887 13181
rect 14829 13141 14841 13175
rect 14875 13172 14887 13175
rect 14918 13172 14924 13184
rect 14875 13144 14924 13172
rect 14875 13141 14887 13144
rect 14829 13135 14887 13141
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 17696 13172 17724 13348
rect 17770 13336 17776 13388
rect 17828 13376 17834 13388
rect 18230 13385 18236 13388
rect 17957 13379 18015 13385
rect 17957 13376 17969 13379
rect 17828 13348 17969 13376
rect 17828 13336 17834 13348
rect 17957 13345 17969 13348
rect 18003 13345 18015 13379
rect 18224 13376 18236 13385
rect 18191 13348 18236 13376
rect 17957 13339 18015 13345
rect 18224 13339 18236 13348
rect 18288 13376 18294 13388
rect 19521 13379 19579 13385
rect 19521 13376 19533 13379
rect 18288 13348 19533 13376
rect 18230 13336 18236 13339
rect 18288 13336 18294 13348
rect 19521 13345 19533 13348
rect 19567 13345 19579 13379
rect 19521 13339 19579 13345
rect 19610 13336 19616 13388
rect 19668 13376 19674 13388
rect 19981 13379 20039 13385
rect 19981 13376 19993 13379
rect 19668 13348 19993 13376
rect 19668 13336 19674 13348
rect 19981 13345 19993 13348
rect 20027 13345 20039 13379
rect 19981 13339 20039 13345
rect 18966 13268 18972 13320
rect 19024 13308 19030 13320
rect 20180 13317 20208 13416
rect 20073 13311 20131 13317
rect 20073 13308 20085 13311
rect 19024 13280 20085 13308
rect 19024 13268 19030 13280
rect 20073 13277 20085 13280
rect 20119 13277 20131 13311
rect 20073 13271 20131 13277
rect 20165 13311 20223 13317
rect 20165 13277 20177 13311
rect 20211 13277 20223 13311
rect 20165 13271 20223 13277
rect 20806 13240 20812 13252
rect 18892 13212 20812 13240
rect 18892 13172 18920 13212
rect 20806 13200 20812 13212
rect 20864 13200 20870 13252
rect 17696 13144 18920 13172
rect 19337 13175 19395 13181
rect 19337 13141 19349 13175
rect 19383 13172 19395 13175
rect 19426 13172 19432 13184
rect 19383 13144 19432 13172
rect 19383 13141 19395 13144
rect 19337 13135 19395 13141
rect 19426 13132 19432 13144
rect 19484 13132 19490 13184
rect 19521 13175 19579 13181
rect 19521 13141 19533 13175
rect 19567 13172 19579 13175
rect 19702 13172 19708 13184
rect 19567 13144 19708 13172
rect 19567 13141 19579 13144
rect 19521 13135 19579 13141
rect 19702 13132 19708 13144
rect 19760 13172 19766 13184
rect 20530 13172 20536 13184
rect 19760 13144 20536 13172
rect 19760 13132 19766 13144
rect 20530 13132 20536 13144
rect 20588 13132 20594 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1489 12971 1547 12977
rect 1489 12937 1501 12971
rect 1535 12968 1547 12971
rect 1670 12968 1676 12980
rect 1535 12940 1676 12968
rect 1535 12937 1547 12940
rect 1489 12931 1547 12937
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 3881 12971 3939 12977
rect 3881 12937 3893 12971
rect 3927 12968 3939 12971
rect 3970 12968 3976 12980
rect 3927 12940 3976 12968
rect 3927 12937 3939 12940
rect 3881 12931 3939 12937
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 4709 12971 4767 12977
rect 4709 12937 4721 12971
rect 4755 12968 4767 12971
rect 5902 12968 5908 12980
rect 4755 12940 5908 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 5902 12928 5908 12940
rect 5960 12928 5966 12980
rect 7193 12971 7251 12977
rect 7193 12937 7205 12971
rect 7239 12968 7251 12971
rect 9214 12968 9220 12980
rect 7239 12940 9220 12968
rect 7239 12937 7251 12940
rect 7193 12931 7251 12937
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 10870 12968 10876 12980
rect 9732 12940 10876 12968
rect 9732 12928 9738 12940
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 12713 12971 12771 12977
rect 12713 12937 12725 12971
rect 12759 12968 12771 12971
rect 13998 12968 14004 12980
rect 12759 12940 14004 12968
rect 12759 12937 12771 12940
rect 12713 12931 12771 12937
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 17218 12968 17224 12980
rect 14292 12940 17224 12968
rect 3510 12860 3516 12912
rect 3568 12900 3574 12912
rect 13170 12900 13176 12912
rect 3568 12872 13176 12900
rect 3568 12860 3574 12872
rect 13170 12860 13176 12872
rect 13228 12860 13234 12912
rect 13265 12903 13323 12909
rect 13265 12869 13277 12903
rect 13311 12900 13323 12903
rect 14292 12900 14320 12940
rect 17218 12928 17224 12940
rect 17276 12928 17282 12980
rect 18966 12968 18972 12980
rect 18927 12940 18972 12968
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 13311 12872 14320 12900
rect 15657 12903 15715 12909
rect 13311 12869 13323 12872
rect 13265 12863 13323 12869
rect 15657 12869 15669 12903
rect 15703 12869 15715 12903
rect 15657 12863 15715 12869
rect 2133 12835 2191 12841
rect 2133 12801 2145 12835
rect 2179 12832 2191 12835
rect 4246 12832 4252 12844
rect 2179 12804 2636 12832
rect 4207 12804 4252 12832
rect 2179 12801 2191 12804
rect 2133 12795 2191 12801
rect 1486 12724 1492 12776
rect 1544 12764 1550 12776
rect 2501 12767 2559 12773
rect 2501 12764 2513 12767
rect 1544 12736 2513 12764
rect 1544 12724 1550 12736
rect 2501 12733 2513 12736
rect 2547 12733 2559 12767
rect 2608 12764 2636 12804
rect 4246 12792 4252 12804
rect 4304 12792 4310 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5534 12832 5540 12844
rect 5399 12804 5540 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 6178 12832 6184 12844
rect 6139 12804 6184 12832
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 6362 12832 6368 12844
rect 6323 12804 6368 12832
rect 6362 12792 6368 12804
rect 6420 12792 6426 12844
rect 7650 12832 7656 12844
rect 7611 12804 7656 12832
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 7837 12835 7895 12841
rect 7837 12801 7849 12835
rect 7883 12832 7895 12835
rect 8662 12832 8668 12844
rect 7883 12804 8668 12832
rect 7883 12801 7895 12804
rect 7837 12795 7895 12801
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 8849 12835 8907 12841
rect 8849 12801 8861 12835
rect 8895 12832 8907 12835
rect 8938 12832 8944 12844
rect 8895 12804 8944 12832
rect 8895 12801 8907 12804
rect 8849 12795 8907 12801
rect 8938 12792 8944 12804
rect 8996 12792 9002 12844
rect 9398 12792 9404 12844
rect 9456 12832 9462 12844
rect 12250 12832 12256 12844
rect 9456 12804 12256 12832
rect 9456 12792 9462 12804
rect 12250 12792 12256 12804
rect 12308 12792 12314 12844
rect 13722 12832 13728 12844
rect 13683 12804 13728 12832
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 13817 12835 13875 12841
rect 13817 12801 13829 12835
rect 13863 12801 13875 12835
rect 13817 12795 13875 12801
rect 2774 12773 2780 12776
rect 2757 12767 2780 12773
rect 2757 12764 2769 12767
rect 2608 12736 2769 12764
rect 2501 12727 2559 12733
rect 2757 12733 2769 12736
rect 2832 12764 2838 12776
rect 2832 12736 2905 12764
rect 2757 12727 2780 12733
rect 2774 12724 2780 12727
rect 2832 12724 2838 12736
rect 4890 12724 4896 12776
rect 4948 12764 4954 12776
rect 9861 12767 9919 12773
rect 4948 12736 8340 12764
rect 4948 12724 4954 12736
rect 5169 12699 5227 12705
rect 5169 12665 5181 12699
rect 5215 12696 5227 12699
rect 5350 12696 5356 12708
rect 5215 12668 5356 12696
rect 5215 12665 5227 12668
rect 5169 12659 5227 12665
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 7561 12699 7619 12705
rect 7561 12665 7573 12699
rect 7607 12696 7619 12699
rect 7607 12668 8248 12696
rect 7607 12665 7619 12668
rect 7561 12659 7619 12665
rect 1854 12628 1860 12640
rect 1815 12600 1860 12628
rect 1854 12588 1860 12600
rect 1912 12588 1918 12640
rect 1946 12588 1952 12640
rect 2004 12628 2010 12640
rect 5074 12628 5080 12640
rect 2004 12600 2049 12628
rect 5035 12600 5080 12628
rect 2004 12588 2010 12600
rect 5074 12588 5080 12600
rect 5132 12588 5138 12640
rect 5721 12631 5779 12637
rect 5721 12597 5733 12631
rect 5767 12628 5779 12631
rect 5994 12628 6000 12640
rect 5767 12600 6000 12628
rect 5767 12597 5779 12600
rect 5721 12591 5779 12597
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 6086 12588 6092 12640
rect 6144 12628 6150 12640
rect 8220 12637 8248 12668
rect 8205 12631 8263 12637
rect 6144 12600 6189 12628
rect 6144 12588 6150 12600
rect 8205 12597 8217 12631
rect 8251 12597 8263 12631
rect 8312 12628 8340 12736
rect 9861 12733 9873 12767
rect 9907 12764 9919 12767
rect 11977 12767 12035 12773
rect 11977 12764 11989 12767
rect 9907 12736 11989 12764
rect 9907 12733 9919 12736
rect 9861 12727 9919 12733
rect 11977 12733 11989 12736
rect 12023 12764 12035 12767
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12023 12736 12909 12764
rect 12023 12733 12035 12736
rect 11977 12727 12035 12733
rect 12897 12733 12909 12736
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 13630 12724 13636 12776
rect 13688 12764 13694 12776
rect 13832 12764 13860 12795
rect 15378 12792 15384 12844
rect 15436 12832 15442 12844
rect 15672 12832 15700 12863
rect 15838 12860 15844 12912
rect 15896 12900 15902 12912
rect 17954 12900 17960 12912
rect 15896 12872 17960 12900
rect 15896 12860 15902 12872
rect 17954 12860 17960 12872
rect 18012 12860 18018 12912
rect 18046 12860 18052 12912
rect 18104 12900 18110 12912
rect 18874 12900 18880 12912
rect 18104 12872 18880 12900
rect 18104 12860 18110 12872
rect 18874 12860 18880 12872
rect 18932 12860 18938 12912
rect 19058 12860 19064 12912
rect 19116 12900 19122 12912
rect 20346 12900 20352 12912
rect 19116 12872 20352 12900
rect 19116 12860 19122 12872
rect 20346 12860 20352 12872
rect 20404 12900 20410 12912
rect 21082 12900 21088 12912
rect 20404 12872 21088 12900
rect 20404 12860 20410 12872
rect 21082 12860 21088 12872
rect 21140 12860 21146 12912
rect 16485 12835 16543 12841
rect 16485 12832 16497 12835
rect 15436 12804 16497 12832
rect 15436 12792 15442 12804
rect 16485 12801 16497 12804
rect 16531 12801 16543 12835
rect 16485 12795 16543 12801
rect 16574 12792 16580 12844
rect 16632 12832 16638 12844
rect 17034 12832 17040 12844
rect 16632 12804 17040 12832
rect 16632 12792 16638 12804
rect 17034 12792 17040 12804
rect 17092 12792 17098 12844
rect 17218 12792 17224 12844
rect 17276 12832 17282 12844
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 17276 12804 17417 12832
rect 17276 12792 17282 12804
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 17494 12792 17500 12844
rect 17552 12832 17558 12844
rect 18509 12835 18567 12841
rect 17552 12804 17597 12832
rect 17552 12792 17558 12804
rect 18509 12801 18521 12835
rect 18555 12832 18567 12835
rect 18598 12832 18604 12844
rect 18555 12804 18604 12832
rect 18555 12801 18567 12804
rect 18509 12795 18567 12801
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 19426 12792 19432 12844
rect 19484 12832 19490 12844
rect 19613 12835 19671 12841
rect 19613 12832 19625 12835
rect 19484 12804 19625 12832
rect 19484 12792 19490 12804
rect 19613 12801 19625 12804
rect 19659 12832 19671 12835
rect 20162 12832 20168 12844
rect 19659 12804 20168 12832
rect 19659 12801 19671 12804
rect 19613 12795 19671 12801
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 20530 12832 20536 12844
rect 20491 12804 20536 12832
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 13688 12736 13860 12764
rect 14277 12767 14335 12773
rect 13688 12724 13694 12736
rect 14277 12733 14289 12767
rect 14323 12733 14335 12767
rect 14277 12727 14335 12733
rect 14544 12767 14602 12773
rect 14544 12733 14556 12767
rect 14590 12764 14602 12767
rect 14826 12764 14832 12776
rect 14590 12736 14832 12764
rect 14590 12733 14602 12736
rect 14544 12727 14602 12733
rect 8573 12699 8631 12705
rect 8573 12665 8585 12699
rect 8619 12696 8631 12699
rect 9217 12699 9275 12705
rect 9217 12696 9229 12699
rect 8619 12668 9229 12696
rect 8619 12665 8631 12668
rect 8573 12659 8631 12665
rect 9217 12665 9229 12668
rect 9263 12665 9275 12699
rect 9217 12659 9275 12665
rect 10134 12656 10140 12708
rect 10192 12696 10198 12708
rect 10413 12699 10471 12705
rect 10413 12696 10425 12699
rect 10192 12668 10425 12696
rect 10192 12656 10198 12668
rect 10413 12665 10425 12668
rect 10459 12665 10471 12699
rect 14292 12696 14320 12727
rect 14826 12724 14832 12736
rect 14884 12724 14890 12776
rect 16114 12764 16120 12776
rect 15028 12736 16120 12764
rect 15028 12696 15056 12736
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 16390 12764 16396 12776
rect 16351 12736 16396 12764
rect 16390 12724 16396 12736
rect 16448 12724 16454 12776
rect 18233 12767 18291 12773
rect 18233 12764 18245 12767
rect 16960 12736 18245 12764
rect 14292 12668 15056 12696
rect 10413 12659 10471 12665
rect 15102 12656 15108 12708
rect 15160 12696 15166 12708
rect 16301 12699 16359 12705
rect 16301 12696 16313 12699
rect 15160 12668 16313 12696
rect 15160 12656 15166 12668
rect 16301 12665 16313 12668
rect 16347 12665 16359 12699
rect 16301 12659 16359 12665
rect 8665 12631 8723 12637
rect 8665 12628 8677 12631
rect 8312 12600 8677 12628
rect 8205 12591 8263 12597
rect 8665 12597 8677 12600
rect 8711 12597 8723 12631
rect 8665 12591 8723 12597
rect 8754 12588 8760 12640
rect 8812 12628 8818 12640
rect 9677 12631 9735 12637
rect 9677 12628 9689 12631
rect 8812 12600 9689 12628
rect 8812 12588 8818 12600
rect 9677 12597 9689 12600
rect 9723 12597 9735 12631
rect 9677 12591 9735 12597
rect 13633 12631 13691 12637
rect 13633 12597 13645 12631
rect 13679 12628 13691 12631
rect 13906 12628 13912 12640
rect 13679 12600 13912 12628
rect 13679 12597 13691 12600
rect 13633 12591 13691 12597
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 15930 12628 15936 12640
rect 15891 12600 15936 12628
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 16960 12637 16988 12736
rect 18233 12733 18245 12736
rect 18279 12733 18291 12767
rect 18233 12727 18291 12733
rect 19337 12767 19395 12773
rect 19337 12733 19349 12767
rect 19383 12764 19395 12767
rect 20254 12764 20260 12776
rect 19383 12736 20260 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 17310 12696 17316 12708
rect 17271 12668 17316 12696
rect 17310 12656 17316 12668
rect 17368 12656 17374 12708
rect 19429 12699 19487 12705
rect 19429 12665 19441 12699
rect 19475 12696 19487 12699
rect 19518 12696 19524 12708
rect 19475 12668 19524 12696
rect 19475 12665 19487 12668
rect 19429 12659 19487 12665
rect 19518 12656 19524 12668
rect 19576 12656 19582 12708
rect 20349 12699 20407 12705
rect 19628 12668 20116 12696
rect 16945 12631 17003 12637
rect 16945 12597 16957 12631
rect 16991 12597 17003 12631
rect 16945 12591 17003 12597
rect 17034 12588 17040 12640
rect 17092 12628 17098 12640
rect 19628 12628 19656 12668
rect 19978 12628 19984 12640
rect 17092 12600 19656 12628
rect 19939 12600 19984 12628
rect 17092 12588 17098 12600
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 20088 12628 20116 12668
rect 20349 12665 20361 12699
rect 20395 12696 20407 12699
rect 20898 12696 20904 12708
rect 20395 12668 20904 12696
rect 20395 12665 20407 12668
rect 20349 12659 20407 12665
rect 20898 12656 20904 12668
rect 20956 12656 20962 12708
rect 20441 12631 20499 12637
rect 20441 12628 20453 12631
rect 20088 12600 20453 12628
rect 20441 12597 20453 12600
rect 20487 12597 20499 12631
rect 20441 12591 20499 12597
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 2961 12427 3019 12433
rect 2961 12424 2973 12427
rect 2832 12396 2973 12424
rect 2832 12384 2838 12396
rect 2961 12393 2973 12396
rect 3007 12393 3019 12427
rect 2961 12387 3019 12393
rect 4246 12384 4252 12436
rect 4304 12424 4310 12436
rect 5997 12427 6055 12433
rect 5997 12424 6009 12427
rect 4304 12396 6009 12424
rect 4304 12384 4310 12396
rect 5997 12393 6009 12396
rect 6043 12393 6055 12427
rect 5997 12387 6055 12393
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 8202 12424 8208 12436
rect 7156 12396 8208 12424
rect 7156 12384 7162 12396
rect 8202 12384 8208 12396
rect 8260 12424 8266 12436
rect 8754 12424 8760 12436
rect 8260 12396 8760 12424
rect 8260 12384 8266 12396
rect 8754 12384 8760 12396
rect 8812 12384 8818 12436
rect 10318 12384 10324 12436
rect 10376 12424 10382 12436
rect 10686 12424 10692 12436
rect 10376 12396 10692 12424
rect 10376 12384 10382 12396
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 11057 12427 11115 12433
rect 11057 12393 11069 12427
rect 11103 12424 11115 12427
rect 12526 12424 12532 12436
rect 11103 12396 12532 12424
rect 11103 12393 11115 12396
rect 11057 12387 11115 12393
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 13688 12396 14289 12424
rect 13688 12384 13694 12396
rect 14277 12393 14289 12396
rect 14323 12393 14335 12427
rect 14277 12387 14335 12393
rect 14737 12427 14795 12433
rect 14737 12393 14749 12427
rect 14783 12424 14795 12427
rect 15010 12424 15016 12436
rect 14783 12396 15016 12424
rect 14783 12393 14795 12396
rect 14737 12387 14795 12393
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 15289 12427 15347 12433
rect 15289 12424 15301 12427
rect 15252 12396 15301 12424
rect 15252 12384 15258 12396
rect 15289 12393 15301 12396
rect 15335 12393 15347 12427
rect 15289 12387 15347 12393
rect 17494 12384 17500 12436
rect 17552 12424 17558 12436
rect 17865 12427 17923 12433
rect 17865 12424 17877 12427
rect 17552 12396 17877 12424
rect 17552 12384 17558 12396
rect 17865 12393 17877 12396
rect 17911 12393 17923 12427
rect 19610 12424 19616 12436
rect 19571 12396 19616 12424
rect 17865 12387 17923 12393
rect 19610 12384 19616 12396
rect 19668 12384 19674 12436
rect 19978 12424 19984 12436
rect 19939 12396 19984 12424
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 20898 12424 20904 12436
rect 20859 12396 20904 12424
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 15746 12356 15752 12368
rect 4120 12328 15752 12356
rect 4120 12316 4126 12328
rect 15746 12316 15752 12328
rect 15804 12316 15810 12368
rect 16752 12359 16810 12365
rect 16752 12325 16764 12359
rect 16798 12356 16810 12359
rect 17402 12356 17408 12368
rect 16798 12328 17408 12356
rect 16798 12325 16810 12328
rect 16752 12319 16810 12325
rect 17402 12316 17408 12328
rect 17460 12356 17466 12368
rect 17586 12356 17592 12368
rect 17460 12328 17592 12356
rect 17460 12316 17466 12328
rect 17586 12316 17592 12328
rect 17644 12316 17650 12368
rect 17770 12316 17776 12368
rect 17828 12356 17834 12368
rect 20438 12356 20444 12368
rect 17828 12328 20444 12356
rect 17828 12316 17834 12328
rect 20438 12316 20444 12328
rect 20496 12316 20502 12368
rect 1848 12291 1906 12297
rect 1848 12257 1860 12291
rect 1894 12288 1906 12291
rect 2682 12288 2688 12300
rect 1894 12260 2688 12288
rect 1894 12257 1906 12260
rect 1848 12251 1906 12257
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 4700 12291 4758 12297
rect 4700 12257 4712 12291
rect 4746 12288 4758 12291
rect 5258 12288 5264 12300
rect 4746 12260 5264 12288
rect 4746 12257 4758 12260
rect 4700 12251 4758 12257
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 6345 12291 6403 12297
rect 6345 12288 6357 12291
rect 5828 12260 6357 12288
rect 1486 12180 1492 12232
rect 1544 12220 1550 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 1544 12192 1593 12220
rect 1544 12180 1550 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 4246 12180 4252 12232
rect 4304 12220 4310 12232
rect 4433 12223 4491 12229
rect 4433 12220 4445 12223
rect 4304 12192 4445 12220
rect 4304 12180 4310 12192
rect 4433 12189 4445 12192
rect 4479 12189 4491 12223
rect 4433 12183 4491 12189
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 5828 12093 5856 12260
rect 6345 12257 6357 12260
rect 6391 12257 6403 12291
rect 8012 12291 8070 12297
rect 8012 12288 8024 12291
rect 6345 12251 6403 12257
rect 7668 12260 8024 12288
rect 5997 12223 6055 12229
rect 5997 12189 6009 12223
rect 6043 12220 6055 12223
rect 6089 12223 6147 12229
rect 6089 12220 6101 12223
rect 6043 12192 6101 12220
rect 6043 12189 6055 12192
rect 5997 12183 6055 12189
rect 6089 12189 6101 12192
rect 6135 12189 6147 12223
rect 6089 12183 6147 12189
rect 7469 12155 7527 12161
rect 7469 12121 7481 12155
rect 7515 12152 7527 12155
rect 7668 12152 7696 12260
rect 8012 12257 8024 12260
rect 8058 12288 8070 12291
rect 9214 12288 9220 12300
rect 8058 12260 9220 12288
rect 8058 12257 8070 12260
rect 8012 12251 8070 12257
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 10134 12248 10140 12300
rect 10192 12288 10198 12300
rect 10410 12288 10416 12300
rect 10192 12260 10416 12288
rect 10192 12248 10198 12260
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 10594 12288 10600 12300
rect 10555 12260 10600 12288
rect 10594 12248 10600 12260
rect 10652 12288 10658 12300
rect 10778 12288 10784 12300
rect 10652 12260 10784 12288
rect 10652 12248 10658 12260
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 11508 12291 11566 12297
rect 11508 12288 11520 12291
rect 10888 12260 11520 12288
rect 7742 12180 7748 12232
rect 7800 12220 7806 12232
rect 7800 12192 7845 12220
rect 7800 12180 7806 12192
rect 8754 12180 8760 12232
rect 8812 12220 8818 12232
rect 10686 12220 10692 12232
rect 8812 12192 10692 12220
rect 8812 12180 8818 12192
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 10888 12229 10916 12260
rect 11508 12257 11520 12260
rect 11554 12288 11566 12291
rect 12342 12288 12348 12300
rect 11554 12260 12348 12288
rect 11554 12257 11566 12260
rect 11508 12251 11566 12257
rect 12342 12248 12348 12260
rect 12400 12248 12406 12300
rect 13164 12291 13222 12297
rect 13164 12288 13176 12291
rect 12728 12260 13176 12288
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12189 10931 12223
rect 10873 12183 10931 12189
rect 11146 12180 11152 12232
rect 11204 12220 11210 12232
rect 11241 12223 11299 12229
rect 11241 12220 11253 12223
rect 11204 12192 11253 12220
rect 11204 12180 11210 12192
rect 11241 12189 11253 12192
rect 11287 12189 11299 12223
rect 11241 12183 11299 12189
rect 11057 12155 11115 12161
rect 11057 12152 11069 12155
rect 7515 12124 7696 12152
rect 8680 12124 11069 12152
rect 7515 12121 7527 12124
rect 7469 12115 7527 12121
rect 5813 12087 5871 12093
rect 5813 12084 5825 12087
rect 4856 12056 5825 12084
rect 4856 12044 4862 12056
rect 5813 12053 5825 12056
rect 5859 12053 5871 12087
rect 5813 12047 5871 12053
rect 5902 12044 5908 12096
rect 5960 12084 5966 12096
rect 8680 12084 8708 12124
rect 11057 12121 11069 12124
rect 11103 12121 11115 12155
rect 11057 12115 11115 12121
rect 12621 12155 12679 12161
rect 12621 12121 12633 12155
rect 12667 12152 12679 12155
rect 12728 12152 12756 12260
rect 13164 12257 13176 12260
rect 13210 12288 13222 12291
rect 14458 12288 14464 12300
rect 13210 12260 14464 12288
rect 13210 12257 13222 12260
rect 13164 12251 13222 12257
rect 14458 12248 14464 12260
rect 14516 12248 14522 12300
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12288 15715 12291
rect 17310 12288 17316 12300
rect 15703 12260 17316 12288
rect 15703 12257 15715 12260
rect 15657 12251 15715 12257
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 18969 12291 19027 12297
rect 18969 12257 18981 12291
rect 19015 12257 19027 12291
rect 20530 12288 20536 12300
rect 18969 12251 19027 12257
rect 19076 12260 20536 12288
rect 12894 12220 12900 12232
rect 12855 12192 12900 12220
rect 12894 12180 12900 12192
rect 12952 12180 12958 12232
rect 15746 12220 15752 12232
rect 15707 12192 15752 12220
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 12667 12124 12756 12152
rect 12667 12121 12679 12124
rect 12621 12115 12679 12121
rect 14458 12112 14464 12164
rect 14516 12152 14522 12164
rect 15010 12152 15016 12164
rect 14516 12124 15016 12152
rect 14516 12112 14522 12124
rect 15010 12112 15016 12124
rect 15068 12112 15074 12164
rect 15378 12112 15384 12164
rect 15436 12152 15442 12164
rect 15856 12152 15884 12183
rect 16114 12180 16120 12232
rect 16172 12220 16178 12232
rect 16485 12223 16543 12229
rect 16485 12220 16497 12223
rect 16172 12192 16497 12220
rect 16172 12180 16178 12192
rect 16485 12189 16497 12192
rect 16531 12189 16543 12223
rect 16485 12183 16543 12189
rect 17494 12180 17500 12232
rect 17552 12220 17558 12232
rect 18984 12220 19012 12251
rect 19076 12229 19104 12260
rect 20530 12248 20536 12260
rect 20588 12248 20594 12300
rect 17552 12192 19012 12220
rect 19061 12223 19119 12229
rect 17552 12180 17558 12192
rect 19061 12189 19073 12223
rect 19107 12189 19119 12223
rect 19061 12183 19119 12189
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 19702 12220 19708 12232
rect 19291 12192 19708 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 19702 12180 19708 12192
rect 19760 12180 19766 12232
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 15436 12124 15884 12152
rect 18601 12155 18659 12161
rect 15436 12112 15442 12124
rect 18601 12121 18613 12155
rect 18647 12152 18659 12155
rect 20088 12152 20116 12183
rect 20162 12180 20168 12232
rect 20220 12220 20226 12232
rect 20220 12192 20265 12220
rect 20220 12180 20226 12192
rect 18647 12124 20116 12152
rect 18647 12121 18659 12124
rect 18601 12115 18659 12121
rect 5960 12056 8708 12084
rect 5960 12044 5966 12056
rect 8938 12044 8944 12096
rect 8996 12084 9002 12096
rect 9125 12087 9183 12093
rect 9125 12084 9137 12087
rect 8996 12056 9137 12084
rect 8996 12044 9002 12056
rect 9125 12053 9137 12056
rect 9171 12053 9183 12087
rect 9125 12047 9183 12053
rect 10229 12087 10287 12093
rect 10229 12053 10241 12087
rect 10275 12084 10287 12087
rect 14550 12084 14556 12096
rect 10275 12056 14556 12084
rect 10275 12053 10287 12056
rect 10229 12047 10287 12053
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 16850 12044 16856 12096
rect 16908 12084 16914 12096
rect 19150 12084 19156 12096
rect 16908 12056 19156 12084
rect 16908 12044 16914 12056
rect 19150 12044 19156 12056
rect 19208 12044 19214 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 1946 11840 1952 11892
rect 2004 11880 2010 11892
rect 2133 11883 2191 11889
rect 2133 11880 2145 11883
rect 2004 11852 2145 11880
rect 2004 11840 2010 11852
rect 2133 11849 2145 11852
rect 2179 11849 2191 11883
rect 4154 11880 4160 11892
rect 4115 11852 4160 11880
rect 2133 11843 2191 11849
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 12434 11880 12440 11892
rect 7576 11852 12440 11880
rect 7193 11815 7251 11821
rect 7193 11812 7205 11815
rect 2976 11784 7205 11812
rect 2682 11744 2688 11756
rect 2643 11716 2688 11744
rect 2682 11704 2688 11716
rect 2740 11704 2746 11756
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11676 2651 11679
rect 2976 11676 3004 11784
rect 7193 11781 7205 11784
rect 7239 11781 7251 11815
rect 7193 11775 7251 11781
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11713 3847 11747
rect 4798 11744 4804 11756
rect 4759 11716 4804 11744
rect 3789 11707 3847 11713
rect 3510 11676 3516 11688
rect 2639 11648 3004 11676
rect 3471 11648 3516 11676
rect 2639 11645 2651 11648
rect 2593 11639 2651 11645
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 3804 11620 3832 11707
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 5350 11704 5356 11756
rect 5408 11744 5414 11756
rect 5721 11747 5779 11753
rect 5721 11744 5733 11747
rect 5408 11716 5733 11744
rect 5408 11704 5414 11716
rect 5721 11713 5733 11716
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 4062 11636 4068 11688
rect 4120 11676 4126 11688
rect 5902 11676 5908 11688
rect 4120 11648 5908 11676
rect 4120 11636 4126 11648
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 6641 11679 6699 11685
rect 6641 11645 6653 11679
rect 6687 11676 6699 11679
rect 7098 11676 7104 11688
rect 6687 11648 7104 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 7576 11685 7604 11852
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12526 11840 12532 11892
rect 12584 11880 12590 11892
rect 12584 11852 14044 11880
rect 12584 11840 12590 11852
rect 9214 11772 9220 11824
rect 9272 11812 9278 11824
rect 14016 11812 14044 11852
rect 14274 11840 14280 11892
rect 14332 11880 14338 11892
rect 14737 11883 14795 11889
rect 14737 11880 14749 11883
rect 14332 11852 14749 11880
rect 14332 11840 14338 11852
rect 14737 11849 14749 11852
rect 14783 11849 14795 11883
rect 16666 11880 16672 11892
rect 14737 11843 14795 11849
rect 14844 11852 16672 11880
rect 14844 11812 14872 11852
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 18601 11883 18659 11889
rect 18601 11849 18613 11883
rect 18647 11880 18659 11883
rect 19242 11880 19248 11892
rect 18647 11852 19248 11880
rect 18647 11849 18659 11852
rect 18601 11843 18659 11849
rect 19242 11840 19248 11852
rect 19300 11840 19306 11892
rect 9272 11784 11652 11812
rect 14016 11784 14872 11812
rect 14936 11784 15424 11812
rect 9272 11772 9278 11784
rect 7837 11747 7895 11753
rect 7837 11713 7849 11747
rect 7883 11744 7895 11747
rect 8021 11747 8079 11753
rect 8021 11744 8033 11747
rect 7883 11716 8033 11744
rect 7883 11713 7895 11716
rect 7837 11707 7895 11713
rect 8021 11713 8033 11716
rect 8067 11713 8079 11747
rect 10594 11744 10600 11756
rect 10555 11716 10600 11744
rect 8021 11707 8079 11713
rect 10594 11704 10600 11716
rect 10652 11704 10658 11756
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 11624 11753 11652 11784
rect 11609 11747 11667 11753
rect 10836 11716 11468 11744
rect 10836 11704 10842 11716
rect 7561 11679 7619 11685
rect 7561 11645 7573 11679
rect 7607 11645 7619 11679
rect 7561 11639 7619 11645
rect 7742 11636 7748 11688
rect 7800 11676 7806 11688
rect 8110 11676 8116 11688
rect 7800 11648 8116 11676
rect 7800 11636 7806 11648
rect 8110 11636 8116 11648
rect 8168 11676 8174 11688
rect 8205 11679 8263 11685
rect 8205 11676 8217 11679
rect 8168 11648 8217 11676
rect 8168 11636 8174 11648
rect 8205 11645 8217 11648
rect 8251 11645 8263 11679
rect 8205 11639 8263 11645
rect 8472 11679 8530 11685
rect 8472 11645 8484 11679
rect 8518 11676 8530 11679
rect 8846 11676 8852 11688
rect 8518 11648 8852 11676
rect 8518 11645 8530 11648
rect 8472 11639 8530 11645
rect 8846 11636 8852 11648
rect 8904 11636 8910 11688
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 9088 11648 10425 11676
rect 9088 11636 9094 11648
rect 10413 11645 10425 11648
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 10686 11636 10692 11688
rect 10744 11676 10750 11688
rect 11440 11685 11468 11716
rect 11609 11713 11621 11747
rect 11655 11713 11667 11747
rect 11609 11707 11667 11713
rect 11974 11704 11980 11756
rect 12032 11744 12038 11756
rect 12894 11744 12900 11756
rect 12032 11716 12900 11744
rect 12032 11704 12038 11716
rect 12894 11704 12900 11716
rect 12952 11744 12958 11756
rect 13081 11747 13139 11753
rect 13081 11744 13093 11747
rect 12952 11716 13093 11744
rect 12952 11704 12958 11716
rect 13081 11713 13093 11716
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 11425 11679 11483 11685
rect 10744 11648 11192 11676
rect 10744 11636 10750 11648
rect 3605 11611 3663 11617
rect 3605 11577 3617 11611
rect 3651 11608 3663 11611
rect 3694 11608 3700 11620
rect 3651 11580 3700 11608
rect 3651 11577 3663 11580
rect 3605 11571 3663 11577
rect 3694 11568 3700 11580
rect 3752 11568 3758 11620
rect 3786 11568 3792 11620
rect 3844 11608 3850 11620
rect 7653 11611 7711 11617
rect 3844 11580 6592 11608
rect 3844 11568 3850 11580
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 3145 11543 3203 11549
rect 3145 11540 3157 11543
rect 2547 11512 3157 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 3145 11509 3157 11512
rect 3191 11509 3203 11543
rect 3145 11503 3203 11509
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4525 11543 4583 11549
rect 4525 11540 4537 11543
rect 4304 11512 4537 11540
rect 4304 11500 4310 11512
rect 4525 11509 4537 11512
rect 4571 11509 4583 11543
rect 4525 11503 4583 11509
rect 4617 11543 4675 11549
rect 4617 11509 4629 11543
rect 4663 11540 4675 11543
rect 5169 11543 5227 11549
rect 5169 11540 5181 11543
rect 4663 11512 5181 11540
rect 4663 11509 4675 11512
rect 4617 11503 4675 11509
rect 5169 11509 5181 11512
rect 5215 11509 5227 11543
rect 5534 11540 5540 11552
rect 5495 11512 5540 11540
rect 5169 11503 5227 11509
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5629 11543 5687 11549
rect 5629 11509 5641 11543
rect 5675 11540 5687 11543
rect 6270 11540 6276 11552
rect 5675 11512 6276 11540
rect 5675 11509 5687 11512
rect 5629 11503 5687 11509
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 6454 11540 6460 11552
rect 6415 11512 6460 11540
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 6564 11540 6592 11580
rect 7653 11577 7665 11611
rect 7699 11608 7711 11611
rect 11164 11608 11192 11648
rect 11425 11645 11437 11679
rect 11471 11645 11483 11679
rect 11425 11639 11483 11645
rect 12066 11636 12072 11688
rect 12124 11676 12130 11688
rect 12250 11676 12256 11688
rect 12124 11648 12256 11676
rect 12124 11636 12130 11648
rect 12250 11636 12256 11648
rect 12308 11636 12314 11688
rect 13348 11679 13406 11685
rect 13348 11645 13360 11679
rect 13394 11676 13406 11679
rect 13630 11676 13636 11688
rect 13394 11648 13636 11676
rect 13394 11645 13406 11648
rect 13348 11639 13406 11645
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 14936 11676 14964 11784
rect 15010 11704 15016 11756
rect 15068 11744 15074 11756
rect 15289 11747 15347 11753
rect 15289 11744 15301 11747
rect 15068 11716 15301 11744
rect 15068 11704 15074 11716
rect 15289 11713 15301 11716
rect 15335 11713 15347 11747
rect 15396 11744 15424 11784
rect 17678 11772 17684 11824
rect 17736 11812 17742 11824
rect 17736 11784 19564 11812
rect 17736 11772 17742 11784
rect 19536 11753 19564 11784
rect 19521 11747 19579 11753
rect 15396 11716 16160 11744
rect 15289 11707 15347 11713
rect 13780 11648 14964 11676
rect 15105 11679 15163 11685
rect 13780 11636 13786 11648
rect 15105 11645 15117 11679
rect 15151 11676 15163 11679
rect 15930 11676 15936 11688
rect 15151 11648 15936 11676
rect 15151 11645 15163 11648
rect 15105 11639 15163 11645
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 16032 11679 16090 11685
rect 16032 11645 16044 11679
rect 16078 11645 16090 11679
rect 16132 11676 16160 11716
rect 19521 11713 19533 11747
rect 19567 11744 19579 11747
rect 20533 11747 20591 11753
rect 20533 11744 20545 11747
rect 19567 11716 20545 11744
rect 19567 11713 19579 11716
rect 19521 11707 19579 11713
rect 20533 11713 20545 11716
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 16574 11676 16580 11688
rect 16132 11648 16580 11676
rect 16032 11639 16090 11645
rect 11517 11611 11575 11617
rect 11517 11608 11529 11611
rect 7699 11580 11100 11608
rect 11164 11580 11529 11608
rect 7699 11577 7711 11580
rect 7653 11571 7711 11577
rect 8021 11543 8079 11549
rect 8021 11540 8033 11543
rect 6564 11512 8033 11540
rect 8021 11509 8033 11512
rect 8067 11540 8079 11543
rect 8938 11540 8944 11552
rect 8067 11512 8944 11540
rect 8067 11509 8079 11512
rect 8021 11503 8079 11509
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9122 11500 9128 11552
rect 9180 11540 9186 11552
rect 9585 11543 9643 11549
rect 9585 11540 9597 11543
rect 9180 11512 9597 11540
rect 9180 11500 9186 11512
rect 9585 11509 9597 11512
rect 9631 11509 9643 11543
rect 10042 11540 10048 11552
rect 10003 11512 10048 11540
rect 9585 11503 9643 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 11072 11549 11100 11580
rect 11517 11577 11529 11580
rect 11563 11577 11575 11611
rect 11517 11571 11575 11577
rect 11606 11568 11612 11620
rect 11664 11608 11670 11620
rect 13814 11608 13820 11620
rect 11664 11580 13820 11608
rect 11664 11568 11670 11580
rect 13814 11568 13820 11580
rect 13872 11608 13878 11620
rect 13872 11580 14504 11608
rect 13872 11568 13878 11580
rect 10505 11543 10563 11549
rect 10505 11540 10517 11543
rect 10468 11512 10517 11540
rect 10468 11500 10474 11512
rect 10505 11509 10517 11512
rect 10551 11509 10563 11543
rect 10505 11503 10563 11509
rect 11057 11543 11115 11549
rect 11057 11509 11069 11543
rect 11103 11509 11115 11543
rect 11057 11503 11115 11509
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 14366 11540 14372 11552
rect 11388 11512 14372 11540
rect 11388 11500 11394 11512
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 14476 11549 14504 11580
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 15197 11611 15255 11617
rect 15197 11608 15209 11611
rect 15068 11580 15209 11608
rect 15068 11568 15074 11580
rect 15197 11577 15209 11580
rect 15243 11577 15255 11611
rect 15197 11571 15255 11577
rect 16047 11608 16075 11639
rect 16574 11636 16580 11648
rect 16632 11636 16638 11688
rect 18414 11676 18420 11688
rect 18375 11648 18420 11676
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 19337 11679 19395 11685
rect 19337 11645 19349 11679
rect 19383 11676 19395 11679
rect 19978 11676 19984 11688
rect 19383 11648 19984 11676
rect 19383 11645 19395 11648
rect 19337 11639 19395 11645
rect 19978 11636 19984 11648
rect 20036 11636 20042 11688
rect 16114 11608 16120 11620
rect 16047 11580 16120 11608
rect 14461 11543 14519 11549
rect 14461 11509 14473 11543
rect 14507 11509 14519 11543
rect 14461 11503 14519 11509
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 16047 11540 16075 11580
rect 16114 11568 16120 11580
rect 16172 11568 16178 11620
rect 16292 11611 16350 11617
rect 16292 11577 16304 11611
rect 16338 11608 16350 11611
rect 16850 11608 16856 11620
rect 16338 11580 16856 11608
rect 16338 11577 16350 11580
rect 16292 11571 16350 11577
rect 16850 11568 16856 11580
rect 16908 11568 16914 11620
rect 17126 11568 17132 11620
rect 17184 11608 17190 11620
rect 19429 11611 19487 11617
rect 19429 11608 19441 11611
rect 17184 11580 19441 11608
rect 17184 11568 17190 11580
rect 19429 11577 19441 11580
rect 19475 11577 19487 11611
rect 19429 11571 19487 11577
rect 20349 11611 20407 11617
rect 20349 11577 20361 11611
rect 20395 11608 20407 11611
rect 20530 11608 20536 11620
rect 20395 11580 20536 11608
rect 20395 11577 20407 11580
rect 20349 11571 20407 11577
rect 20530 11568 20536 11580
rect 20588 11568 20594 11620
rect 17402 11540 17408 11552
rect 15344 11512 16075 11540
rect 17363 11512 17408 11540
rect 15344 11500 15350 11512
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 18874 11500 18880 11552
rect 18932 11540 18938 11552
rect 18969 11543 19027 11549
rect 18969 11540 18981 11543
rect 18932 11512 18981 11540
rect 18932 11500 18938 11512
rect 18969 11509 18981 11512
rect 19015 11509 19027 11543
rect 18969 11503 19027 11509
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 19981 11543 20039 11549
rect 19981 11540 19993 11543
rect 19576 11512 19993 11540
rect 19576 11500 19582 11512
rect 19981 11509 19993 11512
rect 20027 11509 20039 11543
rect 19981 11503 20039 11509
rect 20162 11500 20168 11552
rect 20220 11540 20226 11552
rect 20441 11543 20499 11549
rect 20441 11540 20453 11543
rect 20220 11512 20453 11540
rect 20220 11500 20226 11512
rect 20441 11509 20453 11512
rect 20487 11509 20499 11543
rect 20441 11503 20499 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 2682 11296 2688 11348
rect 2740 11336 2746 11348
rect 2869 11339 2927 11345
rect 2869 11336 2881 11339
rect 2740 11308 2881 11336
rect 2740 11296 2746 11308
rect 2869 11305 2881 11308
rect 2915 11305 2927 11339
rect 2869 11299 2927 11305
rect 5442 11296 5448 11348
rect 5500 11296 5506 11348
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 5721 11339 5779 11345
rect 5721 11336 5733 11339
rect 5592 11308 5733 11336
rect 5592 11296 5598 11308
rect 5721 11305 5733 11308
rect 5767 11305 5779 11339
rect 5721 11299 5779 11305
rect 5994 11296 6000 11348
rect 6052 11336 6058 11348
rect 6181 11339 6239 11345
rect 6181 11336 6193 11339
rect 6052 11308 6193 11336
rect 6052 11296 6058 11308
rect 6181 11305 6193 11308
rect 6227 11305 6239 11339
rect 6181 11299 6239 11305
rect 6270 11296 6276 11348
rect 6328 11336 6334 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 6328 11308 6745 11336
rect 6328 11296 6334 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 6733 11299 6791 11305
rect 7006 11296 7012 11348
rect 7064 11336 7070 11348
rect 8754 11336 8760 11348
rect 7064 11308 8760 11336
rect 7064 11296 7070 11308
rect 8754 11296 8760 11308
rect 8812 11296 8818 11348
rect 8941 11339 8999 11345
rect 8941 11305 8953 11339
rect 8987 11336 8999 11339
rect 9030 11336 9036 11348
rect 8987 11308 9036 11336
rect 8987 11305 8999 11308
rect 8941 11299 8999 11305
rect 9030 11296 9036 11308
rect 9088 11296 9094 11348
rect 10413 11339 10471 11345
rect 10413 11305 10425 11339
rect 10459 11336 10471 11339
rect 12621 11339 12679 11345
rect 10459 11308 12388 11336
rect 10459 11305 10471 11308
rect 10413 11299 10471 11305
rect 1486 11228 1492 11280
rect 1544 11268 1550 11280
rect 4154 11268 4160 11280
rect 1544 11240 4160 11268
rect 1544 11228 1550 11240
rect 1756 11203 1814 11209
rect 1756 11169 1768 11203
rect 1802 11200 1814 11203
rect 2498 11200 2504 11212
rect 1802 11172 2504 11200
rect 1802 11169 1814 11172
rect 1756 11163 1814 11169
rect 2498 11160 2504 11172
rect 2556 11160 2562 11212
rect 4080 11209 4108 11240
rect 4154 11228 4160 11240
rect 4212 11228 4218 11280
rect 5460 11268 5488 11296
rect 5902 11268 5908 11280
rect 5460 11240 5908 11268
rect 5902 11228 5908 11240
rect 5960 11228 5966 11280
rect 7101 11271 7159 11277
rect 7101 11237 7113 11271
rect 7147 11268 7159 11271
rect 9582 11268 9588 11280
rect 7147 11240 9588 11268
rect 7147 11237 7159 11240
rect 7101 11231 7159 11237
rect 9582 11228 9588 11240
rect 9640 11228 9646 11280
rect 10042 11228 10048 11280
rect 10100 11268 10106 11280
rect 11146 11268 11152 11280
rect 10100 11240 11152 11268
rect 10100 11228 10106 11240
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 12360 11268 12388 11308
rect 12621 11305 12633 11339
rect 12667 11336 12679 11339
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 12667 11308 13277 11336
rect 12667 11305 12679 11308
rect 12621 11299 12679 11305
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 13633 11339 13691 11345
rect 13633 11305 13645 11339
rect 13679 11336 13691 11339
rect 13722 11336 13728 11348
rect 13679 11308 13728 11336
rect 13679 11305 13691 11308
rect 13633 11299 13691 11305
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 14737 11339 14795 11345
rect 14737 11305 14749 11339
rect 14783 11336 14795 11339
rect 15102 11336 15108 11348
rect 14783 11308 15108 11336
rect 14783 11305 14795 11308
rect 14737 11299 14795 11305
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 16669 11339 16727 11345
rect 16669 11305 16681 11339
rect 16715 11336 16727 11339
rect 16850 11336 16856 11348
rect 16715 11308 16856 11336
rect 16715 11305 16727 11308
rect 16669 11299 16727 11305
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 17313 11339 17371 11345
rect 17313 11305 17325 11339
rect 17359 11336 17371 11339
rect 17586 11336 17592 11348
rect 17359 11308 17592 11336
rect 17359 11305 17371 11308
rect 17313 11299 17371 11305
rect 17586 11296 17592 11308
rect 17644 11336 17650 11348
rect 17770 11336 17776 11348
rect 17644 11308 17776 11336
rect 17644 11296 17650 11308
rect 17770 11296 17776 11308
rect 17828 11296 17834 11348
rect 18414 11296 18420 11348
rect 18472 11296 18478 11348
rect 18509 11339 18567 11345
rect 18509 11305 18521 11339
rect 18555 11336 18567 11339
rect 18782 11336 18788 11348
rect 18555 11308 18788 11336
rect 18555 11305 18567 11308
rect 18509 11299 18567 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 18877 11339 18935 11345
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 19334 11336 19340 11348
rect 18923 11308 19340 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 19334 11296 19340 11308
rect 19392 11296 19398 11348
rect 20622 11296 20628 11348
rect 20680 11336 20686 11348
rect 20901 11339 20959 11345
rect 20901 11336 20913 11339
rect 20680 11308 20913 11336
rect 20680 11296 20686 11308
rect 20901 11305 20913 11308
rect 20947 11305 20959 11339
rect 20901 11299 20959 11305
rect 12713 11271 12771 11277
rect 12713 11268 12725 11271
rect 12360 11240 12725 11268
rect 12713 11237 12725 11240
rect 12759 11237 12771 11271
rect 12713 11231 12771 11237
rect 14366 11228 14372 11280
rect 14424 11268 14430 11280
rect 17405 11271 17463 11277
rect 17405 11268 17417 11271
rect 14424 11240 17417 11268
rect 14424 11228 14430 11240
rect 17405 11237 17417 11240
rect 17451 11237 17463 11271
rect 17405 11231 17463 11237
rect 4065 11203 4123 11209
rect 4065 11169 4077 11203
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 4332 11203 4390 11209
rect 4332 11169 4344 11203
rect 4378 11200 4390 11203
rect 4798 11200 4804 11212
rect 4378 11172 4804 11200
rect 4378 11169 4390 11172
rect 4332 11163 4390 11169
rect 4798 11160 4804 11172
rect 4856 11200 4862 11212
rect 4856 11172 5396 11200
rect 4856 11160 4862 11172
rect 1486 11132 1492 11144
rect 1447 11104 1492 11132
rect 1486 11092 1492 11104
rect 1544 11092 1550 11144
rect 5368 11132 5396 11172
rect 5442 11160 5448 11212
rect 5500 11200 5506 11212
rect 6089 11203 6147 11209
rect 6089 11200 6101 11203
rect 5500 11172 6101 11200
rect 5500 11160 5506 11172
rect 6089 11169 6101 11172
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 7193 11203 7251 11209
rect 7193 11169 7205 11203
rect 7239 11200 7251 11203
rect 8202 11200 8208 11212
rect 7239 11172 8208 11200
rect 7239 11169 7251 11172
rect 7193 11163 7251 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 10410 11200 10416 11212
rect 9048 11172 10416 11200
rect 9048 11141 9076 11172
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 10781 11203 10839 11209
rect 10781 11169 10793 11203
rect 10827 11169 10839 11203
rect 10781 11163 10839 11169
rect 12161 11203 12219 11209
rect 12161 11169 12173 11203
rect 12207 11200 12219 11203
rect 12207 11172 13584 11200
rect 12207 11169 12219 11172
rect 12161 11163 12219 11169
rect 6273 11135 6331 11141
rect 6273 11132 6285 11135
rect 5368 11104 6285 11132
rect 6273 11101 6285 11104
rect 6319 11132 6331 11135
rect 7285 11135 7343 11141
rect 7285 11132 7297 11135
rect 6319 11104 7297 11132
rect 6319 11101 6331 11104
rect 6273 11095 6331 11101
rect 7285 11101 7297 11104
rect 7331 11101 7343 11135
rect 7285 11095 7343 11101
rect 9033 11135 9091 11141
rect 9033 11101 9045 11135
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 6914 11024 6920 11076
rect 6972 11064 6978 11076
rect 9048 11064 9076 11095
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 9180 11104 9225 11132
rect 9180 11092 9186 11104
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 10318 11132 10324 11144
rect 9916 11104 10324 11132
rect 9916 11092 9922 11104
rect 10318 11092 10324 11104
rect 10376 11132 10382 11144
rect 10796 11132 10824 11163
rect 10376 11104 10824 11132
rect 10873 11135 10931 11141
rect 10376 11092 10382 11104
rect 10873 11101 10885 11135
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 11057 11135 11115 11141
rect 11057 11101 11069 11135
rect 11103 11132 11115 11135
rect 11606 11132 11612 11144
rect 11103 11104 11612 11132
rect 11103 11101 11115 11104
rect 11057 11095 11115 11101
rect 6972 11036 9076 11064
rect 6972 11024 6978 11036
rect 9306 11024 9312 11076
rect 9364 11064 9370 11076
rect 9490 11064 9496 11076
rect 9364 11036 9496 11064
rect 9364 11024 9370 11036
rect 9490 11024 9496 11036
rect 9548 11064 9554 11076
rect 10888 11064 10916 11095
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 12342 11092 12348 11144
rect 12400 11132 12406 11144
rect 12802 11132 12808 11144
rect 12400 11104 12808 11132
rect 12400 11092 12406 11104
rect 12802 11092 12808 11104
rect 12860 11092 12866 11144
rect 9548 11036 10916 11064
rect 9548 11024 9554 11036
rect 11238 11024 11244 11076
rect 11296 11064 11302 11076
rect 11974 11064 11980 11076
rect 11296 11036 11980 11064
rect 11296 11024 11302 11036
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 12253 11067 12311 11073
rect 12253 11033 12265 11067
rect 12299 11064 12311 11067
rect 12894 11064 12900 11076
rect 12299 11036 12900 11064
rect 12299 11033 12311 11036
rect 12253 11027 12311 11033
rect 12894 11024 12900 11036
rect 12952 11024 12958 11076
rect 13556 11064 13584 11172
rect 13998 11160 14004 11212
rect 14056 11200 14062 11212
rect 14461 11203 14519 11209
rect 14461 11200 14473 11203
rect 14056 11172 14473 11200
rect 14056 11160 14062 11172
rect 14461 11169 14473 11172
rect 14507 11169 14519 11203
rect 14461 11163 14519 11169
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11200 14703 11203
rect 15545 11203 15603 11209
rect 15545 11200 15557 11203
rect 14691 11172 15557 11200
rect 14691 11169 14703 11172
rect 14645 11163 14703 11169
rect 15545 11169 15557 11172
rect 15591 11200 15603 11203
rect 18313 11203 18371 11209
rect 18313 11200 18325 11203
rect 15591 11172 17080 11200
rect 15591 11169 15603 11172
rect 15545 11163 15603 11169
rect 13722 11132 13728 11144
rect 13683 11104 13728 11132
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 13872 11104 13917 11132
rect 13872 11092 13878 11104
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 15286 11132 15292 11144
rect 14608 11104 15292 11132
rect 14608 11092 14614 11104
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 17052 11132 17080 11172
rect 18248 11172 18325 11200
rect 17497 11135 17555 11141
rect 17497 11132 17509 11135
rect 17052 11104 17509 11132
rect 17497 11101 17509 11104
rect 17543 11132 17555 11135
rect 17678 11132 17684 11144
rect 17543 11104 17684 11132
rect 17543 11101 17555 11104
rect 17497 11095 17555 11101
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 17954 11092 17960 11144
rect 18012 11132 18018 11144
rect 18248 11132 18276 11172
rect 18313 11169 18325 11172
rect 18359 11169 18371 11203
rect 18432 11200 18460 11296
rect 18693 11271 18751 11277
rect 18693 11237 18705 11271
rect 18739 11268 18751 11271
rect 19245 11271 19303 11277
rect 19245 11268 19257 11271
rect 18739 11240 19257 11268
rect 18739 11237 18751 11240
rect 18693 11231 18751 11237
rect 19245 11237 19257 11240
rect 19291 11237 19303 11271
rect 19245 11231 19303 11237
rect 20070 11228 20076 11280
rect 20128 11268 20134 11280
rect 20257 11271 20315 11277
rect 20257 11268 20269 11271
rect 20128 11240 20269 11268
rect 20128 11228 20134 11240
rect 20257 11237 20269 11240
rect 20303 11237 20315 11271
rect 20257 11231 20315 11237
rect 19337 11203 19395 11209
rect 19337 11200 19349 11203
rect 18432 11172 19349 11200
rect 18313 11163 18371 11169
rect 19337 11169 19349 11172
rect 19383 11169 19395 11203
rect 19981 11203 20039 11209
rect 19981 11200 19993 11203
rect 19337 11163 19395 11169
rect 19444 11172 19993 11200
rect 19444 11132 19472 11172
rect 19981 11169 19993 11172
rect 20027 11169 20039 11203
rect 19981 11163 20039 11169
rect 18012 11104 18276 11132
rect 18708 11104 19472 11132
rect 19521 11135 19579 11141
rect 18012 11092 18018 11104
rect 14277 11067 14335 11073
rect 14277 11064 14289 11067
rect 13556 11036 14289 11064
rect 14277 11033 14289 11036
rect 14323 11064 14335 11067
rect 14826 11064 14832 11076
rect 14323 11036 14832 11064
rect 14323 11033 14335 11036
rect 14277 11027 14335 11033
rect 14826 11024 14832 11036
rect 14884 11024 14890 11076
rect 16574 11024 16580 11076
rect 16632 11064 16638 11076
rect 18708 11064 18736 11104
rect 19521 11101 19533 11135
rect 19567 11132 19579 11135
rect 19610 11132 19616 11144
rect 19567 11104 19616 11132
rect 19567 11101 19579 11104
rect 19521 11095 19579 11101
rect 19610 11092 19616 11104
rect 19668 11092 19674 11144
rect 16632 11036 18736 11064
rect 16632 11024 16638 11036
rect 5350 10956 5356 11008
rect 5408 10996 5414 11008
rect 5445 10999 5503 11005
rect 5445 10996 5457 10999
rect 5408 10968 5457 10996
rect 5408 10956 5414 10968
rect 5445 10965 5457 10968
rect 5491 10965 5503 10999
rect 8570 10996 8576 11008
rect 8531 10968 8576 10996
rect 5445 10959 5503 10965
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 8662 10956 8668 11008
rect 8720 10996 8726 11008
rect 9214 10996 9220 11008
rect 8720 10968 9220 10996
rect 8720 10956 8726 10968
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 14645 10999 14703 11005
rect 14645 10996 14657 10999
rect 10652 10968 14657 10996
rect 10652 10956 10658 10968
rect 14645 10965 14657 10968
rect 14691 10965 14703 10999
rect 14645 10959 14703 10965
rect 14734 10956 14740 11008
rect 14792 10996 14798 11008
rect 15194 10996 15200 11008
rect 14792 10968 15200 10996
rect 14792 10956 14798 10968
rect 15194 10956 15200 10968
rect 15252 10956 15258 11008
rect 16942 10996 16948 11008
rect 16903 10968 16948 10996
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 17862 10956 17868 11008
rect 17920 10996 17926 11008
rect 18693 10999 18751 11005
rect 18693 10996 18705 10999
rect 17920 10968 18705 10996
rect 17920 10956 17926 10968
rect 18693 10965 18705 10968
rect 18739 10965 18751 10999
rect 18693 10959 18751 10965
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 1673 10795 1731 10801
rect 1673 10761 1685 10795
rect 1719 10792 1731 10795
rect 1854 10792 1860 10804
rect 1719 10764 1860 10792
rect 1719 10761 1731 10764
rect 1673 10755 1731 10761
rect 1854 10752 1860 10764
rect 1912 10752 1918 10804
rect 3881 10795 3939 10801
rect 3881 10761 3893 10795
rect 3927 10792 3939 10795
rect 4246 10792 4252 10804
rect 3927 10764 4252 10792
rect 3927 10761 3939 10764
rect 3881 10755 3939 10761
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 4890 10752 4896 10804
rect 4948 10792 4954 10804
rect 5258 10792 5264 10804
rect 4948 10764 5264 10792
rect 4948 10752 4954 10764
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 8665 10795 8723 10801
rect 8665 10761 8677 10795
rect 8711 10792 8723 10795
rect 10134 10792 10140 10804
rect 8711 10764 10140 10792
rect 8711 10761 8723 10764
rect 8665 10755 8723 10761
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 11054 10792 11060 10804
rect 10704 10764 11060 10792
rect 4338 10684 4344 10736
rect 4396 10724 4402 10736
rect 4706 10724 4712 10736
rect 4396 10696 4712 10724
rect 4396 10684 4402 10696
rect 4706 10684 4712 10696
rect 4764 10724 4770 10736
rect 5166 10724 5172 10736
rect 4764 10696 5172 10724
rect 4764 10684 4770 10696
rect 5166 10684 5172 10696
rect 5224 10684 5230 10736
rect 7852 10696 9260 10724
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2682 10656 2688 10668
rect 2363 10628 2688 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 3329 10659 3387 10665
rect 3329 10625 3341 10659
rect 3375 10656 3387 10659
rect 3786 10656 3792 10668
rect 3375 10628 3792 10656
rect 3375 10625 3387 10628
rect 3329 10619 3387 10625
rect 2498 10548 2504 10600
rect 2556 10588 2562 10600
rect 3344 10588 3372 10619
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10656 4583 10659
rect 5350 10656 5356 10668
rect 4571 10628 5356 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10656 5595 10659
rect 5994 10656 6000 10668
rect 5583 10628 6000 10656
rect 5583 10625 5595 10628
rect 5537 10619 5595 10625
rect 5994 10616 6000 10628
rect 6052 10656 6058 10668
rect 6362 10656 6368 10668
rect 6052 10628 6368 10656
rect 6052 10616 6058 10628
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 7650 10616 7656 10668
rect 7708 10656 7714 10668
rect 7852 10665 7880 10696
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7708 10628 7849 10656
rect 7708 10616 7714 10628
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 8570 10616 8576 10668
rect 8628 10656 8634 10668
rect 9232 10665 9260 10696
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 8628 10628 9137 10656
rect 8628 10616 8634 10628
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10656 9275 10659
rect 9306 10656 9312 10668
rect 9263 10628 9312 10656
rect 9263 10625 9275 10628
rect 9217 10619 9275 10625
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 10704 10665 10732 10764
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 12069 10795 12127 10801
rect 12069 10761 12081 10795
rect 12115 10792 12127 10795
rect 12342 10792 12348 10804
rect 12115 10764 12348 10792
rect 12115 10761 12127 10764
rect 12069 10755 12127 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 14553 10795 14611 10801
rect 14553 10761 14565 10795
rect 14599 10792 14611 10795
rect 14734 10792 14740 10804
rect 14599 10764 14740 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 14734 10752 14740 10764
rect 14792 10752 14798 10804
rect 14921 10795 14979 10801
rect 14921 10761 14933 10795
rect 14967 10792 14979 10795
rect 15010 10792 15016 10804
rect 14967 10764 15016 10792
rect 14967 10761 14979 10764
rect 14921 10755 14979 10761
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 15102 10752 15108 10804
rect 15160 10792 15166 10804
rect 17402 10792 17408 10804
rect 15160 10764 17408 10792
rect 15160 10752 15166 10764
rect 17402 10752 17408 10764
rect 17460 10752 17466 10804
rect 18417 10795 18475 10801
rect 18417 10761 18429 10795
rect 18463 10792 18475 10795
rect 18506 10792 18512 10804
rect 18463 10764 18512 10792
rect 18463 10761 18475 10764
rect 18417 10755 18475 10761
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 19245 10795 19303 10801
rect 19245 10792 19257 10795
rect 18932 10764 19257 10792
rect 18932 10752 18938 10764
rect 19245 10761 19257 10764
rect 19291 10761 19303 10795
rect 19245 10755 19303 10761
rect 19978 10752 19984 10804
rect 20036 10752 20042 10804
rect 12526 10684 12532 10736
rect 12584 10724 12590 10736
rect 16574 10724 16580 10736
rect 12584 10696 16580 10724
rect 12584 10684 12590 10696
rect 16574 10684 16580 10696
rect 16632 10684 16638 10736
rect 19996 10724 20024 10752
rect 16684 10696 20024 10724
rect 10229 10659 10287 10665
rect 10229 10656 10241 10659
rect 9456 10628 10241 10656
rect 9456 10616 9462 10628
rect 10229 10625 10241 10628
rect 10275 10625 10287 10659
rect 10229 10619 10287 10625
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10625 10747 10659
rect 12894 10656 12900 10668
rect 12855 10628 12900 10656
rect 10689 10619 10747 10625
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 2556 10560 3372 10588
rect 2556 10548 2562 10560
rect 4246 10548 4252 10600
rect 4304 10588 4310 10600
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 4304 10560 4353 10588
rect 4304 10548 4310 10560
rect 4341 10557 4353 10560
rect 4387 10557 4399 10591
rect 4341 10551 4399 10557
rect 4890 10548 4896 10600
rect 4948 10548 4954 10600
rect 6454 10548 6460 10600
rect 6512 10588 6518 10600
rect 8481 10591 8539 10597
rect 8481 10588 8493 10591
rect 6512 10560 8493 10588
rect 6512 10548 6518 10560
rect 8481 10557 8493 10560
rect 8527 10557 8539 10591
rect 8481 10551 8539 10557
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9824 10560 10057 10588
rect 9824 10548 9830 10560
rect 10045 10557 10057 10560
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 10137 10591 10195 10597
rect 10137 10557 10149 10591
rect 10183 10588 10195 10591
rect 10778 10588 10784 10600
rect 10183 10560 10784 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 2041 10523 2099 10529
rect 2041 10489 2053 10523
rect 2087 10520 2099 10523
rect 3145 10523 3203 10529
rect 2087 10492 2728 10520
rect 2087 10489 2099 10492
rect 2041 10483 2099 10489
rect 1854 10412 1860 10464
rect 1912 10452 1918 10464
rect 2700 10461 2728 10492
rect 3145 10489 3157 10523
rect 3191 10520 3203 10523
rect 4908 10520 4936 10548
rect 3191 10492 4936 10520
rect 3191 10489 3203 10492
rect 3145 10483 3203 10489
rect 5166 10480 5172 10532
rect 5224 10520 5230 10532
rect 5353 10523 5411 10529
rect 5353 10520 5365 10523
rect 5224 10492 5365 10520
rect 5224 10480 5230 10492
rect 5353 10489 5365 10492
rect 5399 10489 5411 10523
rect 8938 10520 8944 10532
rect 5353 10483 5411 10489
rect 7300 10492 8944 10520
rect 2133 10455 2191 10461
rect 2133 10452 2145 10455
rect 1912 10424 2145 10452
rect 1912 10412 1918 10424
rect 2133 10421 2145 10424
rect 2179 10421 2191 10455
rect 2133 10415 2191 10421
rect 2685 10455 2743 10461
rect 2685 10421 2697 10455
rect 2731 10421 2743 10455
rect 3050 10452 3056 10464
rect 3011 10424 3056 10452
rect 2685 10415 2743 10421
rect 3050 10412 3056 10424
rect 3108 10412 3114 10464
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 4249 10455 4307 10461
rect 4249 10452 4261 10455
rect 4120 10424 4261 10452
rect 4120 10412 4126 10424
rect 4249 10421 4261 10424
rect 4295 10421 4307 10455
rect 4249 10415 4307 10421
rect 4798 10412 4804 10464
rect 4856 10452 4862 10464
rect 4893 10455 4951 10461
rect 4893 10452 4905 10455
rect 4856 10424 4905 10452
rect 4856 10412 4862 10424
rect 4893 10421 4905 10424
rect 4939 10421 4951 10455
rect 5258 10452 5264 10464
rect 5219 10424 5264 10452
rect 4893 10415 4951 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 7300 10461 7328 10492
rect 8938 10480 8944 10492
rect 8996 10480 9002 10532
rect 9033 10523 9091 10529
rect 9033 10489 9045 10523
rect 9079 10520 9091 10523
rect 10060 10520 10088 10551
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 10962 10597 10968 10600
rect 10956 10588 10968 10597
rect 10923 10560 10968 10588
rect 10956 10551 10968 10560
rect 10962 10548 10968 10551
rect 11020 10548 11026 10600
rect 12250 10588 12256 10600
rect 11072 10560 12256 10588
rect 11072 10520 11100 10560
rect 12250 10548 12256 10560
rect 12308 10548 12314 10600
rect 12342 10548 12348 10600
rect 12400 10588 12406 10600
rect 13004 10588 13032 10619
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 14185 10659 14243 10665
rect 14185 10656 14197 10659
rect 13872 10628 14197 10656
rect 13872 10616 13878 10628
rect 14185 10625 14197 10628
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 15378 10616 15384 10668
rect 15436 10656 15442 10668
rect 15473 10659 15531 10665
rect 15473 10656 15485 10659
rect 15436 10628 15485 10656
rect 15436 10616 15442 10628
rect 15473 10625 15485 10628
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 15562 10616 15568 10668
rect 15620 10656 15626 10668
rect 16684 10656 16712 10696
rect 15620 10628 16712 10656
rect 16761 10659 16819 10665
rect 15620 10616 15626 10628
rect 16761 10625 16773 10659
rect 16807 10656 16819 10659
rect 16850 10656 16856 10668
rect 16807 10628 16856 10656
rect 16807 10625 16819 10628
rect 16761 10619 16819 10625
rect 16850 10616 16856 10628
rect 16908 10656 16914 10668
rect 17770 10656 17776 10668
rect 16908 10628 17776 10656
rect 16908 10616 16914 10628
rect 17770 10616 17776 10628
rect 17828 10656 17834 10668
rect 18874 10656 18880 10668
rect 17828 10628 18880 10656
rect 17828 10616 17834 10628
rect 18874 10616 18880 10628
rect 18932 10656 18938 10668
rect 18969 10659 19027 10665
rect 18969 10656 18981 10659
rect 18932 10628 18981 10656
rect 18932 10616 18938 10628
rect 18969 10625 18981 10628
rect 19015 10625 19027 10659
rect 18969 10619 19027 10625
rect 19610 10616 19616 10668
rect 19668 10656 19674 10668
rect 19981 10659 20039 10665
rect 19981 10656 19993 10659
rect 19668 10628 19993 10656
rect 19668 10616 19674 10628
rect 19981 10625 19993 10628
rect 20027 10625 20039 10659
rect 19981 10619 20039 10625
rect 12400 10560 13032 10588
rect 14001 10591 14059 10597
rect 12400 10548 12406 10560
rect 14001 10557 14013 10591
rect 14047 10588 14059 10591
rect 14090 10588 14096 10600
rect 14047 10560 14096 10588
rect 14047 10557 14059 10560
rect 14001 10551 14059 10557
rect 14090 10548 14096 10560
rect 14148 10548 14154 10600
rect 14826 10588 14832 10600
rect 14787 10560 14832 10588
rect 14826 10548 14832 10560
rect 14884 10548 14890 10600
rect 15010 10548 15016 10600
rect 15068 10588 15074 10600
rect 15289 10591 15347 10597
rect 15289 10588 15301 10591
rect 15068 10560 15301 10588
rect 15068 10548 15074 10560
rect 15289 10557 15301 10560
rect 15335 10588 15347 10591
rect 15838 10588 15844 10600
rect 15335 10560 15844 10588
rect 15335 10557 15347 10560
rect 15289 10551 15347 10557
rect 15838 10548 15844 10560
rect 15896 10548 15902 10600
rect 16485 10591 16543 10597
rect 16485 10557 16497 10591
rect 16531 10588 16543 10591
rect 16942 10588 16948 10600
rect 16531 10560 16948 10588
rect 16531 10557 16543 10560
rect 16485 10551 16543 10557
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 18138 10548 18144 10600
rect 18196 10588 18202 10600
rect 18690 10588 18696 10600
rect 18196 10560 18696 10588
rect 18196 10548 18202 10560
rect 18690 10548 18696 10560
rect 18748 10548 18754 10600
rect 18785 10591 18843 10597
rect 18785 10557 18797 10591
rect 18831 10588 18843 10591
rect 19518 10588 19524 10600
rect 18831 10560 19524 10588
rect 18831 10557 18843 10560
rect 18785 10551 18843 10557
rect 19518 10548 19524 10560
rect 19576 10548 19582 10600
rect 19702 10548 19708 10600
rect 19760 10588 19766 10600
rect 20441 10591 20499 10597
rect 20441 10588 20453 10591
rect 19760 10560 20453 10588
rect 19760 10548 19766 10560
rect 20441 10557 20453 10560
rect 20487 10557 20499 10591
rect 20441 10551 20499 10557
rect 9079 10492 9720 10520
rect 10060 10492 11100 10520
rect 9079 10489 9091 10492
rect 9033 10483 9091 10489
rect 7285 10455 7343 10461
rect 7285 10421 7297 10455
rect 7331 10421 7343 10455
rect 7285 10415 7343 10421
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 7653 10455 7711 10461
rect 7653 10452 7665 10455
rect 7524 10424 7665 10452
rect 7524 10412 7530 10424
rect 7653 10421 7665 10424
rect 7699 10421 7711 10455
rect 7653 10415 7711 10421
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 8294 10452 8300 10464
rect 7800 10424 7845 10452
rect 8207 10424 8300 10452
rect 7800 10412 7806 10424
rect 8294 10412 8300 10424
rect 8352 10452 8358 10464
rect 8570 10452 8576 10464
rect 8352 10424 8576 10452
rect 8352 10412 8358 10424
rect 8570 10412 8576 10424
rect 8628 10412 8634 10464
rect 9692 10461 9720 10492
rect 11146 10480 11152 10532
rect 11204 10520 11210 10532
rect 16577 10523 16635 10529
rect 16577 10520 16589 10523
rect 11204 10492 16589 10520
rect 11204 10480 11210 10492
rect 16577 10489 16589 10492
rect 16623 10489 16635 10523
rect 16577 10483 16635 10489
rect 16758 10480 16764 10532
rect 16816 10520 16822 10532
rect 17770 10520 17776 10532
rect 16816 10492 17776 10520
rect 16816 10480 16822 10492
rect 17770 10480 17776 10492
rect 17828 10520 17834 10532
rect 19797 10523 19855 10529
rect 17828 10492 19564 10520
rect 17828 10480 17834 10492
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10421 9735 10455
rect 9677 10415 9735 10421
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12526 10452 12532 10464
rect 12483 10424 12532 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 12802 10452 12808 10464
rect 12763 10424 12808 10452
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13354 10412 13360 10464
rect 13412 10452 13418 10464
rect 13633 10455 13691 10461
rect 13633 10452 13645 10455
rect 13412 10424 13645 10452
rect 13412 10412 13418 10424
rect 13633 10421 13645 10424
rect 13679 10421 13691 10455
rect 13633 10415 13691 10421
rect 14093 10455 14151 10461
rect 14093 10421 14105 10455
rect 14139 10452 14151 10455
rect 14461 10455 14519 10461
rect 14461 10452 14473 10455
rect 14139 10424 14473 10452
rect 14139 10421 14151 10424
rect 14093 10415 14151 10421
rect 14461 10421 14473 10424
rect 14507 10421 14519 10455
rect 14461 10415 14519 10421
rect 14550 10412 14556 10464
rect 14608 10452 14614 10464
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 14608 10424 14657 10452
rect 14608 10412 14614 10424
rect 14645 10421 14657 10424
rect 14691 10421 14703 10455
rect 14645 10415 14703 10421
rect 15381 10455 15439 10461
rect 15381 10421 15393 10455
rect 15427 10452 15439 10455
rect 15562 10452 15568 10464
rect 15427 10424 15568 10452
rect 15427 10421 15439 10424
rect 15381 10415 15439 10421
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 16114 10452 16120 10464
rect 16075 10424 16120 10452
rect 16114 10412 16120 10424
rect 16172 10412 16178 10464
rect 16206 10412 16212 10464
rect 16264 10452 16270 10464
rect 18782 10452 18788 10464
rect 16264 10424 18788 10452
rect 16264 10412 16270 10424
rect 18782 10412 18788 10424
rect 18840 10412 18846 10464
rect 18877 10455 18935 10461
rect 18877 10421 18889 10455
rect 18923 10452 18935 10455
rect 19245 10455 19303 10461
rect 19245 10452 19257 10455
rect 18923 10424 19257 10452
rect 18923 10421 18935 10424
rect 18877 10415 18935 10421
rect 19245 10421 19257 10424
rect 19291 10421 19303 10455
rect 19426 10452 19432 10464
rect 19387 10424 19432 10452
rect 19245 10415 19303 10421
rect 19426 10412 19432 10424
rect 19484 10412 19490 10464
rect 19536 10452 19564 10492
rect 19797 10489 19809 10523
rect 19843 10520 19855 10523
rect 20070 10520 20076 10532
rect 19843 10492 20076 10520
rect 19843 10489 19855 10492
rect 19797 10483 19855 10489
rect 20070 10480 20076 10492
rect 20128 10480 20134 10532
rect 20714 10520 20720 10532
rect 20675 10492 20720 10520
rect 20714 10480 20720 10492
rect 20772 10480 20778 10532
rect 19889 10455 19947 10461
rect 19889 10452 19901 10455
rect 19536 10424 19901 10452
rect 19889 10421 19901 10424
rect 19935 10421 19947 10455
rect 19889 10415 19947 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 2225 10251 2283 10257
rect 2225 10217 2237 10251
rect 2271 10248 2283 10251
rect 3881 10251 3939 10257
rect 3881 10248 3893 10251
rect 2271 10220 3893 10248
rect 2271 10217 2283 10220
rect 2225 10211 2283 10217
rect 3881 10217 3893 10220
rect 3927 10217 3939 10251
rect 4062 10248 4068 10260
rect 4023 10220 4068 10248
rect 3881 10211 3939 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 5077 10251 5135 10257
rect 5077 10248 5089 10251
rect 4212 10220 5089 10248
rect 4212 10208 4218 10220
rect 5077 10217 5089 10220
rect 5123 10248 5135 10251
rect 5353 10251 5411 10257
rect 5353 10248 5365 10251
rect 5123 10220 5365 10248
rect 5123 10217 5135 10220
rect 5077 10211 5135 10217
rect 5353 10217 5365 10220
rect 5399 10217 5411 10251
rect 5534 10248 5540 10260
rect 5353 10211 5411 10217
rect 5460 10220 5540 10248
rect 1397 10183 1455 10189
rect 1397 10149 1409 10183
rect 1443 10180 1455 10183
rect 3050 10180 3056 10192
rect 1443 10152 3056 10180
rect 1443 10149 1455 10152
rect 1397 10143 1455 10149
rect 3050 10140 3056 10152
rect 3108 10140 3114 10192
rect 4614 10140 4620 10192
rect 4672 10180 4678 10192
rect 5460 10180 5488 10220
rect 5534 10208 5540 10220
rect 5592 10248 5598 10260
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 5592 10220 6837 10248
rect 5592 10208 5598 10220
rect 6825 10217 6837 10220
rect 6871 10217 6883 10251
rect 7466 10248 7472 10260
rect 7427 10220 7472 10248
rect 6825 10211 6883 10217
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 9306 10248 9312 10260
rect 9267 10220 9312 10248
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 9677 10251 9735 10257
rect 9677 10248 9689 10251
rect 9640 10220 9689 10248
rect 9640 10208 9646 10220
rect 9677 10217 9689 10220
rect 9723 10217 9735 10251
rect 9677 10211 9735 10217
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10183 10220 12756 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 6454 10180 6460 10192
rect 4672 10152 5488 10180
rect 5552 10152 6460 10180
rect 4672 10140 4678 10152
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10112 2927 10115
rect 3326 10112 3332 10124
rect 2915 10084 3332 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 3513 10115 3571 10121
rect 3513 10081 3525 10115
rect 3559 10112 3571 10115
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 3559 10084 4445 10112
rect 3559 10081 3571 10084
rect 3513 10075 3571 10081
rect 4433 10081 4445 10084
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 4525 10115 4583 10121
rect 4525 10081 4537 10115
rect 4571 10112 4583 10115
rect 4706 10112 4712 10124
rect 4571 10084 4712 10112
rect 4571 10081 4583 10084
rect 4525 10075 4583 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 5261 10115 5319 10121
rect 5261 10081 5273 10115
rect 5307 10081 5319 10115
rect 5261 10075 5319 10081
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 5399 10084 5457 10112
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 5445 10081 5457 10084
rect 5491 10081 5503 10115
rect 5445 10075 5503 10081
rect 2314 10044 2320 10056
rect 2275 10016 2320 10044
rect 2314 10004 2320 10016
rect 2372 10004 2378 10056
rect 2498 10044 2504 10056
rect 2459 10016 2504 10044
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4338 10044 4344 10056
rect 4212 10016 4344 10044
rect 4212 10004 4218 10016
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 4614 10044 4620 10056
rect 4575 10016 4620 10044
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 3053 9979 3111 9985
rect 3053 9945 3065 9979
rect 3099 9976 3111 9979
rect 3142 9976 3148 9988
rect 3099 9948 3148 9976
rect 3099 9945 3111 9948
rect 3053 9939 3111 9945
rect 3142 9936 3148 9948
rect 3200 9936 3206 9988
rect 3970 9936 3976 9988
rect 4028 9976 4034 9988
rect 5276 9976 5304 10075
rect 5552 10044 5580 10152
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 12618 10180 12624 10192
rect 6564 10152 12624 10180
rect 5712 10115 5770 10121
rect 5712 10081 5724 10115
rect 5758 10112 5770 10115
rect 5994 10112 6000 10124
rect 5758 10084 6000 10112
rect 5758 10081 5770 10084
rect 5712 10075 5770 10081
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 5460 10016 5580 10044
rect 5460 9976 5488 10016
rect 4028 9948 5212 9976
rect 5276 9948 5488 9976
rect 4028 9936 4034 9948
rect 3881 9911 3939 9917
rect 3881 9877 3893 9911
rect 3927 9908 3939 9911
rect 5074 9908 5080 9920
rect 3927 9880 5080 9908
rect 3927 9877 3939 9880
rect 3881 9871 3939 9877
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 5184 9908 5212 9948
rect 6564 9908 6592 10152
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 12728 10180 12756 10220
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 12860 10220 12909 10248
rect 12860 10208 12866 10220
rect 12897 10217 12909 10220
rect 12943 10217 12955 10251
rect 13354 10248 13360 10260
rect 13315 10220 13360 10248
rect 12897 10211 12955 10217
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 14645 10251 14703 10257
rect 14645 10217 14657 10251
rect 14691 10248 14703 10251
rect 16114 10248 16120 10260
rect 14691 10220 16120 10248
rect 14691 10217 14703 10220
rect 14645 10211 14703 10217
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 16209 10251 16267 10257
rect 16209 10217 16221 10251
rect 16255 10248 16267 10251
rect 17954 10248 17960 10260
rect 16255 10220 17960 10248
rect 16255 10217 16267 10220
rect 16209 10211 16267 10217
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 18138 10248 18144 10260
rect 18099 10220 18144 10248
rect 18138 10208 18144 10220
rect 18196 10208 18202 10260
rect 18966 10208 18972 10260
rect 19024 10248 19030 10260
rect 19024 10220 19257 10248
rect 19024 10208 19030 10220
rect 13722 10180 13728 10192
rect 12728 10152 13728 10180
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 14553 10183 14611 10189
rect 14553 10149 14565 10183
rect 14599 10180 14611 10183
rect 16390 10180 16396 10192
rect 14599 10152 16396 10180
rect 14599 10149 14611 10152
rect 14553 10143 14611 10149
rect 16390 10140 16396 10152
rect 16448 10140 16454 10192
rect 17310 10140 17316 10192
rect 17368 10180 17374 10192
rect 19229 10180 19257 10220
rect 20070 10208 20076 10260
rect 20128 10248 20134 10260
rect 20165 10251 20223 10257
rect 20165 10248 20177 10251
rect 20128 10220 20177 10248
rect 20128 10208 20134 10220
rect 20165 10217 20177 10220
rect 20211 10248 20223 10251
rect 20254 10248 20260 10260
rect 20211 10220 20260 10248
rect 20211 10217 20223 10220
rect 20165 10211 20223 10217
rect 20254 10208 20260 10220
rect 20312 10248 20318 10260
rect 20806 10248 20812 10260
rect 20312 10220 20812 10248
rect 20312 10208 20318 10220
rect 20806 10208 20812 10220
rect 20864 10208 20870 10260
rect 19610 10180 19616 10192
rect 17368 10152 18920 10180
rect 17368 10140 17374 10152
rect 7558 10072 7564 10124
rect 7616 10112 7622 10124
rect 8185 10115 8243 10121
rect 8185 10112 8197 10115
rect 7616 10084 8197 10112
rect 7616 10072 7622 10084
rect 8185 10081 8197 10084
rect 8231 10112 8243 10115
rect 9122 10112 9128 10124
rect 8231 10084 9128 10112
rect 8231 10081 8243 10084
rect 8185 10075 8243 10081
rect 9122 10072 9128 10084
rect 9180 10072 9186 10124
rect 10045 10115 10103 10121
rect 10045 10081 10057 10115
rect 10091 10112 10103 10115
rect 10318 10112 10324 10124
rect 10091 10084 10324 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 11514 10121 11520 10124
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 11112 10084 11253 10112
rect 11112 10072 11118 10084
rect 11241 10081 11253 10084
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 11497 10115 11520 10121
rect 11497 10081 11509 10115
rect 11497 10075 11520 10081
rect 11514 10072 11520 10075
rect 11572 10072 11578 10124
rect 13262 10112 13268 10124
rect 13223 10084 13268 10112
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13630 10072 13636 10124
rect 13688 10112 13694 10124
rect 15010 10112 15016 10124
rect 13688 10084 15016 10112
rect 13688 10072 13694 10084
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 15286 10072 15292 10124
rect 15344 10112 15350 10124
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 15344 10084 15669 10112
rect 15344 10072 15350 10084
rect 15657 10081 15669 10084
rect 15703 10081 15715 10115
rect 16206 10112 16212 10124
rect 15657 10075 15715 10081
rect 15948 10084 16212 10112
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 5184 9880 6592 9908
rect 7944 9908 7972 10007
rect 9030 10004 9036 10056
rect 9088 10044 9094 10056
rect 10229 10047 10287 10053
rect 10229 10044 10241 10047
rect 9088 10016 10241 10044
rect 9088 10004 9094 10016
rect 10229 10013 10241 10016
rect 10275 10013 10287 10047
rect 13538 10044 13544 10056
rect 13499 10016 13544 10044
rect 10229 10007 10287 10013
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 14829 10047 14887 10053
rect 14829 10013 14841 10047
rect 14875 10044 14887 10047
rect 15102 10044 15108 10056
rect 14875 10016 15108 10044
rect 14875 10013 14887 10016
rect 14829 10007 14887 10013
rect 15102 10004 15108 10016
rect 15160 10004 15166 10056
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15948 10053 15976 10084
rect 16206 10072 16212 10084
rect 16264 10112 16270 10124
rect 16557 10115 16615 10121
rect 16557 10112 16569 10115
rect 16264 10084 16569 10112
rect 16264 10072 16270 10084
rect 16557 10081 16569 10084
rect 16603 10081 16615 10115
rect 16557 10075 16615 10081
rect 17957 10115 18015 10121
rect 17957 10081 17969 10115
rect 18003 10112 18015 10115
rect 18414 10112 18420 10124
rect 18003 10084 18420 10112
rect 18003 10081 18015 10084
rect 17957 10075 18015 10081
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 18892 10121 18920 10152
rect 18984 10152 19196 10180
rect 19229 10152 19616 10180
rect 18984 10121 19012 10152
rect 18877 10115 18935 10121
rect 18877 10081 18889 10115
rect 18923 10081 18935 10115
rect 18877 10075 18935 10081
rect 18969 10115 19027 10121
rect 18969 10081 18981 10115
rect 19015 10081 19027 10115
rect 19168 10112 19196 10152
rect 19610 10140 19616 10152
rect 19668 10140 19674 10192
rect 19334 10112 19340 10124
rect 19168 10084 19340 10112
rect 18969 10075 19027 10081
rect 15749 10047 15807 10053
rect 15749 10044 15761 10047
rect 15252 10016 15761 10044
rect 15252 10004 15258 10016
rect 15749 10013 15761 10016
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10013 15991 10047
rect 16298 10044 16304 10056
rect 16259 10016 16304 10044
rect 15933 10007 15991 10013
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 18690 10044 18696 10056
rect 17328 10016 18696 10044
rect 11238 9936 11244 9988
rect 11296 9936 11302 9988
rect 12250 9936 12256 9988
rect 12308 9976 12314 9988
rect 16209 9979 16267 9985
rect 16209 9976 16221 9979
rect 12308 9948 16221 9976
rect 12308 9936 12314 9948
rect 16209 9945 16221 9948
rect 16255 9945 16267 9979
rect 16209 9939 16267 9945
rect 8570 9908 8576 9920
rect 7944 9880 8576 9908
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 11256 9908 11284 9936
rect 8720 9880 11284 9908
rect 8720 9868 8726 9880
rect 11606 9868 11612 9920
rect 11664 9908 11670 9920
rect 12342 9908 12348 9920
rect 11664 9880 12348 9908
rect 11664 9868 11670 9880
rect 12342 9868 12348 9880
rect 12400 9908 12406 9920
rect 12621 9911 12679 9917
rect 12621 9908 12633 9911
rect 12400 9880 12633 9908
rect 12400 9868 12406 9880
rect 12621 9877 12633 9880
rect 12667 9877 12679 9911
rect 14182 9908 14188 9920
rect 14143 9880 14188 9908
rect 12621 9871 12679 9877
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 15289 9911 15347 9917
rect 15289 9877 15301 9911
rect 15335 9908 15347 9911
rect 17328 9908 17356 10016
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 18892 9988 18920 10075
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 19978 10072 19984 10124
rect 20036 10112 20042 10124
rect 20073 10115 20131 10121
rect 20073 10112 20085 10115
rect 20036 10084 20085 10112
rect 20036 10072 20042 10084
rect 20073 10081 20085 10084
rect 20119 10081 20131 10115
rect 20073 10075 20131 10081
rect 19153 10047 19211 10053
rect 19153 10013 19165 10047
rect 19199 10044 19211 10047
rect 19518 10044 19524 10056
rect 19199 10016 19524 10044
rect 19199 10013 19211 10016
rect 19153 10007 19211 10013
rect 19518 10004 19524 10016
rect 19576 10004 19582 10056
rect 20346 10044 20352 10056
rect 20307 10016 20352 10044
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 17678 9976 17684 9988
rect 17639 9948 17684 9976
rect 17678 9936 17684 9948
rect 17736 9936 17742 9988
rect 18874 9936 18880 9988
rect 18932 9936 18938 9988
rect 18506 9908 18512 9920
rect 15335 9880 17356 9908
rect 18467 9880 18512 9908
rect 15335 9877 15347 9880
rect 15289 9871 15347 9877
rect 18506 9868 18512 9880
rect 18564 9868 18570 9920
rect 19705 9911 19763 9917
rect 19705 9877 19717 9911
rect 19751 9908 19763 9911
rect 20070 9908 20076 9920
rect 19751 9880 20076 9908
rect 19751 9877 19763 9880
rect 19705 9871 19763 9877
rect 20070 9868 20076 9880
rect 20128 9868 20134 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 2314 9664 2320 9716
rect 2372 9704 2378 9716
rect 6086 9704 6092 9716
rect 2372 9676 6092 9704
rect 2372 9664 2378 9676
rect 6086 9664 6092 9676
rect 6144 9704 6150 9716
rect 6638 9704 6644 9716
rect 6144 9676 6644 9704
rect 6144 9664 6150 9676
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 8570 9704 8576 9716
rect 7576 9676 8576 9704
rect 4065 9639 4123 9645
rect 4065 9605 4077 9639
rect 4111 9636 4123 9639
rect 4111 9608 6040 9636
rect 4111 9605 4123 9608
rect 4065 9599 4123 9605
rect 6012 9580 6040 9608
rect 1578 9528 1584 9580
rect 1636 9568 1642 9580
rect 1949 9571 2007 9577
rect 1949 9568 1961 9571
rect 1636 9540 1961 9568
rect 1636 9528 1642 9540
rect 1949 9537 1961 9540
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 3786 9528 3792 9580
rect 3844 9568 3850 9580
rect 4985 9571 5043 9577
rect 3844 9540 4936 9568
rect 3844 9528 3850 9540
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9500 1823 9503
rect 2222 9500 2228 9512
rect 1811 9472 2228 9500
rect 1811 9469 1823 9472
rect 1765 9463 1823 9469
rect 2222 9460 2228 9472
rect 2280 9460 2286 9512
rect 2685 9503 2743 9509
rect 2685 9469 2697 9503
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9500 4767 9503
rect 4798 9500 4804 9512
rect 4755 9472 4804 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 1578 9392 1584 9444
rect 1636 9432 1642 9444
rect 2700 9432 2728 9463
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 4908 9500 4936 9540
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5534 9568 5540 9580
rect 5031 9540 5540 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 5994 9568 6000 9580
rect 5955 9540 6000 9568
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 7576 9577 7604 9676
rect 8570 9664 8576 9676
rect 8628 9664 8634 9716
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 11790 9704 11796 9716
rect 10744 9676 11796 9704
rect 10744 9664 10750 9676
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 14182 9664 14188 9716
rect 14240 9704 14246 9716
rect 16206 9704 16212 9716
rect 14240 9676 16068 9704
rect 16167 9676 16212 9704
rect 14240 9664 14246 9676
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 16040 9636 16068 9676
rect 16206 9664 16212 9676
rect 16264 9664 16270 9716
rect 17218 9704 17224 9716
rect 16316 9676 17224 9704
rect 16316 9636 16344 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 17402 9664 17408 9716
rect 17460 9704 17466 9716
rect 20162 9704 20168 9716
rect 17460 9676 20168 9704
rect 17460 9664 17466 9676
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 12768 9608 13768 9636
rect 16040 9608 16344 9636
rect 12768 9596 12774 9608
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 8570 9528 8576 9580
rect 8628 9568 8634 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 8628 9540 9965 9568
rect 8628 9528 8634 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 13078 9568 13084 9580
rect 13039 9540 13084 9568
rect 9953 9531 10011 9537
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 13262 9528 13268 9580
rect 13320 9568 13326 9580
rect 13449 9571 13507 9577
rect 13449 9568 13461 9571
rect 13320 9540 13461 9568
rect 13320 9528 13326 9540
rect 13449 9537 13461 9540
rect 13495 9537 13507 9571
rect 13449 9531 13507 9537
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 4908 9472 5825 9500
rect 5813 9469 5825 9472
rect 5859 9500 5871 9503
rect 7374 9500 7380 9512
rect 5859 9472 7380 9500
rect 5859 9469 5871 9472
rect 5813 9463 5871 9469
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 7817 9503 7875 9509
rect 7817 9500 7829 9503
rect 7708 9472 7829 9500
rect 7708 9460 7714 9472
rect 7817 9469 7829 9472
rect 7863 9469 7875 9503
rect 7817 9463 7875 9469
rect 8386 9460 8392 9512
rect 8444 9500 8450 9512
rect 9582 9500 9588 9512
rect 8444 9472 9588 9500
rect 8444 9460 8450 9472
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 10220 9503 10278 9509
rect 10220 9469 10232 9503
rect 10266 9500 10278 9503
rect 11606 9500 11612 9512
rect 10266 9472 11612 9500
rect 10266 9469 10278 9472
rect 10220 9463 10278 9469
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 13630 9500 13636 9512
rect 13096 9472 13636 9500
rect 1636 9404 2728 9432
rect 1636 9392 1642 9404
rect 2866 9392 2872 9444
rect 2924 9441 2930 9444
rect 2924 9435 2988 9441
rect 2924 9401 2942 9435
rect 2976 9401 2988 9435
rect 2924 9395 2988 9401
rect 2924 9392 2930 9395
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 11514 9432 11520 9444
rect 4120 9404 11520 9432
rect 4120 9392 4126 9404
rect 11514 9392 11520 9404
rect 11572 9392 11578 9444
rect 11790 9392 11796 9444
rect 11848 9432 11854 9444
rect 13096 9432 13124 9472
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 13740 9500 13768 9608
rect 16390 9596 16396 9648
rect 16448 9636 16454 9648
rect 18141 9639 18199 9645
rect 18141 9636 18153 9639
rect 16448 9608 18153 9636
rect 16448 9596 16454 9608
rect 18141 9605 18153 9608
rect 18187 9605 18199 9639
rect 18141 9599 18199 9605
rect 18506 9596 18512 9648
rect 18564 9636 18570 9648
rect 18564 9608 18644 9636
rect 18564 9596 18570 9608
rect 14550 9528 14556 9580
rect 14608 9568 14614 9580
rect 14829 9571 14887 9577
rect 14829 9568 14841 9571
rect 14608 9540 14841 9568
rect 14608 9528 14614 9540
rect 14829 9537 14841 9540
rect 14875 9537 14887 9571
rect 14829 9531 14887 9537
rect 16942 9528 16948 9580
rect 17000 9568 17006 9580
rect 18616 9577 18644 9608
rect 18690 9596 18696 9648
rect 18748 9636 18754 9648
rect 19702 9636 19708 9648
rect 18748 9608 19708 9636
rect 18748 9596 18754 9608
rect 19702 9596 19708 9608
rect 19760 9596 19766 9648
rect 20254 9596 20260 9648
rect 20312 9636 20318 9648
rect 21358 9636 21364 9648
rect 20312 9608 21364 9636
rect 20312 9596 20318 9608
rect 21358 9596 21364 9608
rect 21416 9596 21422 9648
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 17000 9540 17049 9568
rect 17000 9528 17006 9540
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 18601 9571 18659 9577
rect 18601 9537 18613 9571
rect 18647 9537 18659 9571
rect 18601 9531 18659 9537
rect 18785 9571 18843 9577
rect 18785 9537 18797 9571
rect 18831 9568 18843 9571
rect 18966 9568 18972 9580
rect 18831 9540 18972 9568
rect 18831 9537 18843 9540
rect 18785 9531 18843 9537
rect 18966 9528 18972 9540
rect 19024 9528 19030 9580
rect 19797 9571 19855 9577
rect 19797 9537 19809 9571
rect 19843 9568 19855 9571
rect 19886 9568 19892 9580
rect 19843 9540 19892 9568
rect 19843 9537 19855 9540
rect 19797 9531 19855 9537
rect 19886 9528 19892 9540
rect 19944 9528 19950 9580
rect 20346 9528 20352 9580
rect 20404 9568 20410 9580
rect 20717 9571 20775 9577
rect 20717 9568 20729 9571
rect 20404 9540 20729 9568
rect 20404 9528 20410 9540
rect 20717 9537 20729 9540
rect 20763 9537 20775 9571
rect 20717 9531 20775 9537
rect 18690 9500 18696 9512
rect 13740 9472 18696 9500
rect 18690 9460 18696 9472
rect 18748 9500 18754 9512
rect 19334 9500 19340 9512
rect 18748 9472 19340 9500
rect 18748 9460 18754 9472
rect 19334 9460 19340 9472
rect 19392 9460 19398 9512
rect 20162 9460 20168 9512
rect 20220 9460 20226 9512
rect 20622 9500 20628 9512
rect 20583 9472 20628 9500
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 11848 9404 13124 9432
rect 11848 9392 11854 9404
rect 15010 9392 15016 9444
rect 15068 9441 15074 9444
rect 15068 9435 15132 9441
rect 15068 9401 15086 9435
rect 15120 9401 15132 9435
rect 16853 9435 16911 9441
rect 16853 9432 16865 9435
rect 15068 9395 15132 9401
rect 15764 9404 16865 9432
rect 15068 9392 15074 9395
rect 4246 9324 4252 9376
rect 4304 9364 4310 9376
rect 4341 9367 4399 9373
rect 4341 9364 4353 9367
rect 4304 9336 4353 9364
rect 4304 9324 4310 9336
rect 4341 9333 4353 9336
rect 4387 9333 4399 9367
rect 4341 9327 4399 9333
rect 4801 9367 4859 9373
rect 4801 9333 4813 9367
rect 4847 9364 4859 9367
rect 5353 9367 5411 9373
rect 5353 9364 5365 9367
rect 4847 9336 5365 9364
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 5353 9333 5365 9336
rect 5399 9333 5411 9367
rect 5718 9364 5724 9376
rect 5679 9336 5724 9364
rect 5353 9327 5411 9333
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 8941 9367 8999 9373
rect 8941 9364 8953 9367
rect 6788 9336 8953 9364
rect 6788 9324 6794 9336
rect 8941 9333 8953 9336
rect 8987 9364 8999 9367
rect 9950 9364 9956 9376
rect 8987 9336 9956 9364
rect 8987 9333 8999 9336
rect 8941 9327 8999 9333
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11333 9367 11391 9373
rect 11333 9364 11345 9367
rect 11020 9336 11345 9364
rect 11020 9324 11026 9336
rect 11333 9333 11345 9336
rect 11379 9333 11391 9367
rect 11333 9327 11391 9333
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12526 9364 12532 9376
rect 12483 9336 12532 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 12802 9364 12808 9376
rect 12763 9336 12808 9364
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 14369 9367 14427 9373
rect 12952 9336 12997 9364
rect 12952 9324 12958 9336
rect 14369 9333 14381 9367
rect 14415 9364 14427 9367
rect 15764 9364 15792 9404
rect 16853 9401 16865 9404
rect 16899 9401 16911 9435
rect 16853 9395 16911 9401
rect 18509 9435 18567 9441
rect 18509 9401 18521 9435
rect 18555 9432 18567 9435
rect 19426 9432 19432 9444
rect 18555 9404 19432 9432
rect 18555 9401 18567 9404
rect 18509 9395 18567 9401
rect 19426 9392 19432 9404
rect 19484 9392 19490 9444
rect 20180 9432 20208 9460
rect 20180 9404 20668 9432
rect 20640 9376 20668 9404
rect 16482 9364 16488 9376
rect 14415 9336 15792 9364
rect 16443 9336 16488 9364
rect 14415 9333 14427 9336
rect 14369 9327 14427 9333
rect 16482 9324 16488 9336
rect 16540 9324 16546 9376
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 16945 9367 17003 9373
rect 16945 9364 16957 9367
rect 16724 9336 16957 9364
rect 16724 9324 16730 9336
rect 16945 9333 16957 9336
rect 16991 9333 17003 9367
rect 16945 9327 17003 9333
rect 19153 9367 19211 9373
rect 19153 9333 19165 9367
rect 19199 9364 19211 9367
rect 19334 9364 19340 9376
rect 19199 9336 19340 9364
rect 19199 9333 19211 9336
rect 19153 9327 19211 9333
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 19518 9364 19524 9376
rect 19479 9336 19524 9364
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 19613 9367 19671 9373
rect 19613 9333 19625 9367
rect 19659 9364 19671 9367
rect 19702 9364 19708 9376
rect 19659 9336 19708 9364
rect 19659 9333 19671 9336
rect 19613 9327 19671 9333
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 20162 9364 20168 9376
rect 20123 9336 20168 9364
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 20530 9364 20536 9376
rect 20491 9336 20536 9364
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 20622 9324 20628 9376
rect 20680 9324 20686 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 2222 9160 2228 9172
rect 2183 9132 2228 9160
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 4433 9163 4491 9169
rect 4433 9129 4445 9163
rect 4479 9160 4491 9163
rect 4706 9160 4712 9172
rect 4479 9132 4712 9160
rect 4479 9129 4491 9132
rect 4433 9123 4491 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 4801 9163 4859 9169
rect 4801 9129 4813 9163
rect 4847 9160 4859 9163
rect 4890 9160 4896 9172
rect 4847 9132 4896 9160
rect 4847 9129 4859 9132
rect 4801 9123 4859 9129
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 5442 9160 5448 9172
rect 5403 9132 5448 9160
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 7101 9163 7159 9169
rect 7101 9129 7113 9163
rect 7147 9160 7159 9163
rect 7742 9160 7748 9172
rect 7147 9132 7748 9160
rect 7147 9129 7159 9132
rect 7101 9123 7159 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8113 9163 8171 9169
rect 8113 9129 8125 9163
rect 8159 9160 8171 9163
rect 8202 9160 8208 9172
rect 8159 9132 8208 9160
rect 8159 9129 8171 9132
rect 8113 9123 8171 9129
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 9858 9160 9864 9172
rect 8527 9132 9864 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 9858 9120 9864 9132
rect 9916 9120 9922 9172
rect 10134 9160 10140 9172
rect 10095 9132 10140 9160
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10781 9163 10839 9169
rect 10781 9129 10793 9163
rect 10827 9160 10839 9163
rect 12894 9160 12900 9172
rect 10827 9132 12900 9160
rect 10827 9129 10839 9132
rect 10781 9123 10839 9129
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 13078 9120 13084 9172
rect 13136 9160 13142 9172
rect 13265 9163 13323 9169
rect 13265 9160 13277 9163
rect 13136 9132 13277 9160
rect 13136 9120 13142 9132
rect 13265 9129 13277 9132
rect 13311 9129 13323 9163
rect 13265 9123 13323 9129
rect 14921 9163 14979 9169
rect 14921 9129 14933 9163
rect 14967 9160 14979 9163
rect 15010 9160 15016 9172
rect 14967 9132 15016 9160
rect 14967 9129 14979 9132
rect 14921 9123 14979 9129
rect 1765 9095 1823 9101
rect 1765 9061 1777 9095
rect 1811 9092 1823 9095
rect 3326 9092 3332 9104
rect 1811 9064 3332 9092
rect 1811 9061 1823 9064
rect 1765 9055 1823 9061
rect 3326 9052 3332 9064
rect 3384 9052 3390 9104
rect 4246 9052 4252 9104
rect 4304 9092 4310 9104
rect 5074 9092 5080 9104
rect 4304 9064 5080 9092
rect 4304 9052 4310 9064
rect 5074 9052 5080 9064
rect 5132 9052 5138 9104
rect 5350 9052 5356 9104
rect 5408 9092 5414 9104
rect 5905 9095 5963 9101
rect 5905 9092 5917 9095
rect 5408 9064 5917 9092
rect 5408 9052 5414 9064
rect 5905 9061 5917 9064
rect 5951 9061 5963 9095
rect 5905 9055 5963 9061
rect 7374 9052 7380 9104
rect 7432 9092 7438 9104
rect 7561 9095 7619 9101
rect 7561 9092 7573 9095
rect 7432 9064 7573 9092
rect 7432 9052 7438 9064
rect 7561 9061 7573 9064
rect 7607 9061 7619 9095
rect 7561 9055 7619 9061
rect 8938 9052 8944 9104
rect 8996 9092 9002 9104
rect 10045 9095 10103 9101
rect 10045 9092 10057 9095
rect 8996 9064 10057 9092
rect 8996 9052 9002 9064
rect 10045 9061 10057 9064
rect 10091 9061 10103 9095
rect 10045 9055 10103 9061
rect 10870 9052 10876 9104
rect 10928 9092 10934 9104
rect 11241 9095 11299 9101
rect 11241 9092 11253 9095
rect 10928 9064 11253 9092
rect 10928 9052 10934 9064
rect 11241 9061 11253 9064
rect 11287 9061 11299 9095
rect 13280 9092 13308 9123
rect 15010 9120 15016 9132
rect 15068 9120 15074 9172
rect 15286 9160 15292 9172
rect 15247 9132 15292 9160
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15657 9163 15715 9169
rect 15657 9129 15669 9163
rect 15703 9160 15715 9163
rect 16482 9160 16488 9172
rect 15703 9132 16488 9160
rect 15703 9129 15715 9132
rect 15657 9123 15715 9129
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 16761 9163 16819 9169
rect 16761 9129 16773 9163
rect 16807 9160 16819 9163
rect 17770 9160 17776 9172
rect 16807 9132 17776 9160
rect 16807 9129 16819 9132
rect 16761 9123 16819 9129
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 20530 9120 20536 9172
rect 20588 9160 20594 9172
rect 20901 9163 20959 9169
rect 20901 9160 20913 9163
rect 20588 9132 20913 9160
rect 20588 9120 20594 9132
rect 20901 9129 20913 9132
rect 20947 9129 20959 9163
rect 20901 9123 20959 9129
rect 13808 9095 13866 9101
rect 13808 9092 13820 9095
rect 13280 9064 13820 9092
rect 11241 9055 11299 9061
rect 13808 9061 13820 9064
rect 13854 9092 13866 9095
rect 16942 9092 16948 9104
rect 13854 9064 16948 9092
rect 13854 9061 13866 9064
rect 13808 9055 13866 9061
rect 16942 9052 16948 9064
rect 17000 9052 17006 9104
rect 17862 9092 17868 9104
rect 17696 9064 17868 9092
rect 1489 9027 1547 9033
rect 1489 8993 1501 9027
rect 1535 8993 1547 9027
rect 2590 9024 2596 9036
rect 2551 8996 2596 9024
rect 1489 8987 1547 8993
rect 1504 8820 1532 8987
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 5092 9024 5120 9052
rect 5718 9024 5724 9036
rect 5092 8996 5724 9024
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 9024 5871 9027
rect 6178 9024 6184 9036
rect 5859 8996 6184 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 6178 8984 6184 8996
rect 6236 9024 6242 9036
rect 6546 9024 6552 9036
rect 6236 8996 6552 9024
rect 6236 8984 6242 8996
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 7282 8984 7288 9036
rect 7340 9024 7346 9036
rect 7469 9027 7527 9033
rect 7469 9024 7481 9027
rect 7340 8996 7481 9024
rect 7340 8984 7346 8996
rect 7469 8993 7481 8996
rect 7515 8993 7527 9027
rect 7926 9024 7932 9036
rect 7469 8987 7527 8993
rect 7576 8996 7932 9024
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8925 2743 8959
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2685 8919 2743 8925
rect 2700 8888 2728 8919
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 4798 8956 4804 8968
rect 3752 8928 4804 8956
rect 3752 8916 3758 8928
rect 4798 8916 4804 8928
rect 4856 8956 4862 8968
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 4856 8928 4905 8956
rect 4856 8916 4862 8928
rect 4893 8925 4905 8928
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5994 8956 6000 8968
rect 5123 8928 6000 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5994 8916 6000 8928
rect 6052 8956 6058 8968
rect 6089 8959 6147 8965
rect 6089 8956 6101 8959
rect 6052 8928 6101 8956
rect 6052 8916 6058 8928
rect 6089 8925 6101 8928
rect 6135 8925 6147 8959
rect 6089 8919 6147 8925
rect 3142 8888 3148 8900
rect 2700 8860 3148 8888
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 6104 8888 6132 8919
rect 7190 8916 7196 8968
rect 7248 8956 7254 8968
rect 7576 8956 7604 8996
rect 7926 8984 7932 8996
rect 7984 8984 7990 9036
rect 8573 9027 8631 9033
rect 8573 8993 8585 9027
rect 8619 9024 8631 9027
rect 9490 9024 9496 9036
rect 8619 8996 9496 9024
rect 8619 8993 8631 8996
rect 8573 8987 8631 8993
rect 9490 8984 9496 8996
rect 9548 8984 9554 9036
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 10008 8996 10272 9024
rect 10008 8984 10014 8996
rect 7248 8928 7604 8956
rect 7248 8916 7254 8928
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 8757 8959 8815 8965
rect 7708 8928 7753 8956
rect 7708 8916 7714 8928
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 9030 8956 9036 8968
rect 8803 8928 9036 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 8772 8888 8800 8919
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 10134 8956 10140 8968
rect 9180 8928 10140 8956
rect 9180 8916 9186 8928
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10244 8965 10272 8996
rect 10318 8984 10324 9036
rect 10376 9024 10382 9036
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 10376 8996 11161 9024
rect 10376 8984 10382 8996
rect 11149 8993 11161 8996
rect 11195 8993 11207 9027
rect 12141 9027 12199 9033
rect 12141 9024 12153 9027
rect 11149 8987 11207 8993
rect 11440 8996 12153 9024
rect 11440 8965 11468 8996
rect 12141 8993 12153 8996
rect 12187 9024 12199 9027
rect 12894 9024 12900 9036
rect 12187 8996 12900 9024
rect 12187 8993 12199 8996
rect 12141 8987 12199 8993
rect 12894 8984 12900 8996
rect 12952 8984 12958 9036
rect 13630 8984 13636 9036
rect 13688 9024 13694 9036
rect 16669 9027 16727 9033
rect 13688 8996 16620 9024
rect 13688 8984 13694 8996
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8925 11943 8959
rect 11885 8919 11943 8925
rect 13541 8959 13599 8965
rect 13541 8925 13553 8959
rect 13587 8925 13599 8959
rect 15746 8956 15752 8968
rect 15707 8928 15752 8956
rect 13541 8919 13599 8925
rect 4120 8860 5488 8888
rect 6104 8860 8800 8888
rect 9677 8891 9735 8897
rect 4120 8848 4126 8860
rect 5350 8820 5356 8832
rect 1504 8792 5356 8820
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 5460 8820 5488 8860
rect 9677 8857 9689 8891
rect 9723 8888 9735 8891
rect 10502 8888 10508 8900
rect 9723 8860 10508 8888
rect 9723 8857 9735 8860
rect 9677 8851 9735 8857
rect 10502 8848 10508 8860
rect 10560 8848 10566 8900
rect 11054 8848 11060 8900
rect 11112 8888 11118 8900
rect 11900 8888 11928 8919
rect 11112 8860 11928 8888
rect 11112 8848 11118 8860
rect 11790 8820 11796 8832
rect 5460 8792 11796 8820
rect 11790 8780 11796 8792
rect 11848 8780 11854 8832
rect 11900 8820 11928 8860
rect 12250 8820 12256 8832
rect 11900 8792 12256 8820
rect 12250 8780 12256 8792
rect 12308 8820 12314 8832
rect 13556 8820 13584 8919
rect 15746 8916 15752 8928
rect 15804 8916 15810 8968
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 15010 8848 15016 8900
rect 15068 8888 15074 8900
rect 15856 8888 15884 8919
rect 15068 8860 15884 8888
rect 15068 8848 15074 8860
rect 12308 8792 13584 8820
rect 12308 8780 12314 8792
rect 15286 8780 15292 8832
rect 15344 8820 15350 8832
rect 16301 8823 16359 8829
rect 16301 8820 16313 8823
rect 15344 8792 16313 8820
rect 15344 8780 15350 8792
rect 16301 8789 16313 8792
rect 16347 8789 16359 8823
rect 16592 8820 16620 8996
rect 16669 8993 16681 9027
rect 16715 9024 16727 9027
rect 17126 9024 17132 9036
rect 16715 8996 17132 9024
rect 16715 8993 16727 8996
rect 16669 8987 16727 8993
rect 17126 8984 17132 8996
rect 17184 9024 17190 9036
rect 17586 9024 17592 9036
rect 17184 8996 17592 9024
rect 17184 8984 17190 8996
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 16942 8956 16948 8968
rect 16903 8928 16948 8956
rect 16942 8916 16948 8928
rect 17000 8916 17006 8968
rect 16666 8848 16672 8900
rect 16724 8888 16730 8900
rect 17696 8888 17724 9064
rect 17862 9052 17868 9064
rect 17920 9052 17926 9104
rect 18500 9095 18558 9101
rect 18500 9061 18512 9095
rect 18546 9092 18558 9095
rect 19426 9092 19432 9104
rect 18546 9064 19432 9092
rect 18546 9061 18558 9064
rect 18500 9055 18558 9061
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 19610 9052 19616 9104
rect 19668 9092 19674 9104
rect 20165 9095 20223 9101
rect 20165 9092 20177 9095
rect 19668 9064 20177 9092
rect 19668 9052 19674 9064
rect 20165 9061 20177 9064
rect 20211 9061 20223 9095
rect 20165 9055 20223 9061
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 19889 9027 19947 9033
rect 19889 9024 19901 9027
rect 19392 8996 19901 9024
rect 19392 8984 19398 8996
rect 19889 8993 19901 8996
rect 19935 8993 19947 9027
rect 19889 8987 19947 8993
rect 17862 8916 17868 8968
rect 17920 8956 17926 8968
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 17920 8928 18245 8956
rect 17920 8916 17926 8928
rect 18233 8925 18245 8928
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 16724 8860 17724 8888
rect 16724 8848 16730 8860
rect 19613 8823 19671 8829
rect 19613 8820 19625 8823
rect 16592 8792 19625 8820
rect 16301 8783 16359 8789
rect 19613 8789 19625 8792
rect 19659 8820 19671 8823
rect 19886 8820 19892 8832
rect 19659 8792 19892 8820
rect 19659 8789 19671 8792
rect 19613 8783 19671 8789
rect 19886 8780 19892 8792
rect 19944 8780 19950 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2866 8616 2872 8628
rect 2827 8588 2872 8616
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 3142 8616 3148 8628
rect 3103 8588 3148 8616
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 4341 8619 4399 8625
rect 4341 8585 4353 8619
rect 4387 8616 4399 8619
rect 5350 8616 5356 8628
rect 4387 8588 4936 8616
rect 5311 8588 5356 8616
rect 4387 8585 4399 8588
rect 4341 8579 4399 8585
rect 4908 8548 4936 8588
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 10229 8619 10287 8625
rect 10229 8616 10241 8619
rect 5592 8588 10241 8616
rect 5592 8576 5598 8588
rect 10229 8585 10241 8588
rect 10275 8585 10287 8619
rect 12434 8616 12440 8628
rect 10229 8579 10287 8585
rect 10336 8588 12440 8616
rect 7561 8551 7619 8557
rect 2700 8520 3740 8548
rect 4908 8520 5856 8548
rect 2700 8424 2728 8520
rect 3712 8489 3740 8520
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8449 3755 8483
rect 4798 8480 4804 8492
rect 4759 8452 4804 8480
rect 3697 8443 3755 8449
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8480 5043 8483
rect 5626 8480 5632 8492
rect 5031 8452 5632 8480
rect 5031 8449 5043 8452
rect 4985 8443 5043 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5828 8489 5856 8520
rect 7561 8517 7573 8551
rect 7607 8517 7619 8551
rect 8389 8551 8447 8557
rect 8389 8548 8401 8551
rect 7561 8511 7619 8517
rect 8128 8520 8401 8548
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8480 6055 8483
rect 7098 8480 7104 8492
rect 6043 8452 7104 8480
rect 6043 8449 6055 8452
rect 5997 8443 6055 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 1489 8415 1547 8421
rect 1489 8381 1501 8415
rect 1535 8412 1547 8415
rect 1578 8412 1584 8424
rect 1535 8384 1584 8412
rect 1535 8381 1547 8384
rect 1489 8375 1547 8381
rect 1578 8372 1584 8384
rect 1636 8372 1642 8424
rect 1756 8415 1814 8421
rect 1756 8381 1768 8415
rect 1802 8412 1814 8415
rect 2682 8412 2688 8424
rect 1802 8384 2688 8412
rect 1802 8381 1814 8384
rect 1756 8375 1814 8381
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 3605 8415 3663 8421
rect 3605 8381 3617 8415
rect 3651 8412 3663 8415
rect 7576 8412 7604 8511
rect 8128 8489 8156 8520
rect 8389 8517 8401 8520
rect 8435 8517 8447 8551
rect 8389 8511 8447 8517
rect 9953 8551 10011 8557
rect 9953 8517 9965 8551
rect 9999 8548 10011 8551
rect 10045 8551 10103 8557
rect 10045 8548 10057 8551
rect 9999 8520 10057 8548
rect 9999 8517 10011 8520
rect 9953 8511 10011 8517
rect 10045 8517 10057 8520
rect 10091 8517 10103 8551
rect 10045 8511 10103 8517
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 8220 8452 8708 8480
rect 8220 8412 8248 8452
rect 8570 8412 8576 8424
rect 3651 8384 7604 8412
rect 7668 8384 8248 8412
rect 8531 8384 8576 8412
rect 3651 8381 3663 8384
rect 3605 8375 3663 8381
rect 4709 8347 4767 8353
rect 4709 8313 4721 8347
rect 4755 8344 4767 8347
rect 4755 8316 5120 8344
rect 4755 8313 4767 8316
rect 4709 8307 4767 8313
rect 3510 8276 3516 8288
rect 3471 8248 3516 8276
rect 3510 8236 3516 8248
rect 3568 8236 3574 8288
rect 5092 8276 5120 8316
rect 5166 8304 5172 8356
rect 5224 8344 5230 8356
rect 5721 8347 5779 8353
rect 5721 8344 5733 8347
rect 5224 8316 5733 8344
rect 5224 8304 5230 8316
rect 5721 8313 5733 8316
rect 5767 8313 5779 8347
rect 5721 8307 5779 8313
rect 6822 8304 6828 8356
rect 6880 8344 6886 8356
rect 7668 8344 7696 8384
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8680 8412 8708 8452
rect 9582 8440 9588 8492
rect 9640 8480 9646 8492
rect 10336 8480 10364 8588
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 14737 8619 14795 8625
rect 14737 8585 14749 8619
rect 14783 8616 14795 8619
rect 15194 8616 15200 8628
rect 14783 8588 15200 8616
rect 14783 8585 14795 8588
rect 14737 8579 14795 8585
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 15746 8616 15752 8628
rect 15707 8588 15752 8616
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 16945 8619 17003 8625
rect 16945 8585 16957 8619
rect 16991 8616 17003 8619
rect 19426 8616 19432 8628
rect 16991 8588 19104 8616
rect 19387 8588 19432 8616
rect 16991 8585 17003 8588
rect 16945 8579 17003 8585
rect 11241 8551 11299 8557
rect 11241 8517 11253 8551
rect 11287 8517 11299 8551
rect 12158 8548 12164 8560
rect 11241 8511 11299 8517
rect 11716 8520 12164 8548
rect 10781 8483 10839 8489
rect 10781 8480 10793 8483
rect 9640 8452 10364 8480
rect 10428 8452 10793 8480
rect 9640 8440 9646 8452
rect 10045 8415 10103 8421
rect 10045 8412 10057 8415
rect 8680 8384 10057 8412
rect 10045 8381 10057 8384
rect 10091 8412 10103 8415
rect 10428 8412 10456 8452
rect 10781 8449 10793 8452
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 10091 8384 10456 8412
rect 10597 8415 10655 8421
rect 10091 8381 10103 8384
rect 10045 8375 10103 8381
rect 10597 8381 10609 8415
rect 10643 8412 10655 8415
rect 11256 8412 11284 8511
rect 11716 8489 11744 8520
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 10643 8384 11284 8412
rect 10643 8381 10655 8384
rect 10597 8375 10655 8381
rect 7926 8344 7932 8356
rect 6880 8316 7696 8344
rect 7887 8316 7932 8344
rect 6880 8304 6886 8316
rect 7926 8304 7932 8316
rect 7984 8304 7990 8356
rect 8021 8347 8079 8353
rect 8021 8313 8033 8347
rect 8067 8344 8079 8347
rect 8478 8344 8484 8356
rect 8067 8316 8484 8344
rect 8067 8313 8079 8316
rect 8021 8307 8079 8313
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 8840 8347 8898 8353
rect 8840 8313 8852 8347
rect 8886 8344 8898 8347
rect 9674 8344 9680 8356
rect 8886 8316 9680 8344
rect 8886 8313 8898 8316
rect 8840 8307 8898 8313
rect 9674 8304 9680 8316
rect 9732 8344 9738 8356
rect 10962 8344 10968 8356
rect 9732 8316 10968 8344
rect 9732 8304 9738 8316
rect 10962 8304 10968 8316
rect 11020 8344 11026 8356
rect 11808 8344 11836 8443
rect 12250 8440 12256 8492
rect 12308 8480 12314 8492
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 12308 8452 12449 8480
rect 12308 8440 12314 8452
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 13446 8440 13452 8492
rect 13504 8480 13510 8492
rect 13504 8452 14044 8480
rect 13504 8440 13510 8452
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 14016 8412 14044 8452
rect 15010 8440 15016 8492
rect 15068 8480 15074 8492
rect 15289 8483 15347 8489
rect 15289 8480 15301 8483
rect 15068 8452 15301 8480
rect 15068 8440 15074 8452
rect 15289 8449 15301 8452
rect 15335 8449 15347 8483
rect 15289 8443 15347 8449
rect 16393 8483 16451 8489
rect 16393 8449 16405 8483
rect 16439 8480 16451 8483
rect 16942 8480 16948 8492
rect 16439 8452 16948 8480
rect 16439 8449 16451 8452
rect 16393 8443 16451 8449
rect 16942 8440 16948 8452
rect 17000 8440 17006 8492
rect 17494 8480 17500 8492
rect 17455 8452 17500 8480
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 19076 8480 19104 8588
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 19702 8616 19708 8628
rect 19663 8588 19708 8616
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 20901 8619 20959 8625
rect 20901 8585 20913 8619
rect 20947 8616 20959 8619
rect 20990 8616 20996 8628
rect 20947 8588 20996 8616
rect 20947 8585 20959 8588
rect 20901 8579 20959 8585
rect 20990 8576 20996 8588
rect 21048 8576 21054 8628
rect 19444 8548 19472 8576
rect 19978 8548 19984 8560
rect 19444 8520 19984 8548
rect 19978 8508 19984 8520
rect 20036 8548 20042 8560
rect 20036 8520 20300 8548
rect 20036 8508 20042 8520
rect 20272 8489 20300 8520
rect 20165 8483 20223 8489
rect 20165 8480 20177 8483
rect 19076 8452 20177 8480
rect 20165 8449 20177 8452
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 16117 8415 16175 8421
rect 16117 8412 16129 8415
rect 12584 8384 13860 8412
rect 14016 8384 16129 8412
rect 12584 8372 12590 8384
rect 11020 8316 11836 8344
rect 12704 8347 12762 8353
rect 11020 8304 11026 8316
rect 12704 8313 12716 8347
rect 12750 8344 12762 8347
rect 13630 8344 13636 8356
rect 12750 8316 13636 8344
rect 12750 8313 12762 8316
rect 12704 8307 12762 8313
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 13832 8344 13860 8384
rect 16117 8381 16129 8384
rect 16163 8412 16175 8415
rect 16666 8412 16672 8424
rect 16163 8384 16672 8412
rect 16163 8381 16175 8384
rect 16117 8375 16175 8381
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 17402 8412 17408 8424
rect 16868 8384 17408 8412
rect 15197 8347 15255 8353
rect 15197 8344 15209 8347
rect 13832 8316 15209 8344
rect 15197 8313 15209 8316
rect 15243 8313 15255 8347
rect 15197 8307 15255 8313
rect 15286 8304 15292 8356
rect 15344 8304 15350 8356
rect 15378 8304 15384 8356
rect 15436 8344 15442 8356
rect 16209 8347 16267 8353
rect 16209 8344 16221 8347
rect 15436 8316 16221 8344
rect 15436 8304 15442 8316
rect 16209 8313 16221 8316
rect 16255 8344 16267 8347
rect 16868 8344 16896 8384
rect 17402 8372 17408 8384
rect 17460 8372 17466 8424
rect 17862 8372 17868 8424
rect 17920 8412 17926 8424
rect 18046 8412 18052 8424
rect 17920 8384 18052 8412
rect 17920 8372 17926 8384
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 20070 8412 20076 8424
rect 20031 8384 20076 8412
rect 20070 8372 20076 8384
rect 20128 8372 20134 8424
rect 20714 8412 20720 8424
rect 20675 8384 20720 8412
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 16255 8316 16896 8344
rect 17313 8347 17371 8353
rect 16255 8313 16267 8316
rect 16209 8307 16267 8313
rect 17313 8313 17325 8347
rect 17359 8344 17371 8347
rect 17954 8344 17960 8356
rect 17359 8316 17960 8344
rect 17359 8313 17371 8316
rect 17313 8307 17371 8313
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 18322 8353 18328 8356
rect 18316 8344 18328 8353
rect 18283 8316 18328 8344
rect 18316 8307 18328 8316
rect 18380 8344 18386 8356
rect 20346 8344 20352 8356
rect 18380 8316 20352 8344
rect 18322 8304 18328 8307
rect 18380 8304 18386 8316
rect 20346 8304 20352 8316
rect 20404 8304 20410 8356
rect 5534 8276 5540 8288
rect 5092 8248 5540 8276
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 5994 8236 6000 8288
rect 6052 8276 6058 8288
rect 8389 8279 8447 8285
rect 8389 8276 8401 8279
rect 6052 8248 8401 8276
rect 6052 8236 6058 8248
rect 8389 8245 8401 8248
rect 8435 8276 8447 8279
rect 9214 8276 9220 8288
rect 8435 8248 9220 8276
rect 8435 8245 8447 8248
rect 8389 8239 8447 8245
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 10686 8276 10692 8288
rect 10647 8248 10692 8276
rect 10686 8236 10692 8248
rect 10744 8236 10750 8288
rect 11606 8276 11612 8288
rect 11567 8248 11612 8276
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 13817 8279 13875 8285
rect 13817 8276 13829 8279
rect 12952 8248 13829 8276
rect 12952 8236 12958 8248
rect 13817 8245 13829 8248
rect 13863 8245 13875 8279
rect 13817 8239 13875 8245
rect 15105 8279 15163 8285
rect 15105 8245 15117 8279
rect 15151 8276 15163 8279
rect 15304 8276 15332 8304
rect 17402 8276 17408 8288
rect 15151 8248 15332 8276
rect 17363 8248 17408 8276
rect 15151 8245 15163 8248
rect 15105 8239 15163 8245
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 19886 8236 19892 8288
rect 19944 8276 19950 8288
rect 20070 8276 20076 8288
rect 19944 8248 20076 8276
rect 19944 8236 19950 8248
rect 20070 8236 20076 8248
rect 20128 8236 20134 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 2590 8072 2596 8084
rect 2551 8044 2596 8072
rect 2590 8032 2596 8044
rect 2648 8032 2654 8084
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 3568 8044 4077 8072
rect 3568 8032 3574 8044
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 5074 8072 5080 8084
rect 4571 8044 5080 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 5994 8072 6000 8084
rect 5184 8044 6000 8072
rect 1486 7964 1492 8016
rect 1544 8004 1550 8016
rect 3053 8007 3111 8013
rect 3053 8004 3065 8007
rect 1544 7976 3065 8004
rect 1544 7964 1550 7976
rect 3053 7973 3065 7976
rect 3099 7973 3111 8007
rect 3053 7967 3111 7973
rect 2958 7936 2964 7948
rect 2919 7908 2964 7936
rect 2958 7896 2964 7908
rect 3016 7896 3022 7948
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 4706 7936 4712 7948
rect 4479 7908 4712 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 2682 7828 2688 7880
rect 2740 7868 2746 7880
rect 3145 7871 3203 7877
rect 3145 7868 3157 7871
rect 2740 7840 3157 7868
rect 2740 7828 2746 7840
rect 3145 7837 3157 7840
rect 3191 7868 3203 7871
rect 3878 7868 3884 7880
rect 3191 7840 3884 7868
rect 3191 7837 3203 7840
rect 3145 7831 3203 7837
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 3970 7828 3976 7880
rect 4028 7868 4034 7880
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 4028 7840 4629 7868
rect 4028 7828 4034 7840
rect 4617 7837 4629 7840
rect 4663 7868 4675 7871
rect 5184 7868 5212 8044
rect 5994 8032 6000 8044
rect 6052 8032 6058 8084
rect 7098 8072 7104 8084
rect 7059 8044 7104 8072
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7745 8075 7803 8081
rect 7745 8041 7757 8075
rect 7791 8072 7803 8075
rect 8570 8072 8576 8084
rect 7791 8044 8576 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 9214 8072 9220 8084
rect 9175 8044 9220 8072
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 9953 8075 10011 8081
rect 9953 8041 9965 8075
rect 9999 8072 10011 8075
rect 10686 8072 10692 8084
rect 9999 8044 10692 8072
rect 9999 8041 10011 8044
rect 9953 8035 10011 8041
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 12345 8075 12403 8081
rect 12345 8041 12357 8075
rect 12391 8072 12403 8075
rect 12802 8072 12808 8084
rect 12391 8044 12808 8072
rect 12391 8041 12403 8044
rect 12345 8035 12403 8041
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 18233 8075 18291 8081
rect 18233 8072 18245 8075
rect 17552 8044 18245 8072
rect 17552 8032 17558 8044
rect 18233 8041 18245 8044
rect 18279 8072 18291 8075
rect 18322 8072 18328 8084
rect 18279 8044 18328 8072
rect 18279 8041 18291 8044
rect 18233 8035 18291 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 19429 8075 19487 8081
rect 19429 8041 19441 8075
rect 19475 8072 19487 8075
rect 19518 8072 19524 8084
rect 19475 8044 19524 8072
rect 19475 8041 19487 8044
rect 19429 8035 19487 8041
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 19797 8075 19855 8081
rect 19797 8041 19809 8075
rect 19843 8072 19855 8075
rect 20162 8072 20168 8084
rect 19843 8044 20168 8072
rect 19843 8041 19855 8044
rect 19797 8035 19855 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 5350 7964 5356 8016
rect 5408 8004 5414 8016
rect 16022 8004 16028 8016
rect 5408 7976 16028 8004
rect 5408 7964 5414 7976
rect 16022 7964 16028 7976
rect 16080 7964 16086 8016
rect 18046 8004 18052 8016
rect 16868 7976 18052 8004
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 8110 7945 8116 7948
rect 5977 7939 6035 7945
rect 5977 7936 5989 7939
rect 5684 7908 5989 7936
rect 5684 7896 5690 7908
rect 5977 7905 5989 7908
rect 6023 7905 6035 7939
rect 5977 7899 6035 7905
rect 8104 7899 8116 7945
rect 8168 7936 8174 7948
rect 10318 7936 10324 7948
rect 8168 7908 8204 7936
rect 10279 7908 10324 7936
rect 8110 7896 8116 7899
rect 8168 7896 8174 7908
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 10413 7939 10471 7945
rect 10413 7905 10425 7939
rect 10459 7936 10471 7939
rect 10870 7936 10876 7948
rect 10459 7908 10876 7936
rect 10459 7905 10471 7908
rect 10413 7899 10471 7905
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 12710 7936 12716 7948
rect 12671 7908 12716 7936
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 16298 7896 16304 7948
rect 16356 7936 16362 7948
rect 16666 7936 16672 7948
rect 16356 7908 16672 7936
rect 16356 7896 16362 7908
rect 16666 7896 16672 7908
rect 16724 7936 16730 7948
rect 16868 7945 16896 7976
rect 18046 7964 18052 7976
rect 18104 8004 18110 8016
rect 19150 8004 19156 8016
rect 18104 7976 19156 8004
rect 18104 7964 18110 7976
rect 19150 7964 19156 7976
rect 19208 7964 19214 8016
rect 17126 7945 17132 7948
rect 16853 7939 16911 7945
rect 16853 7936 16865 7939
rect 16724 7908 16865 7936
rect 16724 7896 16730 7908
rect 16853 7905 16865 7908
rect 16899 7905 16911 7939
rect 16853 7899 16911 7905
rect 17120 7899 17132 7945
rect 17184 7936 17190 7948
rect 17184 7908 17220 7936
rect 17126 7896 17132 7899
rect 17184 7896 17190 7908
rect 4663 7840 5212 7868
rect 5721 7871 5779 7877
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 2498 7760 2504 7812
rect 2556 7800 2562 7812
rect 5736 7800 5764 7831
rect 6914 7828 6920 7880
rect 6972 7868 6978 7880
rect 7745 7871 7803 7877
rect 7745 7868 7757 7871
rect 6972 7840 7757 7868
rect 6972 7828 6978 7840
rect 7745 7837 7757 7840
rect 7791 7868 7803 7871
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7791 7840 7849 7868
rect 7791 7837 7803 7840
rect 7745 7831 7803 7837
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 10505 7871 10563 7877
rect 10505 7868 10517 7871
rect 9732 7840 10517 7868
rect 9732 7828 9738 7840
rect 10505 7837 10517 7840
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 12158 7828 12164 7880
rect 12216 7868 12222 7880
rect 12805 7871 12863 7877
rect 12805 7868 12817 7871
rect 12216 7840 12817 7868
rect 12216 7828 12222 7840
rect 12805 7837 12817 7840
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 12894 7828 12900 7880
rect 12952 7868 12958 7880
rect 19886 7868 19892 7880
rect 12952 7840 12997 7868
rect 19847 7840 19892 7868
rect 12952 7828 12958 7840
rect 19886 7828 19892 7840
rect 19944 7828 19950 7880
rect 19978 7828 19984 7880
rect 20036 7868 20042 7880
rect 20036 7840 20081 7868
rect 20036 7828 20042 7840
rect 13906 7800 13912 7812
rect 2556 7772 5764 7800
rect 8772 7772 13912 7800
rect 2556 7760 2562 7772
rect 3510 7692 3516 7744
rect 3568 7732 3574 7744
rect 8772 7732 8800 7772
rect 13906 7760 13912 7772
rect 13964 7760 13970 7812
rect 3568 7704 8800 7732
rect 3568 7692 3574 7704
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 1486 7528 1492 7540
rect 1447 7500 1492 7528
rect 1486 7488 1492 7500
rect 1544 7488 1550 7540
rect 3878 7528 3884 7540
rect 3839 7500 3884 7528
rect 3878 7488 3884 7500
rect 3936 7488 3942 7540
rect 5626 7488 5632 7540
rect 5684 7528 5690 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 5684 7500 6377 7528
rect 5684 7488 5690 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 8110 7488 8116 7540
rect 8168 7528 8174 7540
rect 8297 7531 8355 7537
rect 8297 7528 8309 7531
rect 8168 7500 8309 7528
rect 8168 7488 8174 7500
rect 8297 7497 8309 7500
rect 8343 7497 8355 7531
rect 8297 7491 8355 7497
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 3970 7392 3976 7404
rect 2179 7364 2636 7392
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 2498 7324 2504 7336
rect 2459 7296 2504 7324
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 2608 7324 2636 7364
rect 3804 7364 3976 7392
rect 2768 7327 2826 7333
rect 2768 7324 2780 7327
rect 2608 7296 2780 7324
rect 2768 7293 2780 7296
rect 2814 7324 2826 7327
rect 3602 7324 3608 7336
rect 2814 7296 3608 7324
rect 2814 7293 2826 7296
rect 2768 7287 2826 7293
rect 3602 7284 3608 7296
rect 3660 7324 3666 7336
rect 3804 7324 3832 7364
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 6914 7392 6920 7404
rect 6875 7364 6920 7392
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 8312 7392 8340 7491
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 8573 7531 8631 7537
rect 8573 7528 8585 7531
rect 8536 7500 8585 7528
rect 8536 7488 8542 7500
rect 8573 7497 8585 7500
rect 8619 7497 8631 7531
rect 8573 7491 8631 7497
rect 16393 7531 16451 7537
rect 16393 7497 16405 7531
rect 16439 7528 16451 7531
rect 17402 7528 17408 7540
rect 16439 7500 17408 7528
rect 16439 7497 16451 7500
rect 16393 7491 16451 7497
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18049 7531 18107 7537
rect 18049 7528 18061 7531
rect 18012 7500 18061 7528
rect 18012 7488 18018 7500
rect 18049 7497 18061 7500
rect 18095 7497 18107 7531
rect 19886 7528 19892 7540
rect 18049 7491 18107 7497
rect 18340 7500 19196 7528
rect 19847 7500 19892 7528
rect 14274 7420 14280 7472
rect 14332 7460 14338 7472
rect 18340 7460 18368 7500
rect 14332 7432 18368 7460
rect 14332 7420 14338 7432
rect 18414 7420 18420 7472
rect 18472 7460 18478 7472
rect 18874 7460 18880 7472
rect 18472 7432 18880 7460
rect 18472 7420 18478 7432
rect 18874 7420 18880 7432
rect 18932 7460 18938 7472
rect 19058 7460 19064 7472
rect 18932 7432 19064 7460
rect 18932 7420 18938 7432
rect 19058 7420 19064 7432
rect 19116 7420 19122 7472
rect 9125 7395 9183 7401
rect 9125 7392 9137 7395
rect 8312 7364 9137 7392
rect 9125 7361 9137 7364
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17126 7392 17132 7404
rect 17083 7364 17132 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17126 7352 17132 7364
rect 17184 7392 17190 7404
rect 18046 7392 18052 7404
rect 17184 7364 18052 7392
rect 17184 7352 17190 7364
rect 18046 7352 18052 7364
rect 18104 7392 18110 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 18104 7364 18613 7392
rect 18104 7352 18110 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 19168 7392 19196 7500
rect 19886 7488 19892 7500
rect 19944 7488 19950 7540
rect 19337 7395 19395 7401
rect 19337 7392 19349 7395
rect 19168 7364 19349 7392
rect 18601 7355 18659 7361
rect 19337 7361 19349 7364
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 20346 7352 20352 7404
rect 20404 7392 20410 7404
rect 20441 7395 20499 7401
rect 20441 7392 20453 7395
rect 20404 7364 20453 7392
rect 20404 7352 20410 7364
rect 20441 7361 20453 7364
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 3660 7296 3832 7324
rect 3660 7284 3666 7296
rect 3878 7284 3884 7336
rect 3936 7324 3942 7336
rect 4985 7327 5043 7333
rect 4985 7324 4997 7327
rect 3936 7296 4997 7324
rect 3936 7284 3942 7296
rect 4985 7293 4997 7296
rect 5031 7293 5043 7327
rect 4985 7287 5043 7293
rect 5074 7284 5080 7336
rect 5132 7324 5138 7336
rect 5252 7327 5310 7333
rect 5252 7324 5264 7327
rect 5132 7296 5264 7324
rect 5132 7284 5138 7296
rect 5252 7293 5264 7296
rect 5298 7324 5310 7327
rect 6822 7324 6828 7336
rect 5298 7296 6828 7324
rect 5298 7293 5310 7296
rect 5252 7287 5310 7293
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 9030 7284 9036 7336
rect 9088 7324 9094 7336
rect 16853 7327 16911 7333
rect 16853 7324 16865 7327
rect 9088 7296 16865 7324
rect 9088 7284 9094 7296
rect 16853 7293 16865 7296
rect 16899 7293 16911 7327
rect 19153 7327 19211 7333
rect 16853 7287 16911 7293
rect 18248 7296 18543 7324
rect 1949 7259 2007 7265
rect 1949 7225 1961 7259
rect 1995 7256 2007 7259
rect 2682 7256 2688 7268
rect 1995 7228 2688 7256
rect 1995 7225 2007 7228
rect 1949 7219 2007 7225
rect 2682 7216 2688 7228
rect 2740 7256 2746 7268
rect 3786 7256 3792 7268
rect 2740 7228 3792 7256
rect 2740 7216 2746 7228
rect 3786 7216 3792 7228
rect 3844 7216 3850 7268
rect 7098 7216 7104 7268
rect 7156 7265 7162 7268
rect 7156 7259 7220 7265
rect 7156 7225 7174 7259
rect 7208 7225 7220 7259
rect 7156 7219 7220 7225
rect 8941 7259 8999 7265
rect 8941 7225 8953 7259
rect 8987 7256 8999 7259
rect 12066 7256 12072 7268
rect 8987 7228 12072 7256
rect 8987 7225 8999 7228
rect 8941 7219 8999 7225
rect 7156 7216 7162 7219
rect 12066 7216 12072 7228
rect 12124 7256 12130 7268
rect 16761 7259 16819 7265
rect 16761 7256 16773 7259
rect 12124 7228 16773 7256
rect 12124 7216 12130 7228
rect 16761 7225 16773 7228
rect 16807 7225 16819 7259
rect 18248 7256 18276 7296
rect 18414 7256 18420 7268
rect 16761 7219 16819 7225
rect 16868 7228 18276 7256
rect 18375 7228 18420 7256
rect 1854 7188 1860 7200
rect 1767 7160 1860 7188
rect 1854 7148 1860 7160
rect 1912 7188 1918 7200
rect 4154 7188 4160 7200
rect 1912 7160 4160 7188
rect 1912 7148 1918 7160
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 4525 7191 4583 7197
rect 4525 7157 4537 7191
rect 4571 7188 4583 7191
rect 5350 7188 5356 7200
rect 4571 7160 5356 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 8386 7148 8392 7200
rect 8444 7188 8450 7200
rect 9030 7188 9036 7200
rect 8444 7160 9036 7188
rect 8444 7148 8450 7160
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 16868 7188 16896 7228
rect 18414 7216 18420 7228
rect 18472 7216 18478 7268
rect 18515 7256 18543 7296
rect 19153 7293 19165 7327
rect 19199 7324 19211 7327
rect 19794 7324 19800 7336
rect 19199 7296 19800 7324
rect 19199 7293 19211 7296
rect 19153 7287 19211 7293
rect 19794 7284 19800 7296
rect 19852 7284 19858 7336
rect 20257 7259 20315 7265
rect 20257 7256 20269 7259
rect 18515 7228 20269 7256
rect 20257 7225 20269 7228
rect 20303 7225 20315 7259
rect 20257 7219 20315 7225
rect 12032 7160 16896 7188
rect 12032 7148 12038 7160
rect 17678 7148 17684 7200
rect 17736 7188 17742 7200
rect 18509 7191 18567 7197
rect 18509 7188 18521 7191
rect 17736 7160 18521 7188
rect 17736 7148 17742 7160
rect 18509 7157 18521 7160
rect 18555 7188 18567 7191
rect 19058 7188 19064 7200
rect 18555 7160 19064 7188
rect 18555 7157 18567 7160
rect 18509 7151 18567 7157
rect 19058 7148 19064 7160
rect 19116 7148 19122 7200
rect 20349 7191 20407 7197
rect 20349 7157 20361 7191
rect 20395 7188 20407 7191
rect 20438 7188 20444 7200
rect 20395 7160 20444 7188
rect 20395 7157 20407 7160
rect 20349 7151 20407 7157
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 18046 6984 18052 6996
rect 18007 6956 18052 6984
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 1578 6876 1584 6928
rect 1636 6916 1642 6928
rect 2498 6916 2504 6928
rect 1636 6888 2504 6916
rect 1636 6876 1642 6888
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 1688 6780 1716 6888
rect 2498 6876 2504 6888
rect 2556 6916 2562 6928
rect 3878 6916 3884 6928
rect 2556 6888 3884 6916
rect 2556 6876 2562 6888
rect 3878 6876 3884 6888
rect 3936 6876 3942 6928
rect 4525 6919 4583 6925
rect 4525 6885 4537 6919
rect 4571 6916 4583 6919
rect 4798 6916 4804 6928
rect 4571 6888 4804 6916
rect 4571 6885 4583 6888
rect 4525 6879 4583 6885
rect 4798 6876 4804 6888
rect 4856 6916 4862 6928
rect 5258 6916 5264 6928
rect 4856 6888 5264 6916
rect 4856 6876 4862 6888
rect 5258 6876 5264 6888
rect 5316 6876 5322 6928
rect 6638 6876 6644 6928
rect 6696 6876 6702 6928
rect 1848 6851 1906 6857
rect 1848 6817 1860 6851
rect 1894 6848 1906 6851
rect 2222 6848 2228 6860
rect 1894 6820 2228 6848
rect 1894 6817 1906 6820
rect 1848 6811 1906 6817
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 5534 6848 5540 6860
rect 5495 6820 5540 6848
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 6546 6848 6552 6860
rect 6507 6820 6552 6848
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 6656 6848 6684 6876
rect 7558 6848 7564 6860
rect 6656 6820 7564 6848
rect 7558 6808 7564 6820
rect 7616 6808 7622 6860
rect 7653 6851 7711 6857
rect 7653 6817 7665 6851
rect 7699 6848 7711 6851
rect 11146 6848 11152 6860
rect 7699 6820 11152 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 16666 6848 16672 6860
rect 16627 6820 16672 6848
rect 16666 6808 16672 6820
rect 16724 6808 16730 6860
rect 16936 6851 16994 6857
rect 16936 6817 16948 6851
rect 16982 6848 16994 6851
rect 19242 6848 19248 6860
rect 16982 6820 19248 6848
rect 16982 6817 16994 6820
rect 16936 6811 16994 6817
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 19420 6851 19478 6857
rect 19420 6817 19432 6851
rect 19466 6848 19478 6851
rect 19702 6848 19708 6860
rect 19466 6820 19708 6848
rect 19466 6817 19478 6820
rect 19420 6811 19478 6817
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 3326 6780 3332 6792
rect 1627 6752 1716 6780
rect 3287 6752 3332 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 4304 6752 4629 6780
rect 4304 6740 4310 6752
rect 4617 6749 4629 6752
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6780 4859 6783
rect 5074 6780 5080 6792
rect 4847 6752 5080 6780
rect 4847 6749 4859 6752
rect 4801 6743 4859 6749
rect 5074 6740 5080 6752
rect 5132 6740 5138 6792
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 2961 6715 3019 6721
rect 2961 6681 2973 6715
rect 3007 6712 3019 6715
rect 3234 6712 3240 6724
rect 3007 6684 3240 6712
rect 3007 6681 3019 6684
rect 2961 6675 3019 6681
rect 3234 6672 3240 6684
rect 3292 6672 3298 6724
rect 4157 6715 4215 6721
rect 4157 6681 4169 6715
rect 4203 6712 4215 6715
rect 5644 6712 5672 6743
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 6641 6783 6699 6789
rect 5776 6752 5821 6780
rect 5776 6740 5782 6752
rect 6641 6749 6653 6783
rect 6687 6749 6699 6783
rect 6822 6780 6828 6792
rect 6783 6752 6828 6780
rect 6641 6743 6699 6749
rect 4203 6684 5672 6712
rect 6656 6712 6684 6743
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6780 7895 6783
rect 9674 6780 9680 6792
rect 7883 6752 9680 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 19150 6780 19156 6792
rect 19111 6752 19156 6780
rect 19150 6740 19156 6752
rect 19208 6740 19214 6792
rect 20162 6740 20168 6792
rect 20220 6780 20226 6792
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20220 6752 20913 6780
rect 20220 6740 20226 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 7193 6715 7251 6721
rect 7193 6712 7205 6715
rect 6656 6684 7205 6712
rect 4203 6681 4215 6684
rect 4157 6675 4215 6681
rect 7193 6681 7205 6684
rect 7239 6681 7251 6715
rect 7193 6675 7251 6681
rect 5166 6644 5172 6656
rect 5127 6616 5172 6644
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 5626 6604 5632 6656
rect 5684 6644 5690 6656
rect 6181 6647 6239 6653
rect 6181 6644 6193 6647
rect 5684 6616 6193 6644
rect 5684 6604 5690 6616
rect 6181 6613 6193 6616
rect 6227 6613 6239 6647
rect 6181 6607 6239 6613
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 17954 6644 17960 6656
rect 7524 6616 17960 6644
rect 7524 6604 7530 6616
rect 17954 6604 17960 6616
rect 18012 6604 18018 6656
rect 20533 6647 20591 6653
rect 20533 6613 20545 6647
rect 20579 6644 20591 6647
rect 20622 6644 20628 6656
rect 20579 6616 20628 6644
rect 20579 6613 20591 6616
rect 20533 6607 20591 6613
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 2958 6440 2964 6452
rect 2919 6412 2964 6440
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 4985 6443 5043 6449
rect 4985 6409 4997 6443
rect 5031 6440 5043 6443
rect 5534 6440 5540 6452
rect 5031 6412 5540 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 20346 6440 20352 6452
rect 19300 6412 20352 6440
rect 19300 6400 19306 6412
rect 20346 6400 20352 6412
rect 20404 6440 20410 6452
rect 20717 6443 20775 6449
rect 20717 6440 20729 6443
rect 20404 6412 20729 6440
rect 20404 6400 20410 6412
rect 20717 6409 20729 6412
rect 20763 6409 20775 6443
rect 20717 6403 20775 6409
rect 3602 6304 3608 6316
rect 3563 6276 3608 6304
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 5074 6264 5080 6316
rect 5132 6304 5138 6316
rect 5537 6307 5595 6313
rect 5537 6304 5549 6307
rect 5132 6276 5549 6304
rect 5132 6264 5138 6276
rect 5537 6273 5549 6276
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 19150 6264 19156 6316
rect 19208 6304 19214 6316
rect 19337 6307 19395 6313
rect 19337 6304 19349 6307
rect 19208 6276 19349 6304
rect 19208 6264 19214 6276
rect 19337 6273 19349 6276
rect 19383 6273 19395 6307
rect 19337 6267 19395 6273
rect 3326 6236 3332 6248
rect 3287 6208 3332 6236
rect 3326 6196 3332 6208
rect 3384 6196 3390 6248
rect 5350 6236 5356 6248
rect 5311 6208 5356 6236
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 10042 6168 10048 6180
rect 4120 6140 10048 6168
rect 4120 6128 4126 6140
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 19604 6171 19662 6177
rect 19604 6137 19616 6171
rect 19650 6168 19662 6171
rect 20622 6168 20628 6180
rect 19650 6140 20628 6168
rect 19650 6137 19662 6140
rect 19604 6131 19662 6137
rect 20622 6128 20628 6140
rect 20680 6128 20686 6180
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 3421 6103 3479 6109
rect 3421 6100 3433 6103
rect 3384 6072 3433 6100
rect 3384 6060 3390 6072
rect 3421 6069 3433 6072
rect 3467 6100 3479 6103
rect 3694 6100 3700 6112
rect 3467 6072 3700 6100
rect 3467 6069 3479 6072
rect 3421 6063 3479 6069
rect 3694 6060 3700 6072
rect 3752 6060 3758 6112
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 4890 6100 4896 6112
rect 4212 6072 4896 6100
rect 4212 6060 4218 6072
rect 4890 6060 4896 6072
rect 4948 6100 4954 6112
rect 5445 6103 5503 6109
rect 5445 6100 5457 6103
rect 4948 6072 5457 6100
rect 4948 6060 4954 6072
rect 5445 6069 5457 6072
rect 5491 6069 5503 6103
rect 5445 6063 5503 6069
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 8294 5896 8300 5908
rect 4028 5868 8300 5896
rect 4028 5856 4034 5868
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 19794 5896 19800 5908
rect 19755 5868 19800 5896
rect 19794 5856 19800 5868
rect 19852 5856 19858 5908
rect 20162 5896 20168 5908
rect 20123 5868 20168 5896
rect 20162 5856 20168 5868
rect 20220 5856 20226 5908
rect 20254 5692 20260 5704
rect 20215 5664 20260 5692
rect 20254 5652 20260 5664
rect 20312 5652 20318 5704
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20404 5664 20449 5692
rect 20404 5652 20410 5664
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 5902 5312 5908 5364
rect 5960 5352 5966 5364
rect 17954 5352 17960 5364
rect 5960 5324 17960 5352
rect 5960 5312 5966 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 20073 5355 20131 5361
rect 20073 5321 20085 5355
rect 20119 5352 20131 5355
rect 20254 5352 20260 5364
rect 20119 5324 20260 5352
rect 20119 5321 20131 5324
rect 20073 5315 20131 5321
rect 20254 5312 20260 5324
rect 20312 5312 20318 5364
rect 4062 5244 4068 5296
rect 4120 5284 4126 5296
rect 11974 5284 11980 5296
rect 4120 5256 11980 5284
rect 4120 5244 4126 5256
rect 11974 5244 11980 5256
rect 12032 5244 12038 5296
rect 20622 5216 20628 5228
rect 20583 5188 20628 5216
rect 20622 5176 20628 5188
rect 20680 5176 20686 5228
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 19889 5015 19947 5021
rect 19889 5012 19901 5015
rect 4120 4984 19901 5012
rect 4120 4972 4126 4984
rect 19889 4981 19901 4984
rect 19935 5012 19947 5015
rect 20441 5015 20499 5021
rect 20441 5012 20453 5015
rect 19935 4984 20453 5012
rect 19935 4981 19947 4984
rect 19889 4975 19947 4981
rect 20441 4981 20453 4984
rect 20487 4981 20499 5015
rect 20441 4975 20499 4981
rect 20530 4972 20536 5024
rect 20588 5012 20594 5024
rect 20588 4984 20633 5012
rect 20588 4972 20594 4984
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 6362 3068 6368 3120
rect 6420 3108 6426 3120
rect 6420 3080 15516 3108
rect 6420 3068 6426 3080
rect 4982 3040 4988 3052
rect 4943 3012 4988 3040
rect 4982 3000 4988 3012
rect 5040 3000 5046 3052
rect 5810 3040 5816 3052
rect 5771 3012 5816 3040
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 15488 3049 15516 3080
rect 15473 3043 15531 3049
rect 15473 3009 15485 3043
rect 15519 3009 15531 3043
rect 15473 3003 15531 3009
rect 4709 2975 4767 2981
rect 4709 2941 4721 2975
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 5629 2975 5687 2981
rect 5629 2941 5641 2975
rect 5675 2972 5687 2975
rect 11146 2972 11152 2984
rect 5675 2944 11152 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 4724 2904 4752 2935
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 15197 2975 15255 2981
rect 15197 2941 15209 2975
rect 15243 2972 15255 2975
rect 15838 2972 15844 2984
rect 15243 2944 15844 2972
rect 15243 2941 15255 2944
rect 15197 2935 15255 2941
rect 15838 2932 15844 2944
rect 15896 2932 15902 2984
rect 20438 2904 20444 2916
rect 4724 2876 20444 2904
rect 20438 2864 20444 2876
rect 20496 2864 20502 2916
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 2774 960 2780 1012
rect 2832 1000 2838 1012
rect 4706 1000 4712 1012
rect 2832 972 4712 1000
rect 2832 960 2838 972
rect 4706 960 4712 972
rect 4764 960 4770 1012
<< via1 >>
rect 3700 20952 3752 21004
rect 6092 20952 6144 21004
rect 14372 20272 14424 20324
rect 14924 20272 14976 20324
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 2780 20000 2832 20052
rect 11152 20000 11204 20052
rect 11612 20000 11664 20052
rect 12164 20000 12216 20052
rect 12716 20000 12768 20052
rect 13268 20000 13320 20052
rect 204 19932 256 19984
rect 2504 19932 2556 19984
rect 3240 19932 3292 19984
rect 12440 19932 12492 19984
rect 17040 20000 17092 20052
rect 17500 20000 17552 20052
rect 18328 20000 18380 20052
rect 18788 20000 18840 20052
rect 19616 20043 19668 20052
rect 19616 20009 19625 20043
rect 19625 20009 19659 20043
rect 19659 20009 19668 20043
rect 19616 20000 19668 20009
rect 20168 20043 20220 20052
rect 20168 20009 20177 20043
rect 20177 20009 20211 20043
rect 20211 20009 20220 20043
rect 20168 20000 20220 20009
rect 20628 20000 20680 20052
rect 17868 19932 17920 19984
rect 3332 19864 3384 19916
rect 8484 19864 8536 19916
rect 9588 19864 9640 19916
rect 3148 19796 3200 19848
rect 3700 19796 3752 19848
rect 8852 19839 8904 19848
rect 8852 19805 8861 19839
rect 8861 19805 8895 19839
rect 8895 19805 8904 19839
rect 8852 19796 8904 19805
rect 4160 19728 4212 19780
rect 7564 19728 7616 19780
rect 10416 19864 10468 19916
rect 11152 19864 11204 19916
rect 11612 19864 11664 19916
rect 13268 19907 13320 19916
rect 13268 19873 13277 19907
rect 13277 19873 13311 19907
rect 13311 19873 13320 19907
rect 13268 19864 13320 19873
rect 14188 19907 14240 19916
rect 14188 19873 14197 19907
rect 14197 19873 14231 19907
rect 14231 19873 14240 19907
rect 14188 19864 14240 19873
rect 14740 19907 14792 19916
rect 14740 19873 14749 19907
rect 14749 19873 14783 19907
rect 14783 19873 14792 19907
rect 14740 19864 14792 19873
rect 15016 19864 15068 19916
rect 16028 19864 16080 19916
rect 16764 19864 16816 19916
rect 9956 19796 10008 19848
rect 10508 19839 10560 19848
rect 10508 19805 10517 19839
rect 10517 19805 10551 19839
rect 10551 19805 10560 19839
rect 10508 19796 10560 19805
rect 11796 19796 11848 19848
rect 13360 19839 13412 19848
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 16580 19796 16632 19848
rect 18512 19864 18564 19916
rect 19432 19907 19484 19916
rect 17960 19796 18012 19848
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 19340 19796 19392 19848
rect 19616 19796 19668 19848
rect 16672 19728 16724 19780
rect 19064 19771 19116 19780
rect 19064 19737 19073 19771
rect 19073 19737 19107 19771
rect 19107 19737 19116 19771
rect 19064 19728 19116 19737
rect 2596 19703 2648 19712
rect 2596 19669 2605 19703
rect 2605 19669 2639 19703
rect 2639 19669 2648 19703
rect 2596 19660 2648 19669
rect 3148 19703 3200 19712
rect 3148 19669 3157 19703
rect 3157 19669 3191 19703
rect 3191 19669 3200 19703
rect 3148 19660 3200 19669
rect 8300 19703 8352 19712
rect 8300 19669 8309 19703
rect 8309 19669 8343 19703
rect 8343 19669 8352 19703
rect 8300 19660 8352 19669
rect 9496 19660 9548 19712
rect 11060 19660 11112 19712
rect 14096 19660 14148 19712
rect 18604 19660 18656 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 3424 19499 3476 19508
rect 3424 19465 3433 19499
rect 3433 19465 3467 19499
rect 3467 19465 3476 19499
rect 3424 19456 3476 19465
rect 6092 19499 6144 19508
rect 6092 19465 6101 19499
rect 6101 19465 6135 19499
rect 6135 19465 6144 19499
rect 6092 19456 6144 19465
rect 8852 19456 8904 19508
rect 9956 19456 10008 19508
rect 2136 19252 2188 19304
rect 2320 19295 2372 19304
rect 2320 19261 2329 19295
rect 2329 19261 2363 19295
rect 2363 19261 2372 19295
rect 2320 19252 2372 19261
rect 3976 19295 4028 19304
rect 3976 19261 3985 19295
rect 3985 19261 4019 19295
rect 4019 19261 4028 19295
rect 3976 19252 4028 19261
rect 5540 19252 5592 19304
rect 5908 19295 5960 19304
rect 5908 19261 5917 19295
rect 5917 19261 5951 19295
rect 5951 19261 5960 19295
rect 5908 19252 5960 19261
rect 1032 19184 1084 19236
rect 6644 19184 6696 19236
rect 2872 19116 2924 19168
rect 4160 19116 4212 19168
rect 4252 19116 4304 19168
rect 4988 19116 5040 19168
rect 7288 19252 7340 19304
rect 9404 19388 9456 19440
rect 8300 19320 8352 19372
rect 14740 19320 14792 19372
rect 15476 19363 15528 19372
rect 15476 19329 15485 19363
rect 15485 19329 15519 19363
rect 15519 19329 15528 19363
rect 15476 19320 15528 19329
rect 8668 19252 8720 19304
rect 10048 19252 10100 19304
rect 13176 19252 13228 19304
rect 14096 19295 14148 19304
rect 14096 19261 14105 19295
rect 14105 19261 14139 19295
rect 14139 19261 14148 19295
rect 14096 19252 14148 19261
rect 7656 19116 7708 19168
rect 8944 19116 8996 19168
rect 9220 19159 9272 19168
rect 9220 19125 9229 19159
rect 9229 19125 9263 19159
rect 9263 19125 9272 19159
rect 9220 19116 9272 19125
rect 9312 19116 9364 19168
rect 11704 19184 11756 19236
rect 12808 19184 12860 19236
rect 11796 19159 11848 19168
rect 11796 19125 11805 19159
rect 11805 19125 11839 19159
rect 11839 19125 11848 19159
rect 11796 19116 11848 19125
rect 12440 19116 12492 19168
rect 14556 19184 14608 19236
rect 13544 19116 13596 19168
rect 16580 19252 16632 19304
rect 18236 19320 18288 19372
rect 18512 19320 18564 19372
rect 18604 19320 18656 19372
rect 19248 19295 19300 19304
rect 19248 19261 19257 19295
rect 19257 19261 19291 19295
rect 19291 19261 19300 19295
rect 19248 19252 19300 19261
rect 15568 19184 15620 19236
rect 19340 19184 19392 19236
rect 19524 19227 19576 19236
rect 19524 19193 19533 19227
rect 19533 19193 19567 19227
rect 19567 19193 19576 19227
rect 19524 19184 19576 19193
rect 20076 19252 20128 19304
rect 20536 19295 20588 19304
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 22100 19184 22152 19236
rect 15200 19159 15252 19168
rect 15200 19125 15209 19159
rect 15209 19125 15243 19159
rect 15243 19125 15252 19159
rect 15200 19116 15252 19125
rect 15936 19116 15988 19168
rect 17316 19159 17368 19168
rect 17316 19125 17325 19159
rect 17325 19125 17359 19159
rect 17359 19125 17368 19159
rect 17316 19116 17368 19125
rect 17408 19159 17460 19168
rect 17408 19125 17417 19159
rect 17417 19125 17451 19159
rect 17451 19125 17460 19159
rect 17408 19116 17460 19125
rect 17592 19116 17644 19168
rect 19156 19116 19208 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 2780 18912 2832 18964
rect 3792 18912 3844 18964
rect 4252 18955 4304 18964
rect 4252 18921 4261 18955
rect 4261 18921 4295 18955
rect 4295 18921 4304 18955
rect 4252 18912 4304 18921
rect 5908 18844 5960 18896
rect 8760 18912 8812 18964
rect 9404 18912 9456 18964
rect 13360 18912 13412 18964
rect 15292 18912 15344 18964
rect 2504 18819 2556 18828
rect 2504 18785 2513 18819
rect 2513 18785 2547 18819
rect 2547 18785 2556 18819
rect 2504 18776 2556 18785
rect 3608 18776 3660 18828
rect 4896 18776 4948 18828
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 8852 18776 8904 18828
rect 9404 18776 9456 18828
rect 3884 18708 3936 18760
rect 3976 18708 4028 18760
rect 7564 18708 7616 18760
rect 9680 18751 9732 18760
rect 2964 18640 3016 18692
rect 3240 18683 3292 18692
rect 3240 18649 3249 18683
rect 3249 18649 3283 18683
rect 3283 18649 3292 18683
rect 3240 18640 3292 18649
rect 3700 18640 3752 18692
rect 5080 18640 5132 18692
rect 7656 18640 7708 18692
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 13084 18844 13136 18896
rect 13544 18844 13596 18896
rect 15476 18844 15528 18896
rect 11060 18776 11112 18828
rect 16028 18776 16080 18828
rect 18236 18912 18288 18964
rect 17500 18844 17552 18896
rect 12624 18751 12676 18760
rect 12624 18717 12633 18751
rect 12633 18717 12667 18751
rect 12667 18717 12676 18751
rect 12624 18708 12676 18717
rect 12808 18751 12860 18760
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 13176 18751 13228 18760
rect 13176 18717 13185 18751
rect 13185 18717 13219 18751
rect 13219 18717 13228 18751
rect 13176 18708 13228 18717
rect 15292 18708 15344 18760
rect 10784 18572 10836 18624
rect 14280 18640 14332 18692
rect 12440 18572 12492 18624
rect 12532 18572 12584 18624
rect 13912 18572 13964 18624
rect 14556 18615 14608 18624
rect 14556 18581 14565 18615
rect 14565 18581 14599 18615
rect 14599 18581 14608 18615
rect 14556 18572 14608 18581
rect 19432 18572 19484 18624
rect 20168 18615 20220 18624
rect 20168 18581 20177 18615
rect 20177 18581 20211 18615
rect 20211 18581 20220 18615
rect 20168 18572 20220 18581
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 3056 18368 3108 18420
rect 3976 18368 4028 18420
rect 4160 18368 4212 18420
rect 3516 18300 3568 18352
rect 6736 18300 6788 18352
rect 2504 18232 2556 18284
rect 3792 18232 3844 18284
rect 4896 18275 4948 18284
rect 3516 18164 3568 18216
rect 4160 18164 4212 18216
rect 4896 18241 4905 18275
rect 4905 18241 4939 18275
rect 4939 18241 4948 18275
rect 4896 18232 4948 18241
rect 5632 18232 5684 18284
rect 6368 18232 6420 18284
rect 6460 18232 6512 18284
rect 7288 18232 7340 18284
rect 4804 18164 4856 18216
rect 6828 18164 6880 18216
rect 6092 18096 6144 18148
rect 6184 18096 6236 18148
rect 6920 18096 6972 18148
rect 9220 18368 9272 18420
rect 7472 18232 7524 18284
rect 7748 18232 7800 18284
rect 8852 18275 8904 18284
rect 8852 18241 8861 18275
rect 8861 18241 8895 18275
rect 8895 18241 8904 18275
rect 13268 18368 13320 18420
rect 15476 18368 15528 18420
rect 15936 18411 15988 18420
rect 15936 18377 15945 18411
rect 15945 18377 15979 18411
rect 15979 18377 15988 18411
rect 15936 18368 15988 18377
rect 17316 18368 17368 18420
rect 18880 18368 18932 18420
rect 20812 18411 20864 18420
rect 20812 18377 20821 18411
rect 20821 18377 20855 18411
rect 20855 18377 20864 18411
rect 20812 18368 20864 18377
rect 11704 18300 11756 18352
rect 12256 18300 12308 18352
rect 13176 18300 13228 18352
rect 8852 18232 8904 18241
rect 8576 18207 8628 18216
rect 8576 18173 8585 18207
rect 8585 18173 8619 18207
rect 8619 18173 8628 18207
rect 8576 18164 8628 18173
rect 8944 18164 8996 18216
rect 7012 18071 7064 18080
rect 7012 18037 7021 18071
rect 7021 18037 7055 18071
rect 7055 18037 7064 18071
rect 7012 18028 7064 18037
rect 8668 18139 8720 18148
rect 8668 18105 8677 18139
rect 8677 18105 8711 18139
rect 8711 18105 8720 18139
rect 8668 18096 8720 18105
rect 11244 18232 11296 18284
rect 11980 18232 12032 18284
rect 12808 18232 12860 18284
rect 16764 18300 16816 18352
rect 19340 18300 19392 18352
rect 17500 18275 17552 18284
rect 9680 18164 9732 18216
rect 10232 18164 10284 18216
rect 10784 18164 10836 18216
rect 12532 18164 12584 18216
rect 13544 18164 13596 18216
rect 9772 18096 9824 18148
rect 10600 18096 10652 18148
rect 12072 18096 12124 18148
rect 13452 18096 13504 18148
rect 14556 18139 14608 18148
rect 14556 18105 14590 18139
rect 14590 18105 14608 18139
rect 14556 18096 14608 18105
rect 15844 18096 15896 18148
rect 17500 18241 17509 18275
rect 17509 18241 17543 18275
rect 17543 18241 17552 18275
rect 17500 18232 17552 18241
rect 19156 18232 19208 18284
rect 20168 18275 20220 18284
rect 20168 18241 20177 18275
rect 20177 18241 20211 18275
rect 20211 18241 20220 18275
rect 20168 18232 20220 18241
rect 17592 18164 17644 18216
rect 19524 18164 19576 18216
rect 20260 18164 20312 18216
rect 9220 18028 9272 18080
rect 10876 18028 10928 18080
rect 11796 18071 11848 18080
rect 11796 18037 11805 18071
rect 11805 18037 11839 18071
rect 11839 18037 11848 18071
rect 11796 18028 11848 18037
rect 16304 18071 16356 18080
rect 16304 18037 16313 18071
rect 16313 18037 16347 18071
rect 16347 18037 16356 18071
rect 16304 18028 16356 18037
rect 16488 18028 16540 18080
rect 17592 18028 17644 18080
rect 18880 18028 18932 18080
rect 19432 18028 19484 18080
rect 19984 18071 20036 18080
rect 19984 18037 19993 18071
rect 19993 18037 20027 18071
rect 20027 18037 20036 18071
rect 19984 18028 20036 18037
rect 20168 18028 20220 18080
rect 20536 18028 20588 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 2504 17867 2556 17876
rect 2504 17833 2513 17867
rect 2513 17833 2547 17867
rect 2547 17833 2556 17867
rect 2504 17824 2556 17833
rect 3792 17824 3844 17876
rect 7564 17824 7616 17876
rect 7656 17824 7708 17876
rect 8300 17824 8352 17876
rect 9496 17824 9548 17876
rect 9772 17824 9824 17876
rect 11152 17824 11204 17876
rect 11796 17824 11848 17876
rect 12808 17824 12860 17876
rect 6000 17756 6052 17808
rect 6828 17756 6880 17808
rect 9220 17756 9272 17808
rect 9312 17756 9364 17808
rect 12532 17756 12584 17808
rect 12624 17756 12676 17808
rect 15200 17824 15252 17876
rect 16212 17824 16264 17876
rect 17408 17824 17460 17876
rect 18604 17867 18656 17876
rect 18604 17833 18613 17867
rect 18613 17833 18647 17867
rect 18647 17833 18656 17867
rect 18604 17824 18656 17833
rect 2320 17731 2372 17740
rect 2320 17697 2329 17731
rect 2329 17697 2363 17731
rect 2363 17697 2372 17731
rect 2320 17688 2372 17697
rect 2964 17688 3016 17740
rect 4252 17688 4304 17740
rect 5908 17731 5960 17740
rect 5908 17697 5942 17731
rect 5942 17697 5960 17731
rect 5908 17688 5960 17697
rect 7472 17688 7524 17740
rect 7656 17731 7708 17740
rect 7656 17697 7665 17731
rect 7665 17697 7699 17731
rect 7699 17697 7708 17731
rect 7656 17688 7708 17697
rect 8576 17688 8628 17740
rect 8944 17731 8996 17740
rect 8944 17697 8953 17731
rect 8953 17697 8987 17731
rect 8987 17697 8996 17731
rect 8944 17688 8996 17697
rect 2596 17620 2648 17672
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 4804 17620 4856 17672
rect 6828 17620 6880 17672
rect 9772 17688 9824 17740
rect 10508 17688 10560 17740
rect 10968 17688 11020 17740
rect 11704 17688 11756 17740
rect 13268 17688 13320 17740
rect 9680 17663 9732 17672
rect 7472 17552 7524 17604
rect 9680 17629 9689 17663
rect 9689 17629 9723 17663
rect 9723 17629 9732 17663
rect 9680 17620 9732 17629
rect 11796 17663 11848 17672
rect 11796 17629 11805 17663
rect 11805 17629 11839 17663
rect 11839 17629 11848 17663
rect 11796 17620 11848 17629
rect 11888 17663 11940 17672
rect 11888 17629 11897 17663
rect 11897 17629 11931 17663
rect 11931 17629 11940 17663
rect 11888 17620 11940 17629
rect 12072 17620 12124 17672
rect 12624 17620 12676 17672
rect 14372 17688 14424 17740
rect 13728 17620 13780 17672
rect 5632 17484 5684 17536
rect 8852 17552 8904 17604
rect 19616 17824 19668 17876
rect 19156 17756 19208 17808
rect 19892 17756 19944 17808
rect 15016 17688 15068 17740
rect 17132 17688 17184 17740
rect 17684 17688 17736 17740
rect 17868 17731 17920 17740
rect 17868 17697 17877 17731
rect 17877 17697 17911 17731
rect 17911 17697 17920 17731
rect 17868 17688 17920 17697
rect 18696 17688 18748 17740
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 17316 17620 17368 17672
rect 17500 17663 17552 17672
rect 17500 17629 17509 17663
rect 17509 17629 17543 17663
rect 17543 17629 17552 17663
rect 17500 17620 17552 17629
rect 8300 17527 8352 17536
rect 8300 17493 8309 17527
rect 8309 17493 8343 17527
rect 8343 17493 8352 17527
rect 8300 17484 8352 17493
rect 14556 17552 14608 17604
rect 18880 17620 18932 17672
rect 11796 17484 11848 17536
rect 12072 17484 12124 17536
rect 13176 17484 13228 17536
rect 13360 17484 13412 17536
rect 17960 17484 18012 17536
rect 19708 17484 19760 17536
rect 19892 17484 19944 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 1952 17323 2004 17332
rect 1952 17289 1961 17323
rect 1961 17289 1995 17323
rect 1995 17289 2004 17323
rect 1952 17280 2004 17289
rect 2780 17280 2832 17332
rect 4160 17280 4212 17332
rect 4804 17280 4856 17332
rect 5908 17280 5960 17332
rect 6828 17323 6880 17332
rect 6828 17289 6837 17323
rect 6837 17289 6871 17323
rect 6871 17289 6880 17323
rect 6828 17280 6880 17289
rect 9588 17280 9640 17332
rect 11060 17280 11112 17332
rect 11612 17280 11664 17332
rect 2688 17212 2740 17264
rect 3792 17144 3844 17196
rect 5632 17212 5684 17264
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 7012 17144 7064 17196
rect 7564 17144 7616 17196
rect 7748 17144 7800 17196
rect 9496 17212 9548 17264
rect 10324 17187 10376 17196
rect 2136 16940 2188 16992
rect 3700 16940 3752 16992
rect 3976 16983 4028 16992
rect 3976 16949 3985 16983
rect 3985 16949 4019 16983
rect 4019 16949 4028 16983
rect 3976 16940 4028 16949
rect 5448 17008 5500 17060
rect 7104 17008 7156 17060
rect 8208 17119 8260 17128
rect 8208 17085 8217 17119
rect 8217 17085 8251 17119
rect 8251 17085 8260 17119
rect 8852 17119 8904 17128
rect 8208 17076 8260 17085
rect 8852 17085 8861 17119
rect 8861 17085 8895 17119
rect 8895 17085 8904 17119
rect 8852 17076 8904 17085
rect 10324 17153 10333 17187
rect 10333 17153 10367 17187
rect 10367 17153 10376 17187
rect 10324 17144 10376 17153
rect 10876 17144 10928 17196
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 12532 17212 12584 17264
rect 13360 17187 13412 17196
rect 13360 17153 13369 17187
rect 13369 17153 13403 17187
rect 13403 17153 13412 17187
rect 13360 17144 13412 17153
rect 13820 17144 13872 17196
rect 14004 17144 14056 17196
rect 14372 17187 14424 17196
rect 14372 17153 14381 17187
rect 14381 17153 14415 17187
rect 14415 17153 14424 17187
rect 14372 17144 14424 17153
rect 15384 17280 15436 17332
rect 16580 17280 16632 17332
rect 17592 17280 17644 17332
rect 15752 17212 15804 17264
rect 15016 17144 15068 17196
rect 17132 17187 17184 17196
rect 8668 17008 8720 17060
rect 8760 17008 8812 17060
rect 9220 17008 9272 17060
rect 8944 16940 8996 16992
rect 9496 16940 9548 16992
rect 9772 16940 9824 16992
rect 9956 17008 10008 17060
rect 14648 17076 14700 17128
rect 17132 17153 17141 17187
rect 17141 17153 17175 17187
rect 17175 17153 17184 17187
rect 17132 17144 17184 17153
rect 17776 17144 17828 17196
rect 16856 17076 16908 17128
rect 15108 17008 15160 17060
rect 17868 17008 17920 17060
rect 11520 16940 11572 16992
rect 11888 16940 11940 16992
rect 12072 16940 12124 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 13176 16940 13228 16992
rect 13544 16940 13596 16992
rect 16488 16940 16540 16992
rect 18788 17008 18840 17060
rect 19248 17280 19300 17332
rect 19892 17280 19944 17332
rect 20168 17280 20220 17332
rect 19156 17212 19208 17264
rect 19340 17144 19392 17196
rect 19800 17144 19852 17196
rect 19984 17144 20036 17196
rect 19524 17119 19576 17128
rect 19524 17085 19533 17119
rect 19533 17085 19567 17119
rect 19567 17085 19576 17119
rect 19524 17076 19576 17085
rect 19616 17076 19668 17128
rect 20536 17119 20588 17128
rect 20536 17085 20545 17119
rect 20545 17085 20579 17119
rect 20579 17085 20588 17119
rect 20536 17076 20588 17085
rect 19156 16940 19208 16992
rect 19432 16983 19484 16992
rect 19432 16949 19441 16983
rect 19441 16949 19475 16983
rect 19475 16949 19484 16983
rect 19432 16940 19484 16949
rect 19616 16940 19668 16992
rect 20260 16940 20312 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1952 16779 2004 16788
rect 1952 16745 1961 16779
rect 1961 16745 1995 16779
rect 1995 16745 2004 16779
rect 1952 16736 2004 16745
rect 2596 16779 2648 16788
rect 2596 16745 2605 16779
rect 2605 16745 2639 16779
rect 2639 16745 2648 16779
rect 2596 16736 2648 16745
rect 3148 16736 3200 16788
rect 5448 16779 5500 16788
rect 5448 16745 5457 16779
rect 5457 16745 5491 16779
rect 5491 16745 5500 16779
rect 5448 16736 5500 16745
rect 10324 16736 10376 16788
rect 10876 16736 10928 16788
rect 14372 16736 14424 16788
rect 15016 16736 15068 16788
rect 18052 16736 18104 16788
rect 19524 16736 19576 16788
rect 4160 16668 4212 16720
rect 4712 16668 4764 16720
rect 3792 16600 3844 16652
rect 4804 16600 4856 16652
rect 7380 16668 7432 16720
rect 7472 16668 7524 16720
rect 7564 16600 7616 16652
rect 3056 16575 3108 16584
rect 3056 16541 3065 16575
rect 3065 16541 3099 16575
rect 3099 16541 3108 16575
rect 3056 16532 3108 16541
rect 3240 16575 3292 16584
rect 3240 16541 3249 16575
rect 3249 16541 3283 16575
rect 3283 16541 3292 16575
rect 3240 16532 3292 16541
rect 7380 16532 7432 16584
rect 8300 16600 8352 16652
rect 9680 16600 9732 16652
rect 9864 16600 9916 16652
rect 10508 16668 10560 16720
rect 10232 16600 10284 16652
rect 12256 16668 12308 16720
rect 12900 16668 12952 16720
rect 16028 16668 16080 16720
rect 17776 16668 17828 16720
rect 5264 16464 5316 16516
rect 5724 16464 5776 16516
rect 7472 16507 7524 16516
rect 7472 16473 7481 16507
rect 7481 16473 7515 16507
rect 7515 16473 7524 16507
rect 7472 16464 7524 16473
rect 5080 16396 5132 16448
rect 10324 16575 10376 16584
rect 9588 16464 9640 16516
rect 10324 16541 10333 16575
rect 10333 16541 10367 16575
rect 10367 16541 10376 16575
rect 10324 16532 10376 16541
rect 11888 16600 11940 16652
rect 9680 16439 9732 16448
rect 9680 16405 9689 16439
rect 9689 16405 9723 16439
rect 9723 16405 9732 16439
rect 9680 16396 9732 16405
rect 14096 16600 14148 16652
rect 15108 16600 15160 16652
rect 15292 16600 15344 16652
rect 13360 16464 13412 16516
rect 15568 16532 15620 16584
rect 15660 16532 15712 16584
rect 12716 16439 12768 16448
rect 12716 16405 12725 16439
rect 12725 16405 12759 16439
rect 12759 16405 12768 16439
rect 13728 16464 13780 16516
rect 15200 16464 15252 16516
rect 15936 16532 15988 16584
rect 15292 16439 15344 16448
rect 12716 16396 12768 16405
rect 15292 16405 15301 16439
rect 15301 16405 15335 16439
rect 15335 16405 15344 16439
rect 15292 16396 15344 16405
rect 19064 16600 19116 16652
rect 19248 16600 19300 16652
rect 19984 16600 20036 16652
rect 20904 16575 20956 16584
rect 20904 16541 20913 16575
rect 20913 16541 20947 16575
rect 20947 16541 20956 16575
rect 20904 16532 20956 16541
rect 18604 16396 18656 16448
rect 18972 16396 19024 16448
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 2228 16056 2280 16108
rect 4160 16192 4212 16244
rect 4252 16192 4304 16244
rect 4804 16192 4856 16244
rect 7656 16192 7708 16244
rect 11796 16192 11848 16244
rect 13820 16192 13872 16244
rect 15568 16235 15620 16244
rect 4252 16056 4304 16108
rect 5264 16056 5316 16108
rect 7656 16056 7708 16108
rect 7748 16056 7800 16108
rect 8208 16056 8260 16108
rect 15568 16201 15577 16235
rect 15577 16201 15611 16235
rect 15611 16201 15620 16235
rect 15568 16192 15620 16201
rect 5080 15988 5132 16040
rect 8576 15988 8628 16040
rect 9680 15988 9732 16040
rect 9864 15988 9916 16040
rect 10876 15988 10928 16040
rect 12532 16031 12584 16040
rect 3240 15920 3292 15972
rect 3700 15920 3752 15972
rect 5448 15920 5500 15972
rect 572 15852 624 15904
rect 2780 15852 2832 15904
rect 4896 15852 4948 15904
rect 7196 15852 7248 15904
rect 7656 15852 7708 15904
rect 9772 15920 9824 15972
rect 12532 15997 12541 16031
rect 12541 15997 12575 16031
rect 12575 15997 12584 16031
rect 12532 15988 12584 15997
rect 14464 16031 14516 16040
rect 14464 15997 14487 16031
rect 14487 15997 14516 16031
rect 15844 16031 15896 16040
rect 14464 15988 14516 15997
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 16856 16056 16908 16108
rect 18604 16056 18656 16108
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 8392 15895 8444 15904
rect 8392 15861 8401 15895
rect 8401 15861 8435 15895
rect 8435 15861 8444 15895
rect 8392 15852 8444 15861
rect 11244 15852 11296 15904
rect 11888 15852 11940 15904
rect 12256 15852 12308 15904
rect 12532 15852 12584 15904
rect 12716 15920 12768 15972
rect 15476 15920 15528 15972
rect 19524 15988 19576 16040
rect 20536 16031 20588 16040
rect 20536 15997 20545 16031
rect 20545 15997 20579 16031
rect 20579 15997 20588 16031
rect 20536 15988 20588 15997
rect 19432 15920 19484 15972
rect 20812 15963 20864 15972
rect 20812 15929 20821 15963
rect 20821 15929 20855 15963
rect 20855 15929 20864 15963
rect 20812 15920 20864 15929
rect 13728 15852 13780 15904
rect 16396 15852 16448 15904
rect 18972 15852 19024 15904
rect 19064 15852 19116 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 2780 15648 2832 15700
rect 3976 15648 4028 15700
rect 5356 15648 5408 15700
rect 3056 15580 3108 15632
rect 3700 15580 3752 15632
rect 5264 15580 5316 15632
rect 2412 15512 2464 15564
rect 3240 15444 3292 15496
rect 4160 15444 4212 15496
rect 4712 15487 4764 15496
rect 4712 15453 4721 15487
rect 4721 15453 4755 15487
rect 4755 15453 4764 15487
rect 4712 15444 4764 15453
rect 5540 15487 5592 15496
rect 5540 15453 5549 15487
rect 5549 15453 5583 15487
rect 5583 15453 5592 15487
rect 5540 15444 5592 15453
rect 6184 15648 6236 15700
rect 10416 15648 10468 15700
rect 10876 15648 10928 15700
rect 8300 15580 8352 15632
rect 7196 15512 7248 15564
rect 8116 15512 8168 15564
rect 9772 15512 9824 15564
rect 10324 15512 10376 15564
rect 7472 15444 7524 15496
rect 8208 15487 8260 15496
rect 8208 15453 8217 15487
rect 8217 15453 8251 15487
rect 8251 15453 8260 15487
rect 8208 15444 8260 15453
rect 5356 15376 5408 15428
rect 7656 15376 7708 15428
rect 7840 15376 7892 15428
rect 8576 15376 8628 15428
rect 11244 15580 11296 15632
rect 11704 15555 11756 15564
rect 11704 15521 11713 15555
rect 11713 15521 11747 15555
rect 11747 15521 11756 15555
rect 11704 15512 11756 15521
rect 12808 15648 12860 15700
rect 14096 15691 14148 15700
rect 14096 15657 14105 15691
rect 14105 15657 14139 15691
rect 14139 15657 14148 15691
rect 14096 15648 14148 15657
rect 15292 15648 15344 15700
rect 18052 15648 18104 15700
rect 18788 15691 18840 15700
rect 18788 15657 18797 15691
rect 18797 15657 18831 15691
rect 18831 15657 18840 15691
rect 18788 15648 18840 15657
rect 20904 15648 20956 15700
rect 16212 15580 16264 15632
rect 14464 15512 14516 15564
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 12808 15487 12860 15496
rect 11888 15444 11940 15453
rect 12808 15453 12817 15487
rect 12817 15453 12851 15487
rect 12851 15453 12860 15487
rect 12808 15444 12860 15453
rect 12992 15487 13044 15496
rect 12992 15453 13001 15487
rect 13001 15453 13035 15487
rect 13035 15453 13044 15487
rect 12992 15444 13044 15453
rect 13268 15444 13320 15496
rect 14556 15487 14608 15496
rect 14556 15453 14565 15487
rect 14565 15453 14599 15487
rect 14599 15453 14608 15487
rect 14556 15444 14608 15453
rect 16028 15512 16080 15564
rect 16488 15512 16540 15564
rect 16396 15487 16448 15496
rect 16396 15453 16405 15487
rect 16405 15453 16439 15487
rect 16439 15453 16448 15487
rect 16396 15444 16448 15453
rect 4712 15308 4764 15360
rect 4896 15308 4948 15360
rect 5540 15308 5592 15360
rect 11612 15308 11664 15360
rect 15476 15376 15528 15428
rect 17500 15512 17552 15564
rect 18604 15512 18656 15564
rect 19064 15512 19116 15564
rect 20168 15555 20220 15564
rect 16672 15444 16724 15496
rect 17592 15444 17644 15496
rect 18696 15444 18748 15496
rect 19248 15487 19300 15496
rect 19248 15453 19257 15487
rect 19257 15453 19291 15487
rect 19291 15453 19300 15487
rect 19248 15444 19300 15453
rect 20168 15521 20177 15555
rect 20177 15521 20211 15555
rect 20211 15521 20220 15555
rect 20168 15512 20220 15521
rect 20260 15487 20312 15496
rect 18512 15376 18564 15428
rect 19156 15376 19208 15428
rect 20260 15453 20269 15487
rect 20269 15453 20303 15487
rect 20303 15453 20312 15487
rect 20260 15444 20312 15453
rect 16304 15308 16356 15360
rect 17316 15308 17368 15360
rect 19616 15308 19668 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 7288 15104 7340 15156
rect 7656 15104 7708 15156
rect 7840 15147 7892 15156
rect 7840 15113 7849 15147
rect 7849 15113 7883 15147
rect 7883 15113 7892 15147
rect 7840 15104 7892 15113
rect 3700 15036 3752 15088
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 2228 15011 2280 15020
rect 2228 14977 2237 15011
rect 2237 14977 2271 15011
rect 2271 14977 2280 15011
rect 2228 14968 2280 14977
rect 5816 14968 5868 15020
rect 7748 14968 7800 15020
rect 9956 15104 10008 15156
rect 11704 15104 11756 15156
rect 12808 15104 12860 15156
rect 14280 15147 14332 15156
rect 14280 15113 14289 15147
rect 14289 15113 14323 15147
rect 14323 15113 14332 15147
rect 14280 15104 14332 15113
rect 14556 15104 14608 15156
rect 14740 15104 14792 15156
rect 15568 15104 15620 15156
rect 17960 15104 18012 15156
rect 19432 15147 19484 15156
rect 19432 15113 19441 15147
rect 19441 15113 19475 15147
rect 19475 15113 19484 15147
rect 19432 15104 19484 15113
rect 20260 15104 20312 15156
rect 20628 15104 20680 15156
rect 9864 14968 9916 15020
rect 10324 14968 10376 15020
rect 10876 14968 10928 15020
rect 8208 14900 8260 14952
rect 8300 14900 8352 14952
rect 12900 14968 12952 15020
rect 13176 14968 13228 15020
rect 13636 14968 13688 15020
rect 11612 14900 11664 14952
rect 13820 14900 13872 14952
rect 14740 14968 14792 15020
rect 15200 15011 15252 15020
rect 15200 14977 15209 15011
rect 15209 14977 15243 15011
rect 15243 14977 15252 15011
rect 15200 14968 15252 14977
rect 15844 14968 15896 15020
rect 3240 14832 3292 14884
rect 7564 14832 7616 14884
rect 9128 14832 9180 14884
rect 4804 14807 4856 14816
rect 4804 14773 4813 14807
rect 4813 14773 4847 14807
rect 4847 14773 4856 14807
rect 4804 14764 4856 14773
rect 5356 14764 5408 14816
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 7656 14764 7708 14816
rect 8852 14807 8904 14816
rect 8852 14773 8861 14807
rect 8861 14773 8895 14807
rect 8895 14773 8904 14807
rect 8852 14764 8904 14773
rect 12532 14832 12584 14884
rect 13728 14832 13780 14884
rect 17776 14900 17828 14952
rect 9772 14807 9824 14816
rect 9772 14773 9781 14807
rect 9781 14773 9815 14807
rect 9815 14773 9824 14807
rect 9772 14764 9824 14773
rect 10416 14764 10468 14816
rect 10876 14807 10928 14816
rect 10876 14773 10885 14807
rect 10885 14773 10919 14807
rect 10919 14773 10928 14807
rect 10876 14764 10928 14773
rect 12624 14807 12676 14816
rect 12624 14773 12633 14807
rect 12633 14773 12667 14807
rect 12667 14773 12676 14807
rect 12624 14764 12676 14773
rect 12992 14807 13044 14816
rect 12992 14773 13001 14807
rect 13001 14773 13035 14807
rect 13035 14773 13044 14807
rect 12992 14764 13044 14773
rect 15476 14764 15528 14816
rect 15844 14764 15896 14816
rect 16120 14764 16172 14816
rect 16396 14832 16448 14884
rect 17500 14832 17552 14884
rect 18512 14832 18564 14884
rect 19708 14832 19760 14884
rect 16856 14764 16908 14816
rect 17408 14807 17460 14816
rect 17408 14773 17417 14807
rect 17417 14773 17451 14807
rect 17451 14773 17460 14807
rect 17408 14764 17460 14773
rect 17960 14764 18012 14816
rect 19340 14764 19392 14816
rect 20352 14764 20404 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 4160 14560 4212 14612
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 7104 14560 7156 14612
rect 1860 14424 1912 14476
rect 2412 14424 2464 14476
rect 2872 14424 2924 14476
rect 3700 14356 3752 14408
rect 4252 14424 4304 14476
rect 5080 14424 5132 14476
rect 7564 14492 7616 14544
rect 8300 14560 8352 14612
rect 9680 14560 9732 14612
rect 9772 14560 9824 14612
rect 12532 14560 12584 14612
rect 12624 14560 12676 14612
rect 15660 14560 15712 14612
rect 16396 14603 16448 14612
rect 16396 14569 16405 14603
rect 16405 14569 16439 14603
rect 16439 14569 16448 14603
rect 16396 14560 16448 14569
rect 18512 14560 18564 14612
rect 18696 14560 18748 14612
rect 18972 14603 19024 14612
rect 18972 14569 18981 14603
rect 18981 14569 19015 14603
rect 19015 14569 19024 14603
rect 18972 14560 19024 14569
rect 19616 14603 19668 14612
rect 19616 14569 19625 14603
rect 19625 14569 19659 14603
rect 19659 14569 19668 14603
rect 19616 14560 19668 14569
rect 5540 14424 5592 14476
rect 9128 14492 9180 14544
rect 10140 14492 10192 14544
rect 12716 14492 12768 14544
rect 16304 14535 16356 14544
rect 16304 14501 16313 14535
rect 16313 14501 16347 14535
rect 16347 14501 16356 14535
rect 16304 14492 16356 14501
rect 17408 14492 17460 14544
rect 9772 14424 9824 14476
rect 9956 14424 10008 14476
rect 12532 14467 12584 14476
rect 7748 14356 7800 14408
rect 8852 14356 8904 14408
rect 10232 14399 10284 14408
rect 10232 14365 10241 14399
rect 10241 14365 10275 14399
rect 10275 14365 10284 14399
rect 10232 14356 10284 14365
rect 10508 14356 10560 14408
rect 12532 14433 12566 14467
rect 12566 14433 12584 14467
rect 12532 14424 12584 14433
rect 14004 14424 14056 14476
rect 15016 14424 15068 14476
rect 12256 14399 12308 14408
rect 12256 14365 12265 14399
rect 12265 14365 12299 14399
rect 12299 14365 12308 14399
rect 12256 14356 12308 14365
rect 13728 14288 13780 14340
rect 14556 14288 14608 14340
rect 7564 14220 7616 14272
rect 7748 14263 7800 14272
rect 7748 14229 7757 14263
rect 7757 14229 7791 14263
rect 7791 14229 7800 14263
rect 7748 14220 7800 14229
rect 10968 14220 11020 14272
rect 11704 14220 11756 14272
rect 13636 14263 13688 14272
rect 13636 14229 13645 14263
rect 13645 14229 13679 14263
rect 13679 14229 13688 14263
rect 13636 14220 13688 14229
rect 15108 14220 15160 14272
rect 16488 14424 16540 14476
rect 18788 14424 18840 14476
rect 16948 14399 17000 14408
rect 16948 14365 16957 14399
rect 16957 14365 16991 14399
rect 16991 14365 17000 14399
rect 16948 14356 17000 14365
rect 20628 14424 20680 14476
rect 19340 14356 19392 14408
rect 16672 14288 16724 14340
rect 18880 14288 18932 14340
rect 19984 14220 20036 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 2780 14016 2832 14068
rect 3148 14059 3200 14068
rect 3148 14025 3157 14059
rect 3157 14025 3191 14059
rect 3191 14025 3200 14059
rect 3148 14016 3200 14025
rect 3516 14016 3568 14068
rect 5080 14059 5132 14068
rect 5080 14025 5089 14059
rect 5089 14025 5123 14059
rect 5123 14025 5132 14059
rect 5080 14016 5132 14025
rect 5356 14059 5408 14068
rect 5356 14025 5365 14059
rect 5365 14025 5399 14059
rect 5399 14025 5408 14059
rect 5356 14016 5408 14025
rect 8668 14059 8720 14068
rect 8668 14025 8677 14059
rect 8677 14025 8711 14059
rect 8711 14025 8720 14059
rect 8668 14016 8720 14025
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 5080 13880 5132 13932
rect 6000 13880 6052 13932
rect 10876 14016 10928 14068
rect 13084 14016 13136 14068
rect 15016 14059 15068 14068
rect 9588 13880 9640 13932
rect 10140 13923 10192 13932
rect 10140 13889 10149 13923
rect 10149 13889 10183 13923
rect 10183 13889 10192 13923
rect 10140 13880 10192 13889
rect 10232 13923 10284 13932
rect 10232 13889 10241 13923
rect 10241 13889 10275 13923
rect 10275 13889 10284 13923
rect 10968 13923 11020 13932
rect 10232 13880 10284 13889
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 14556 13948 14608 14000
rect 15016 14025 15025 14059
rect 15025 14025 15059 14059
rect 15059 14025 15068 14059
rect 15016 14016 15068 14025
rect 15108 14016 15160 14068
rect 17868 14016 17920 14068
rect 17960 14016 18012 14068
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 2412 13855 2464 13864
rect 2412 13821 2421 13855
rect 2421 13821 2455 13855
rect 2455 13821 2464 13855
rect 2412 13812 2464 13821
rect 2964 13855 3016 13864
rect 2964 13821 2973 13855
rect 2973 13821 3007 13855
rect 3007 13821 3016 13855
rect 2964 13812 3016 13821
rect 4252 13812 4304 13864
rect 6828 13812 6880 13864
rect 7288 13855 7340 13864
rect 7288 13821 7297 13855
rect 7297 13821 7331 13855
rect 7331 13821 7340 13855
rect 7288 13812 7340 13821
rect 7564 13855 7616 13864
rect 7564 13821 7598 13855
rect 7598 13821 7616 13855
rect 7564 13812 7616 13821
rect 8944 13812 8996 13864
rect 10324 13812 10376 13864
rect 12256 13880 12308 13932
rect 13636 13855 13688 13864
rect 13636 13821 13670 13855
rect 13670 13821 13688 13855
rect 16396 13880 16448 13932
rect 17500 13923 17552 13932
rect 17500 13889 17509 13923
rect 17509 13889 17543 13923
rect 17543 13889 17552 13923
rect 17500 13880 17552 13889
rect 13636 13812 13688 13821
rect 16304 13812 16356 13864
rect 17132 13812 17184 13864
rect 17224 13855 17276 13864
rect 17224 13821 17233 13855
rect 17233 13821 17267 13855
rect 17267 13821 17276 13855
rect 17224 13812 17276 13821
rect 3976 13787 4028 13796
rect 3976 13753 4010 13787
rect 4010 13753 4028 13787
rect 3976 13744 4028 13753
rect 5540 13744 5592 13796
rect 8852 13744 8904 13796
rect 9588 13744 9640 13796
rect 7748 13676 7800 13728
rect 9220 13719 9272 13728
rect 9220 13685 9229 13719
rect 9229 13685 9263 13719
rect 9263 13685 9272 13719
rect 9220 13676 9272 13685
rect 14372 13744 14424 13796
rect 15016 13744 15068 13796
rect 15936 13744 15988 13796
rect 17868 13744 17920 13796
rect 19248 14016 19300 14068
rect 18236 13991 18288 14000
rect 18236 13957 18245 13991
rect 18245 13957 18279 13991
rect 18279 13957 18288 13991
rect 18236 13948 18288 13957
rect 19708 13880 19760 13932
rect 19432 13812 19484 13864
rect 20444 13812 20496 13864
rect 10140 13676 10192 13728
rect 10508 13676 10560 13728
rect 10784 13676 10836 13728
rect 11796 13719 11848 13728
rect 11796 13685 11805 13719
rect 11805 13685 11839 13719
rect 11839 13685 11848 13719
rect 11796 13676 11848 13685
rect 12900 13676 12952 13728
rect 15200 13676 15252 13728
rect 15292 13676 15344 13728
rect 16304 13676 16356 13728
rect 16488 13676 16540 13728
rect 17776 13676 17828 13728
rect 18604 13676 18656 13728
rect 18972 13676 19024 13728
rect 19248 13676 19300 13728
rect 19892 13676 19944 13728
rect 20260 13719 20312 13728
rect 20260 13685 20269 13719
rect 20269 13685 20303 13719
rect 20303 13685 20312 13719
rect 20260 13676 20312 13685
rect 20720 13676 20772 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 1768 13515 1820 13524
rect 1768 13481 1777 13515
rect 1777 13481 1811 13515
rect 1811 13481 1820 13515
rect 1768 13472 1820 13481
rect 6092 13472 6144 13524
rect 9404 13472 9456 13524
rect 9864 13472 9916 13524
rect 12992 13515 13044 13524
rect 2964 13404 3016 13456
rect 4712 13404 4764 13456
rect 5356 13404 5408 13456
rect 6644 13404 6696 13456
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 4160 13336 4212 13388
rect 4252 13336 4304 13388
rect 6276 13336 6328 13388
rect 4712 13268 4764 13320
rect 5540 13268 5592 13320
rect 5908 13311 5960 13320
rect 5908 13277 5917 13311
rect 5917 13277 5951 13311
rect 5951 13277 5960 13311
rect 5908 13268 5960 13277
rect 6000 13311 6052 13320
rect 6000 13277 6009 13311
rect 6009 13277 6043 13311
rect 6043 13277 6052 13311
rect 7564 13336 7616 13388
rect 8668 13404 8720 13456
rect 10140 13336 10192 13388
rect 11336 13336 11388 13388
rect 12992 13481 13001 13515
rect 13001 13481 13035 13515
rect 13035 13481 13044 13515
rect 12992 13472 13044 13481
rect 13176 13472 13228 13524
rect 15292 13515 15344 13524
rect 15292 13481 15301 13515
rect 15301 13481 15335 13515
rect 15335 13481 15344 13515
rect 15292 13472 15344 13481
rect 15752 13515 15804 13524
rect 15752 13481 15761 13515
rect 15761 13481 15795 13515
rect 15795 13481 15804 13515
rect 15752 13472 15804 13481
rect 16028 13472 16080 13524
rect 16396 13472 16448 13524
rect 20536 13472 20588 13524
rect 15200 13404 15252 13456
rect 12716 13336 12768 13388
rect 6000 13268 6052 13277
rect 7288 13268 7340 13320
rect 9128 13268 9180 13320
rect 4804 13200 4856 13252
rect 8852 13243 8904 13252
rect 8852 13209 8861 13243
rect 8861 13209 8895 13243
rect 8895 13209 8904 13243
rect 8852 13200 8904 13209
rect 7656 13132 7708 13184
rect 12532 13268 12584 13320
rect 14464 13311 14516 13320
rect 12900 13243 12952 13252
rect 12900 13209 12909 13243
rect 12909 13209 12943 13243
rect 12943 13209 12952 13243
rect 12900 13200 12952 13209
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 14556 13268 14608 13320
rect 15016 13336 15068 13388
rect 19892 13404 19944 13456
rect 16120 13268 16172 13320
rect 12256 13132 12308 13184
rect 13728 13132 13780 13184
rect 13912 13132 13964 13184
rect 14280 13132 14332 13184
rect 14924 13132 14976 13184
rect 17776 13336 17828 13388
rect 18236 13379 18288 13388
rect 18236 13345 18270 13379
rect 18270 13345 18288 13379
rect 18236 13336 18288 13345
rect 19616 13336 19668 13388
rect 18972 13268 19024 13320
rect 20812 13200 20864 13252
rect 19432 13132 19484 13184
rect 19708 13132 19760 13184
rect 20536 13132 20588 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 1676 12928 1728 12980
rect 3976 12928 4028 12980
rect 5908 12928 5960 12980
rect 9220 12928 9272 12980
rect 9680 12928 9732 12980
rect 10876 12928 10928 12980
rect 14004 12928 14056 12980
rect 3516 12860 3568 12912
rect 13176 12860 13228 12912
rect 17224 12928 17276 12980
rect 18972 12971 19024 12980
rect 18972 12937 18981 12971
rect 18981 12937 19015 12971
rect 19015 12937 19024 12971
rect 18972 12928 19024 12937
rect 4252 12835 4304 12844
rect 1492 12724 1544 12776
rect 4252 12801 4261 12835
rect 4261 12801 4295 12835
rect 4295 12801 4304 12835
rect 4252 12792 4304 12801
rect 5540 12792 5592 12844
rect 6184 12835 6236 12844
rect 6184 12801 6193 12835
rect 6193 12801 6227 12835
rect 6227 12801 6236 12835
rect 6184 12792 6236 12801
rect 6368 12835 6420 12844
rect 6368 12801 6377 12835
rect 6377 12801 6411 12835
rect 6411 12801 6420 12835
rect 6368 12792 6420 12801
rect 7656 12835 7708 12844
rect 7656 12801 7665 12835
rect 7665 12801 7699 12835
rect 7699 12801 7708 12835
rect 7656 12792 7708 12801
rect 8668 12792 8720 12844
rect 8944 12792 8996 12844
rect 9404 12792 9456 12844
rect 12256 12792 12308 12844
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 2780 12767 2832 12776
rect 2780 12733 2803 12767
rect 2803 12733 2832 12767
rect 2780 12724 2832 12733
rect 4896 12724 4948 12776
rect 5356 12656 5408 12708
rect 1860 12631 1912 12640
rect 1860 12597 1869 12631
rect 1869 12597 1903 12631
rect 1903 12597 1912 12631
rect 1860 12588 1912 12597
rect 1952 12631 2004 12640
rect 1952 12597 1961 12631
rect 1961 12597 1995 12631
rect 1995 12597 2004 12631
rect 5080 12631 5132 12640
rect 1952 12588 2004 12597
rect 5080 12597 5089 12631
rect 5089 12597 5123 12631
rect 5123 12597 5132 12631
rect 5080 12588 5132 12597
rect 6000 12588 6052 12640
rect 6092 12631 6144 12640
rect 6092 12597 6101 12631
rect 6101 12597 6135 12631
rect 6135 12597 6144 12631
rect 6092 12588 6144 12597
rect 13636 12724 13688 12776
rect 15384 12792 15436 12844
rect 15844 12860 15896 12912
rect 17960 12860 18012 12912
rect 18052 12860 18104 12912
rect 18880 12860 18932 12912
rect 19064 12860 19116 12912
rect 20352 12860 20404 12912
rect 21088 12860 21140 12912
rect 16580 12792 16632 12844
rect 17040 12792 17092 12844
rect 17224 12792 17276 12844
rect 17500 12835 17552 12844
rect 17500 12801 17509 12835
rect 17509 12801 17543 12835
rect 17543 12801 17552 12835
rect 17500 12792 17552 12801
rect 18604 12792 18656 12844
rect 19432 12792 19484 12844
rect 20168 12792 20220 12844
rect 20536 12835 20588 12844
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 10140 12656 10192 12708
rect 14832 12724 14884 12776
rect 16120 12724 16172 12776
rect 16396 12767 16448 12776
rect 16396 12733 16405 12767
rect 16405 12733 16439 12767
rect 16439 12733 16448 12767
rect 16396 12724 16448 12733
rect 15108 12656 15160 12708
rect 8760 12588 8812 12640
rect 13912 12588 13964 12640
rect 15936 12631 15988 12640
rect 15936 12597 15945 12631
rect 15945 12597 15979 12631
rect 15979 12597 15988 12631
rect 15936 12588 15988 12597
rect 20260 12724 20312 12776
rect 17316 12699 17368 12708
rect 17316 12665 17325 12699
rect 17325 12665 17359 12699
rect 17359 12665 17368 12699
rect 17316 12656 17368 12665
rect 19524 12656 19576 12708
rect 17040 12588 17092 12640
rect 19984 12631 20036 12640
rect 19984 12597 19993 12631
rect 19993 12597 20027 12631
rect 20027 12597 20036 12631
rect 19984 12588 20036 12597
rect 20904 12656 20956 12708
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2780 12384 2832 12436
rect 4252 12384 4304 12436
rect 7104 12384 7156 12436
rect 8208 12384 8260 12436
rect 8760 12384 8812 12436
rect 10324 12384 10376 12436
rect 10692 12384 10744 12436
rect 12532 12384 12584 12436
rect 13636 12384 13688 12436
rect 15016 12384 15068 12436
rect 15200 12384 15252 12436
rect 17500 12384 17552 12436
rect 19616 12427 19668 12436
rect 19616 12393 19625 12427
rect 19625 12393 19659 12427
rect 19659 12393 19668 12427
rect 19616 12384 19668 12393
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 20904 12427 20956 12436
rect 20904 12393 20913 12427
rect 20913 12393 20947 12427
rect 20947 12393 20956 12427
rect 20904 12384 20956 12393
rect 4068 12316 4120 12368
rect 15752 12316 15804 12368
rect 17408 12316 17460 12368
rect 17592 12316 17644 12368
rect 17776 12316 17828 12368
rect 20444 12316 20496 12368
rect 2688 12248 2740 12300
rect 5264 12248 5316 12300
rect 1492 12180 1544 12232
rect 4252 12180 4304 12232
rect 4804 12044 4856 12096
rect 9220 12248 9272 12300
rect 10140 12248 10192 12300
rect 10416 12248 10468 12300
rect 10600 12291 10652 12300
rect 10600 12257 10609 12291
rect 10609 12257 10643 12291
rect 10643 12257 10652 12291
rect 10600 12248 10652 12257
rect 10784 12248 10836 12300
rect 7748 12223 7800 12232
rect 7748 12189 7757 12223
rect 7757 12189 7791 12223
rect 7791 12189 7800 12223
rect 7748 12180 7800 12189
rect 8760 12180 8812 12232
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 12348 12248 12400 12300
rect 11152 12180 11204 12232
rect 5908 12044 5960 12096
rect 14464 12248 14516 12300
rect 17316 12248 17368 12300
rect 12900 12223 12952 12232
rect 12900 12189 12909 12223
rect 12909 12189 12943 12223
rect 12943 12189 12952 12223
rect 12900 12180 12952 12189
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 14464 12112 14516 12164
rect 15016 12112 15068 12164
rect 15384 12112 15436 12164
rect 16120 12180 16172 12232
rect 17500 12180 17552 12232
rect 20536 12248 20588 12300
rect 19708 12180 19760 12232
rect 20168 12223 20220 12232
rect 20168 12189 20177 12223
rect 20177 12189 20211 12223
rect 20211 12189 20220 12223
rect 20168 12180 20220 12189
rect 8944 12044 8996 12096
rect 14556 12044 14608 12096
rect 16856 12044 16908 12096
rect 19156 12044 19208 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 1952 11840 2004 11892
rect 4160 11883 4212 11892
rect 4160 11849 4169 11883
rect 4169 11849 4203 11883
rect 4203 11849 4212 11883
rect 4160 11840 4212 11849
rect 2688 11747 2740 11756
rect 2688 11713 2697 11747
rect 2697 11713 2731 11747
rect 2731 11713 2740 11747
rect 2688 11704 2740 11713
rect 4804 11747 4856 11756
rect 3516 11679 3568 11688
rect 3516 11645 3525 11679
rect 3525 11645 3559 11679
rect 3559 11645 3568 11679
rect 3516 11636 3568 11645
rect 4804 11713 4813 11747
rect 4813 11713 4847 11747
rect 4847 11713 4856 11747
rect 4804 11704 4856 11713
rect 5356 11704 5408 11756
rect 4068 11636 4120 11688
rect 5908 11636 5960 11688
rect 7104 11636 7156 11688
rect 12440 11840 12492 11892
rect 12532 11840 12584 11892
rect 9220 11772 9272 11824
rect 14280 11840 14332 11892
rect 16672 11840 16724 11892
rect 19248 11840 19300 11892
rect 10600 11747 10652 11756
rect 10600 11713 10609 11747
rect 10609 11713 10643 11747
rect 10643 11713 10652 11747
rect 10600 11704 10652 11713
rect 10784 11704 10836 11756
rect 7748 11636 7800 11688
rect 8116 11636 8168 11688
rect 8852 11636 8904 11688
rect 9036 11636 9088 11688
rect 10692 11636 10744 11688
rect 11980 11704 12032 11756
rect 12900 11704 12952 11756
rect 3700 11568 3752 11620
rect 3792 11568 3844 11620
rect 4252 11500 4304 11552
rect 5540 11543 5592 11552
rect 5540 11509 5549 11543
rect 5549 11509 5583 11543
rect 5583 11509 5592 11543
rect 5540 11500 5592 11509
rect 6276 11500 6328 11552
rect 6460 11543 6512 11552
rect 6460 11509 6469 11543
rect 6469 11509 6503 11543
rect 6503 11509 6512 11543
rect 6460 11500 6512 11509
rect 12072 11636 12124 11688
rect 12256 11636 12308 11688
rect 13636 11636 13688 11688
rect 13728 11636 13780 11688
rect 15016 11704 15068 11756
rect 17684 11772 17736 11824
rect 15936 11636 15988 11688
rect 8944 11500 8996 11552
rect 9128 11500 9180 11552
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 10416 11500 10468 11552
rect 11612 11568 11664 11620
rect 13820 11568 13872 11620
rect 11336 11500 11388 11552
rect 14372 11500 14424 11552
rect 15016 11568 15068 11620
rect 16580 11636 16632 11688
rect 18420 11679 18472 11688
rect 18420 11645 18429 11679
rect 18429 11645 18463 11679
rect 18463 11645 18472 11679
rect 18420 11636 18472 11645
rect 19984 11636 20036 11688
rect 15292 11500 15344 11552
rect 16120 11568 16172 11620
rect 16856 11568 16908 11620
rect 17132 11568 17184 11620
rect 20536 11568 20588 11620
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 18880 11500 18932 11552
rect 19524 11500 19576 11552
rect 20168 11500 20220 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2688 11296 2740 11348
rect 5448 11296 5500 11348
rect 5540 11296 5592 11348
rect 6000 11296 6052 11348
rect 6276 11296 6328 11348
rect 7012 11296 7064 11348
rect 8760 11296 8812 11348
rect 9036 11296 9088 11348
rect 1492 11228 1544 11280
rect 2504 11160 2556 11212
rect 4160 11228 4212 11280
rect 5908 11228 5960 11280
rect 9588 11228 9640 11280
rect 10048 11228 10100 11280
rect 11152 11228 11204 11280
rect 13728 11296 13780 11348
rect 15108 11296 15160 11348
rect 16856 11296 16908 11348
rect 17592 11296 17644 11348
rect 17776 11296 17828 11348
rect 18420 11296 18472 11348
rect 18788 11296 18840 11348
rect 19340 11296 19392 11348
rect 20628 11296 20680 11348
rect 14372 11228 14424 11280
rect 4804 11160 4856 11212
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 5448 11160 5500 11212
rect 8208 11160 8260 11212
rect 10416 11160 10468 11212
rect 6920 11024 6972 11076
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 9864 11092 9916 11144
rect 10324 11092 10376 11144
rect 9312 11024 9364 11076
rect 9496 11024 9548 11076
rect 11612 11092 11664 11144
rect 12348 11092 12400 11144
rect 12808 11135 12860 11144
rect 12808 11101 12817 11135
rect 12817 11101 12851 11135
rect 12851 11101 12860 11135
rect 12808 11092 12860 11101
rect 11244 11024 11296 11076
rect 11980 11067 12032 11076
rect 11980 11033 11989 11067
rect 11989 11033 12023 11067
rect 12023 11033 12032 11067
rect 11980 11024 12032 11033
rect 12900 11024 12952 11076
rect 14004 11160 14056 11212
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 13820 11135 13872 11144
rect 13820 11101 13829 11135
rect 13829 11101 13863 11135
rect 13863 11101 13872 11135
rect 13820 11092 13872 11101
rect 14556 11092 14608 11144
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 17684 11092 17736 11144
rect 17960 11092 18012 11144
rect 20076 11228 20128 11280
rect 14832 11024 14884 11076
rect 16580 11024 16632 11076
rect 19616 11092 19668 11144
rect 5356 10956 5408 11008
rect 8576 10999 8628 11008
rect 8576 10965 8585 10999
rect 8585 10965 8619 10999
rect 8619 10965 8628 10999
rect 8576 10956 8628 10965
rect 8668 10956 8720 11008
rect 9220 10956 9272 11008
rect 10600 10956 10652 11008
rect 14740 10956 14792 11008
rect 15200 10956 15252 11008
rect 16948 10999 17000 11008
rect 16948 10965 16957 10999
rect 16957 10965 16991 10999
rect 16991 10965 17000 10999
rect 16948 10956 17000 10965
rect 17868 10956 17920 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 1860 10752 1912 10804
rect 4252 10752 4304 10804
rect 4896 10752 4948 10804
rect 5264 10752 5316 10804
rect 10140 10752 10192 10804
rect 4344 10684 4396 10736
rect 4712 10684 4764 10736
rect 5172 10684 5224 10736
rect 2688 10616 2740 10668
rect 2504 10548 2556 10600
rect 3792 10616 3844 10668
rect 5356 10616 5408 10668
rect 6000 10616 6052 10668
rect 6368 10616 6420 10668
rect 7656 10616 7708 10668
rect 8576 10616 8628 10668
rect 9312 10616 9364 10668
rect 9404 10616 9456 10668
rect 11060 10752 11112 10804
rect 12348 10752 12400 10804
rect 14740 10752 14792 10804
rect 15016 10752 15068 10804
rect 15108 10752 15160 10804
rect 17408 10752 17460 10804
rect 18512 10752 18564 10804
rect 18880 10752 18932 10804
rect 19984 10752 20036 10804
rect 12532 10684 12584 10736
rect 16580 10684 16632 10736
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 4252 10548 4304 10600
rect 4896 10548 4948 10600
rect 6460 10548 6512 10600
rect 9772 10548 9824 10600
rect 1860 10412 1912 10464
rect 5172 10480 5224 10532
rect 3056 10455 3108 10464
rect 3056 10421 3065 10455
rect 3065 10421 3099 10455
rect 3099 10421 3108 10455
rect 3056 10412 3108 10421
rect 4068 10412 4120 10464
rect 4804 10412 4856 10464
rect 5264 10455 5316 10464
rect 5264 10421 5273 10455
rect 5273 10421 5307 10455
rect 5307 10421 5316 10455
rect 5264 10412 5316 10421
rect 8944 10480 8996 10532
rect 10784 10548 10836 10600
rect 10968 10591 11020 10600
rect 10968 10557 11002 10591
rect 11002 10557 11020 10591
rect 10968 10548 11020 10557
rect 12256 10548 12308 10600
rect 12348 10548 12400 10600
rect 13820 10616 13872 10668
rect 15384 10616 15436 10668
rect 15568 10616 15620 10668
rect 16856 10616 16908 10668
rect 17776 10616 17828 10668
rect 18880 10616 18932 10668
rect 19616 10616 19668 10668
rect 14096 10548 14148 10600
rect 14832 10591 14884 10600
rect 14832 10557 14841 10591
rect 14841 10557 14875 10591
rect 14875 10557 14884 10591
rect 14832 10548 14884 10557
rect 15016 10548 15068 10600
rect 15844 10548 15896 10600
rect 16948 10548 17000 10600
rect 18144 10548 18196 10600
rect 18696 10548 18748 10600
rect 19524 10548 19576 10600
rect 19708 10548 19760 10600
rect 7472 10412 7524 10464
rect 7748 10455 7800 10464
rect 7748 10421 7757 10455
rect 7757 10421 7791 10455
rect 7791 10421 7800 10455
rect 8300 10455 8352 10464
rect 7748 10412 7800 10421
rect 8300 10421 8309 10455
rect 8309 10421 8343 10455
rect 8343 10421 8352 10455
rect 8300 10412 8352 10421
rect 8576 10412 8628 10464
rect 11152 10480 11204 10532
rect 16764 10480 16816 10532
rect 17776 10480 17828 10532
rect 12532 10412 12584 10464
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 13360 10412 13412 10464
rect 14556 10412 14608 10464
rect 15568 10412 15620 10464
rect 16120 10455 16172 10464
rect 16120 10421 16129 10455
rect 16129 10421 16163 10455
rect 16163 10421 16172 10455
rect 16120 10412 16172 10421
rect 16212 10412 16264 10464
rect 18788 10412 18840 10464
rect 19432 10455 19484 10464
rect 19432 10421 19441 10455
rect 19441 10421 19475 10455
rect 19475 10421 19484 10455
rect 19432 10412 19484 10421
rect 20076 10480 20128 10532
rect 20720 10523 20772 10532
rect 20720 10489 20729 10523
rect 20729 10489 20763 10523
rect 20763 10489 20772 10523
rect 20720 10480 20772 10489
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 4068 10251 4120 10260
rect 4068 10217 4077 10251
rect 4077 10217 4111 10251
rect 4111 10217 4120 10251
rect 4068 10208 4120 10217
rect 4160 10208 4212 10260
rect 3056 10140 3108 10192
rect 4620 10140 4672 10192
rect 5540 10208 5592 10260
rect 7472 10251 7524 10260
rect 7472 10217 7481 10251
rect 7481 10217 7515 10251
rect 7515 10217 7524 10251
rect 7472 10208 7524 10217
rect 9312 10251 9364 10260
rect 9312 10217 9321 10251
rect 9321 10217 9355 10251
rect 9355 10217 9364 10251
rect 9312 10208 9364 10217
rect 9588 10208 9640 10260
rect 3332 10072 3384 10124
rect 4712 10072 4764 10124
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 2504 10047 2556 10056
rect 2504 10013 2513 10047
rect 2513 10013 2547 10047
rect 2547 10013 2556 10047
rect 2504 10004 2556 10013
rect 4160 10004 4212 10056
rect 4344 10004 4396 10056
rect 4620 10047 4672 10056
rect 4620 10013 4629 10047
rect 4629 10013 4663 10047
rect 4663 10013 4672 10047
rect 4620 10004 4672 10013
rect 3148 9936 3200 9988
rect 3976 9936 4028 9988
rect 6460 10140 6512 10192
rect 6000 10072 6052 10124
rect 5080 9868 5132 9920
rect 12624 10140 12676 10192
rect 12808 10208 12860 10260
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 16120 10208 16172 10260
rect 17960 10208 18012 10260
rect 18144 10251 18196 10260
rect 18144 10217 18153 10251
rect 18153 10217 18187 10251
rect 18187 10217 18196 10251
rect 18144 10208 18196 10217
rect 18972 10208 19024 10260
rect 13728 10140 13780 10192
rect 16396 10140 16448 10192
rect 17316 10140 17368 10192
rect 20076 10208 20128 10260
rect 20260 10208 20312 10260
rect 20812 10208 20864 10260
rect 7564 10072 7616 10124
rect 9128 10072 9180 10124
rect 10324 10072 10376 10124
rect 11060 10072 11112 10124
rect 11520 10115 11572 10124
rect 11520 10081 11543 10115
rect 11543 10081 11572 10115
rect 11520 10072 11572 10081
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 13636 10072 13688 10124
rect 15016 10072 15068 10124
rect 15292 10072 15344 10124
rect 9036 10004 9088 10056
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 15108 10004 15160 10056
rect 15200 10004 15252 10056
rect 16212 10072 16264 10124
rect 18420 10072 18472 10124
rect 19616 10140 19668 10192
rect 16304 10047 16356 10056
rect 16304 10013 16313 10047
rect 16313 10013 16347 10047
rect 16347 10013 16356 10047
rect 16304 10004 16356 10013
rect 11244 9936 11296 9988
rect 12256 9936 12308 9988
rect 8576 9868 8628 9920
rect 8668 9868 8720 9920
rect 11612 9868 11664 9920
rect 12348 9868 12400 9920
rect 14188 9911 14240 9920
rect 14188 9877 14197 9911
rect 14197 9877 14231 9911
rect 14231 9877 14240 9911
rect 14188 9868 14240 9877
rect 18696 10004 18748 10056
rect 19340 10072 19392 10124
rect 19984 10072 20036 10124
rect 19524 10004 19576 10056
rect 20352 10047 20404 10056
rect 20352 10013 20361 10047
rect 20361 10013 20395 10047
rect 20395 10013 20404 10047
rect 20352 10004 20404 10013
rect 17684 9979 17736 9988
rect 17684 9945 17693 9979
rect 17693 9945 17727 9979
rect 17727 9945 17736 9979
rect 17684 9936 17736 9945
rect 18880 9936 18932 9988
rect 18512 9911 18564 9920
rect 18512 9877 18521 9911
rect 18521 9877 18555 9911
rect 18555 9877 18564 9911
rect 18512 9868 18564 9877
rect 20076 9868 20128 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 2320 9664 2372 9716
rect 6092 9664 6144 9716
rect 6644 9664 6696 9716
rect 1584 9528 1636 9580
rect 3792 9528 3844 9580
rect 2228 9460 2280 9512
rect 1584 9392 1636 9444
rect 4804 9460 4856 9512
rect 5540 9528 5592 9580
rect 6000 9571 6052 9580
rect 6000 9537 6009 9571
rect 6009 9537 6043 9571
rect 6043 9537 6052 9571
rect 6000 9528 6052 9537
rect 8576 9664 8628 9716
rect 10692 9664 10744 9716
rect 11796 9664 11848 9716
rect 14188 9664 14240 9716
rect 16212 9707 16264 9716
rect 12716 9596 12768 9648
rect 16212 9673 16221 9707
rect 16221 9673 16255 9707
rect 16255 9673 16264 9707
rect 16212 9664 16264 9673
rect 17224 9664 17276 9716
rect 17408 9664 17460 9716
rect 20168 9664 20220 9716
rect 8576 9528 8628 9580
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 13268 9528 13320 9580
rect 7380 9460 7432 9512
rect 7656 9460 7708 9512
rect 8392 9460 8444 9512
rect 9588 9460 9640 9512
rect 11612 9460 11664 9512
rect 2872 9392 2924 9444
rect 4068 9392 4120 9444
rect 11520 9392 11572 9444
rect 11796 9392 11848 9444
rect 13636 9460 13688 9512
rect 16396 9596 16448 9648
rect 18512 9596 18564 9648
rect 14556 9528 14608 9580
rect 16948 9528 17000 9580
rect 18696 9596 18748 9648
rect 19708 9596 19760 9648
rect 20260 9596 20312 9648
rect 21364 9596 21416 9648
rect 18972 9528 19024 9580
rect 19892 9528 19944 9580
rect 20352 9528 20404 9580
rect 18696 9460 18748 9512
rect 19340 9460 19392 9512
rect 20168 9460 20220 9512
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 15016 9392 15068 9444
rect 4252 9324 4304 9376
rect 5724 9367 5776 9376
rect 5724 9333 5733 9367
rect 5733 9333 5767 9367
rect 5767 9333 5776 9367
rect 5724 9324 5776 9333
rect 6736 9324 6788 9376
rect 9956 9324 10008 9376
rect 10968 9324 11020 9376
rect 12532 9324 12584 9376
rect 12808 9367 12860 9376
rect 12808 9333 12817 9367
rect 12817 9333 12851 9367
rect 12851 9333 12860 9367
rect 12808 9324 12860 9333
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 19432 9392 19484 9444
rect 16488 9367 16540 9376
rect 16488 9333 16497 9367
rect 16497 9333 16531 9367
rect 16531 9333 16540 9367
rect 16488 9324 16540 9333
rect 16672 9324 16724 9376
rect 19340 9324 19392 9376
rect 19524 9367 19576 9376
rect 19524 9333 19533 9367
rect 19533 9333 19567 9367
rect 19567 9333 19576 9367
rect 19524 9324 19576 9333
rect 19708 9324 19760 9376
rect 20168 9367 20220 9376
rect 20168 9333 20177 9367
rect 20177 9333 20211 9367
rect 20211 9333 20220 9367
rect 20168 9324 20220 9333
rect 20536 9367 20588 9376
rect 20536 9333 20545 9367
rect 20545 9333 20579 9367
rect 20579 9333 20588 9367
rect 20536 9324 20588 9333
rect 20628 9324 20680 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2228 9163 2280 9172
rect 2228 9129 2237 9163
rect 2237 9129 2271 9163
rect 2271 9129 2280 9163
rect 2228 9120 2280 9129
rect 4712 9120 4764 9172
rect 4896 9120 4948 9172
rect 5448 9163 5500 9172
rect 5448 9129 5457 9163
rect 5457 9129 5491 9163
rect 5491 9129 5500 9163
rect 5448 9120 5500 9129
rect 7748 9120 7800 9172
rect 8208 9120 8260 9172
rect 9864 9120 9916 9172
rect 10140 9163 10192 9172
rect 10140 9129 10149 9163
rect 10149 9129 10183 9163
rect 10183 9129 10192 9163
rect 10140 9120 10192 9129
rect 12900 9120 12952 9172
rect 13084 9120 13136 9172
rect 3332 9052 3384 9104
rect 4252 9052 4304 9104
rect 5080 9052 5132 9104
rect 5356 9052 5408 9104
rect 7380 9052 7432 9104
rect 8944 9052 8996 9104
rect 10876 9052 10928 9104
rect 15016 9120 15068 9172
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 15292 9120 15344 9129
rect 16488 9120 16540 9172
rect 17776 9120 17828 9172
rect 20536 9120 20588 9172
rect 16948 9052 17000 9104
rect 2596 9027 2648 9036
rect 2596 8993 2605 9027
rect 2605 8993 2639 9027
rect 2639 8993 2648 9027
rect 2596 8984 2648 8993
rect 5724 8984 5776 9036
rect 6184 8984 6236 9036
rect 6552 8984 6604 9036
rect 7288 8984 7340 9036
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 3700 8916 3752 8968
rect 4804 8916 4856 8968
rect 6000 8916 6052 8968
rect 3148 8848 3200 8900
rect 4068 8848 4120 8900
rect 7196 8916 7248 8968
rect 7932 8984 7984 9036
rect 9496 8984 9548 9036
rect 9956 8984 10008 9036
rect 7656 8959 7708 8968
rect 7656 8925 7665 8959
rect 7665 8925 7699 8959
rect 7699 8925 7708 8959
rect 7656 8916 7708 8925
rect 9036 8916 9088 8968
rect 9128 8916 9180 8968
rect 10140 8916 10192 8968
rect 10324 8984 10376 9036
rect 12900 8984 12952 9036
rect 13636 8984 13688 9036
rect 15752 8959 15804 8968
rect 5356 8780 5408 8832
rect 10508 8848 10560 8900
rect 11060 8848 11112 8900
rect 11796 8780 11848 8832
rect 12256 8780 12308 8832
rect 15752 8925 15761 8959
rect 15761 8925 15795 8959
rect 15795 8925 15804 8959
rect 15752 8916 15804 8925
rect 15016 8848 15068 8900
rect 15292 8780 15344 8832
rect 17132 8984 17184 9036
rect 17592 8984 17644 9036
rect 16948 8959 17000 8968
rect 16948 8925 16957 8959
rect 16957 8925 16991 8959
rect 16991 8925 17000 8959
rect 16948 8916 17000 8925
rect 16672 8848 16724 8900
rect 17868 9052 17920 9104
rect 19432 9052 19484 9104
rect 19616 9052 19668 9104
rect 19340 8984 19392 9036
rect 17868 8916 17920 8968
rect 19892 8780 19944 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 3148 8619 3200 8628
rect 3148 8585 3157 8619
rect 3157 8585 3191 8619
rect 3191 8585 3200 8619
rect 3148 8576 3200 8585
rect 5356 8619 5408 8628
rect 5356 8585 5365 8619
rect 5365 8585 5399 8619
rect 5399 8585 5408 8619
rect 5356 8576 5408 8585
rect 5540 8576 5592 8628
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 5632 8440 5684 8492
rect 7104 8440 7156 8492
rect 1584 8372 1636 8424
rect 2688 8372 2740 8424
rect 8576 8415 8628 8424
rect 3516 8279 3568 8288
rect 3516 8245 3525 8279
rect 3525 8245 3559 8279
rect 3559 8245 3568 8279
rect 3516 8236 3568 8245
rect 5172 8304 5224 8356
rect 6828 8304 6880 8356
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 9588 8440 9640 8492
rect 12440 8576 12492 8628
rect 15200 8576 15252 8628
rect 15752 8619 15804 8628
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 19432 8619 19484 8628
rect 12164 8508 12216 8560
rect 7932 8347 7984 8356
rect 7932 8313 7941 8347
rect 7941 8313 7975 8347
rect 7975 8313 7984 8347
rect 7932 8304 7984 8313
rect 8484 8304 8536 8356
rect 9680 8304 9732 8356
rect 10968 8304 11020 8356
rect 12256 8440 12308 8492
rect 13452 8440 13504 8492
rect 12532 8372 12584 8424
rect 15016 8440 15068 8492
rect 16948 8440 17000 8492
rect 17500 8483 17552 8492
rect 17500 8449 17509 8483
rect 17509 8449 17543 8483
rect 17543 8449 17552 8483
rect 17500 8440 17552 8449
rect 19432 8585 19441 8619
rect 19441 8585 19475 8619
rect 19475 8585 19484 8619
rect 19432 8576 19484 8585
rect 19708 8619 19760 8628
rect 19708 8585 19717 8619
rect 19717 8585 19751 8619
rect 19751 8585 19760 8619
rect 19708 8576 19760 8585
rect 20996 8576 21048 8628
rect 19984 8508 20036 8560
rect 13636 8304 13688 8356
rect 16672 8372 16724 8424
rect 15292 8304 15344 8356
rect 15384 8304 15436 8356
rect 17408 8372 17460 8424
rect 17868 8372 17920 8424
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 20076 8415 20128 8424
rect 20076 8381 20085 8415
rect 20085 8381 20119 8415
rect 20119 8381 20128 8415
rect 20076 8372 20128 8381
rect 20720 8415 20772 8424
rect 20720 8381 20729 8415
rect 20729 8381 20763 8415
rect 20763 8381 20772 8415
rect 20720 8372 20772 8381
rect 17960 8304 18012 8356
rect 18328 8347 18380 8356
rect 18328 8313 18362 8347
rect 18362 8313 18380 8347
rect 18328 8304 18380 8313
rect 20352 8304 20404 8356
rect 5540 8236 5592 8288
rect 6000 8236 6052 8288
rect 9220 8236 9272 8288
rect 10692 8279 10744 8288
rect 10692 8245 10701 8279
rect 10701 8245 10735 8279
rect 10735 8245 10744 8279
rect 10692 8236 10744 8245
rect 11612 8279 11664 8288
rect 11612 8245 11621 8279
rect 11621 8245 11655 8279
rect 11655 8245 11664 8279
rect 11612 8236 11664 8245
rect 12900 8236 12952 8288
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 19892 8236 19944 8288
rect 20076 8236 20128 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 2596 8075 2648 8084
rect 2596 8041 2605 8075
rect 2605 8041 2639 8075
rect 2639 8041 2648 8075
rect 2596 8032 2648 8041
rect 3516 8032 3568 8084
rect 5080 8032 5132 8084
rect 1492 7964 1544 8016
rect 2964 7939 3016 7948
rect 2964 7905 2973 7939
rect 2973 7905 3007 7939
rect 3007 7905 3016 7939
rect 2964 7896 3016 7905
rect 4712 7896 4764 7948
rect 2688 7828 2740 7880
rect 3884 7828 3936 7880
rect 3976 7828 4028 7880
rect 6000 8032 6052 8084
rect 7104 8075 7156 8084
rect 7104 8041 7113 8075
rect 7113 8041 7147 8075
rect 7147 8041 7156 8075
rect 7104 8032 7156 8041
rect 8576 8032 8628 8084
rect 9220 8075 9272 8084
rect 9220 8041 9229 8075
rect 9229 8041 9263 8075
rect 9263 8041 9272 8075
rect 9220 8032 9272 8041
rect 10692 8032 10744 8084
rect 12808 8032 12860 8084
rect 17500 8032 17552 8084
rect 18328 8032 18380 8084
rect 19524 8032 19576 8084
rect 20168 8032 20220 8084
rect 5356 7964 5408 8016
rect 16028 7964 16080 8016
rect 5632 7896 5684 7948
rect 8116 7939 8168 7948
rect 8116 7905 8150 7939
rect 8150 7905 8168 7939
rect 10324 7939 10376 7948
rect 8116 7896 8168 7905
rect 10324 7905 10333 7939
rect 10333 7905 10367 7939
rect 10367 7905 10376 7939
rect 10324 7896 10376 7905
rect 10876 7896 10928 7948
rect 12716 7939 12768 7948
rect 12716 7905 12725 7939
rect 12725 7905 12759 7939
rect 12759 7905 12768 7939
rect 12716 7896 12768 7905
rect 16304 7896 16356 7948
rect 16672 7896 16724 7948
rect 18052 7964 18104 8016
rect 19156 7964 19208 8016
rect 17132 7939 17184 7948
rect 17132 7905 17166 7939
rect 17166 7905 17184 7939
rect 17132 7896 17184 7905
rect 2504 7760 2556 7812
rect 6920 7828 6972 7880
rect 9680 7828 9732 7880
rect 12164 7828 12216 7880
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 19892 7871 19944 7880
rect 12900 7828 12952 7837
rect 19892 7837 19901 7871
rect 19901 7837 19935 7871
rect 19935 7837 19944 7871
rect 19892 7828 19944 7837
rect 19984 7871 20036 7880
rect 19984 7837 19993 7871
rect 19993 7837 20027 7871
rect 20027 7837 20036 7871
rect 19984 7828 20036 7837
rect 3516 7692 3568 7744
rect 13912 7760 13964 7812
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 1492 7531 1544 7540
rect 1492 7497 1501 7531
rect 1501 7497 1535 7531
rect 1535 7497 1544 7531
rect 1492 7488 1544 7497
rect 3884 7531 3936 7540
rect 3884 7497 3893 7531
rect 3893 7497 3927 7531
rect 3927 7497 3936 7531
rect 3884 7488 3936 7497
rect 5632 7488 5684 7540
rect 8116 7488 8168 7540
rect 2504 7327 2556 7336
rect 2504 7293 2513 7327
rect 2513 7293 2547 7327
rect 2547 7293 2556 7327
rect 2504 7284 2556 7293
rect 3608 7284 3660 7336
rect 3976 7352 4028 7404
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 8484 7488 8536 7540
rect 17408 7488 17460 7540
rect 17960 7488 18012 7540
rect 19892 7531 19944 7540
rect 14280 7420 14332 7472
rect 18420 7420 18472 7472
rect 18880 7420 18932 7472
rect 19064 7420 19116 7472
rect 17132 7352 17184 7404
rect 18052 7352 18104 7404
rect 19892 7497 19901 7531
rect 19901 7497 19935 7531
rect 19935 7497 19944 7531
rect 19892 7488 19944 7497
rect 20352 7352 20404 7404
rect 3884 7284 3936 7336
rect 5080 7284 5132 7336
rect 6828 7284 6880 7336
rect 9036 7284 9088 7336
rect 2688 7216 2740 7268
rect 3792 7216 3844 7268
rect 7104 7216 7156 7268
rect 12072 7216 12124 7268
rect 18420 7259 18472 7268
rect 1860 7191 1912 7200
rect 1860 7157 1869 7191
rect 1869 7157 1903 7191
rect 1903 7157 1912 7191
rect 1860 7148 1912 7157
rect 4160 7148 4212 7200
rect 5356 7148 5408 7200
rect 8392 7148 8444 7200
rect 9036 7191 9088 7200
rect 9036 7157 9045 7191
rect 9045 7157 9079 7191
rect 9079 7157 9088 7191
rect 9036 7148 9088 7157
rect 11980 7148 12032 7200
rect 18420 7225 18429 7259
rect 18429 7225 18463 7259
rect 18463 7225 18472 7259
rect 18420 7216 18472 7225
rect 19800 7284 19852 7336
rect 17684 7148 17736 7200
rect 19064 7148 19116 7200
rect 20444 7148 20496 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 18052 6987 18104 6996
rect 18052 6953 18061 6987
rect 18061 6953 18095 6987
rect 18095 6953 18104 6987
rect 18052 6944 18104 6953
rect 1584 6876 1636 6928
rect 2504 6876 2556 6928
rect 3884 6876 3936 6928
rect 4804 6876 4856 6928
rect 5264 6876 5316 6928
rect 6644 6876 6696 6928
rect 2228 6808 2280 6860
rect 5540 6851 5592 6860
rect 5540 6817 5549 6851
rect 5549 6817 5583 6851
rect 5583 6817 5592 6851
rect 5540 6808 5592 6817
rect 6552 6851 6604 6860
rect 6552 6817 6561 6851
rect 6561 6817 6595 6851
rect 6595 6817 6604 6851
rect 6552 6808 6604 6817
rect 7564 6851 7616 6860
rect 7564 6817 7573 6851
rect 7573 6817 7607 6851
rect 7607 6817 7616 6851
rect 7564 6808 7616 6817
rect 11152 6808 11204 6860
rect 16672 6851 16724 6860
rect 16672 6817 16681 6851
rect 16681 6817 16715 6851
rect 16715 6817 16724 6851
rect 16672 6808 16724 6817
rect 19248 6808 19300 6860
rect 19708 6808 19760 6860
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3332 6740 3384 6749
rect 4252 6740 4304 6792
rect 5080 6740 5132 6792
rect 3240 6672 3292 6724
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6828 6783 6880 6792
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 9680 6740 9732 6792
rect 19156 6783 19208 6792
rect 19156 6749 19165 6783
rect 19165 6749 19199 6783
rect 19199 6749 19208 6783
rect 19156 6740 19208 6749
rect 20168 6740 20220 6792
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 5632 6604 5684 6656
rect 7472 6604 7524 6656
rect 17960 6604 18012 6656
rect 20628 6604 20680 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 2964 6443 3016 6452
rect 2964 6409 2973 6443
rect 2973 6409 3007 6443
rect 3007 6409 3016 6443
rect 2964 6400 3016 6409
rect 5540 6400 5592 6452
rect 19248 6400 19300 6452
rect 20352 6400 20404 6452
rect 3608 6307 3660 6316
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 5080 6264 5132 6316
rect 19156 6264 19208 6316
rect 3332 6239 3384 6248
rect 3332 6205 3341 6239
rect 3341 6205 3375 6239
rect 3375 6205 3384 6239
rect 3332 6196 3384 6205
rect 5356 6239 5408 6248
rect 5356 6205 5365 6239
rect 5365 6205 5399 6239
rect 5399 6205 5408 6239
rect 5356 6196 5408 6205
rect 4068 6128 4120 6180
rect 10048 6128 10100 6180
rect 20628 6128 20680 6180
rect 3332 6060 3384 6112
rect 3700 6060 3752 6112
rect 4160 6060 4212 6112
rect 4896 6060 4948 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 3976 5856 4028 5908
rect 8300 5856 8352 5908
rect 19800 5899 19852 5908
rect 19800 5865 19809 5899
rect 19809 5865 19843 5899
rect 19843 5865 19852 5899
rect 19800 5856 19852 5865
rect 20168 5899 20220 5908
rect 20168 5865 20177 5899
rect 20177 5865 20211 5899
rect 20211 5865 20220 5899
rect 20168 5856 20220 5865
rect 20260 5695 20312 5704
rect 20260 5661 20269 5695
rect 20269 5661 20303 5695
rect 20303 5661 20312 5695
rect 20260 5652 20312 5661
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20352 5652 20404 5661
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 5908 5312 5960 5364
rect 17960 5312 18012 5364
rect 20260 5312 20312 5364
rect 4068 5244 4120 5296
rect 11980 5244 12032 5296
rect 20628 5219 20680 5228
rect 20628 5185 20637 5219
rect 20637 5185 20671 5219
rect 20671 5185 20680 5219
rect 20628 5176 20680 5185
rect 4068 4972 4120 5024
rect 20536 5015 20588 5024
rect 20536 4981 20545 5015
rect 20545 4981 20579 5015
rect 20579 4981 20588 5015
rect 20536 4972 20588 4981
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 6368 3068 6420 3120
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 4988 3000 5040 3009
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 11152 2932 11204 2984
rect 15844 2932 15896 2984
rect 20444 2864 20496 2916
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 2780 960 2832 1012
rect 4712 960 4764 1012
<< metal2 >>
rect 202 22320 258 22800
rect 570 22320 626 22800
rect 1030 22320 1086 22800
rect 1398 22320 1454 22800
rect 1858 22320 1914 22800
rect 2226 22320 2282 22800
rect 2686 22320 2742 22800
rect 3054 22536 3110 22545
rect 3054 22471 3110 22480
rect 216 19990 244 22320
rect 204 19984 256 19990
rect 204 19926 256 19932
rect 584 15910 612 22320
rect 1044 19242 1072 22320
rect 1032 19236 1084 19242
rect 1032 19178 1084 19184
rect 1412 19145 1440 22320
rect 1398 19136 1454 19145
rect 1398 19071 1454 19080
rect 1872 19009 1900 22320
rect 2240 20074 2268 22320
rect 2240 20046 2544 20074
rect 2516 19990 2544 20046
rect 2504 19984 2556 19990
rect 2504 19926 2556 19932
rect 1950 19816 2006 19825
rect 1950 19751 2006 19760
rect 1964 19514 1992 19751
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 2136 19304 2188 19310
rect 2136 19246 2188 19252
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 1858 19000 1914 19009
rect 1858 18935 1914 18944
rect 1950 18864 2006 18873
rect 1950 18799 2006 18808
rect 1964 18426 1992 18799
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1950 18320 2006 18329
rect 1950 18255 2006 18264
rect 1964 17882 1992 18255
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 1950 17368 2006 17377
rect 1950 17303 1952 17312
rect 2004 17303 2006 17312
rect 1952 17274 2004 17280
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 572 15904 624 15910
rect 572 15846 624 15852
rect 1780 15026 1808 17070
rect 2148 16998 2176 19246
rect 2332 18057 2360 19246
rect 2410 19136 2466 19145
rect 2410 19071 2466 19080
rect 2318 18048 2374 18057
rect 2318 17983 2374 17992
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2136 16992 2188 16998
rect 1950 16960 2006 16969
rect 2136 16934 2188 16940
rect 1950 16895 2006 16904
rect 1964 16794 1992 16895
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 1950 16552 2006 16561
rect 1950 16487 2006 16496
rect 1964 16250 1992 16487
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 1950 16008 2006 16017
rect 1950 15943 2006 15952
rect 1964 15706 1992 15943
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1950 15600 2006 15609
rect 1950 15535 2006 15544
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1964 14618 1992 15535
rect 2240 15026 2268 16050
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 1766 14104 1822 14113
rect 1766 14039 1822 14048
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1504 12238 1532 12718
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1504 11286 1532 12174
rect 1492 11280 1544 11286
rect 1492 11222 1544 11228
rect 1504 11150 1532 11222
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1504 9466 1532 11086
rect 1596 9586 1624 13330
rect 1688 12986 1716 13806
rect 1780 13530 1808 14039
rect 1872 13938 1900 14418
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 2332 13297 2360 17682
rect 2424 15570 2452 19071
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 2516 18290 2544 18770
rect 2608 18329 2636 19654
rect 2594 18320 2650 18329
rect 2504 18284 2556 18290
rect 2594 18255 2650 18264
rect 2504 18226 2556 18232
rect 2504 17876 2556 17882
rect 2504 17818 2556 17824
rect 2516 17785 2544 17818
rect 2502 17776 2558 17785
rect 2502 17711 2558 17720
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2608 16794 2636 17614
rect 2700 17270 2728 22320
rect 2962 22128 3018 22137
rect 2962 22063 3018 22072
rect 2778 21584 2834 21593
rect 2778 21519 2834 21528
rect 2792 20058 2820 21519
rect 2870 20632 2926 20641
rect 2870 20567 2926 20576
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2778 19272 2834 19281
rect 2778 19207 2834 19216
rect 2792 18970 2820 19207
rect 2884 19174 2912 20567
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2976 18698 3004 22063
rect 2964 18692 3016 18698
rect 2964 18634 3016 18640
rect 3068 18426 3096 22471
rect 3146 22320 3202 22800
rect 3514 22320 3570 22800
rect 3974 22320 4030 22800
rect 4342 22320 4398 22800
rect 4802 22320 4858 22800
rect 5262 22320 5318 22800
rect 5630 22320 5686 22800
rect 6090 22320 6146 22800
rect 6458 22320 6514 22800
rect 6918 22320 6974 22800
rect 7378 22320 7434 22800
rect 7746 22320 7802 22800
rect 8206 22320 8262 22800
rect 8574 22320 8630 22800
rect 9034 22320 9090 22800
rect 9494 22320 9550 22800
rect 9862 22320 9918 22800
rect 10322 22320 10378 22800
rect 10690 22320 10746 22800
rect 11150 22320 11206 22800
rect 11610 22320 11666 22800
rect 11978 22320 12034 22800
rect 12438 22320 12494 22800
rect 12806 22320 12862 22800
rect 13266 22320 13322 22800
rect 13634 22320 13690 22800
rect 14094 22320 14150 22800
rect 14554 22320 14610 22800
rect 14922 22320 14978 22800
rect 15382 22320 15438 22800
rect 15750 22320 15806 22800
rect 16210 22320 16266 22800
rect 16670 22320 16726 22800
rect 17038 22320 17094 22800
rect 17498 22320 17554 22800
rect 17866 22320 17922 22800
rect 18326 22320 18382 22800
rect 18786 22320 18842 22800
rect 19154 22320 19210 22800
rect 19614 22320 19670 22800
rect 19982 22320 20038 22800
rect 20442 22320 20498 22800
rect 20718 22536 20774 22545
rect 20718 22471 20774 22480
rect 3160 19854 3188 22320
rect 3422 20224 3478 20233
rect 3422 20159 3478 20168
rect 3240 19984 3292 19990
rect 3240 19926 3292 19932
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3160 19281 3188 19654
rect 3146 19272 3202 19281
rect 3146 19207 3202 19216
rect 3252 18816 3280 19926
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 3160 18788 3280 18816
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 2778 17912 2834 17921
rect 2778 17847 2834 17856
rect 2792 17338 2820 17847
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2688 17264 2740 17270
rect 2688 17206 2740 17212
rect 2596 16788 2648 16794
rect 2596 16730 2648 16736
rect 2778 16144 2834 16153
rect 2778 16079 2834 16088
rect 2792 15910 2820 16079
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 2792 15706 2820 15846
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2412 14476 2464 14482
rect 2412 14418 2464 14424
rect 2424 13870 2452 14418
rect 2792 14074 2820 14991
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 2318 13288 2374 13297
rect 2318 13223 2374 13232
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1872 10810 1900 12582
rect 1964 11898 1992 12582
rect 2792 12442 2820 12718
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 1952 11892 2004 11898
rect 1952 11834 2004 11840
rect 2700 11762 2728 12242
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 2700 11354 2728 11698
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 2516 10606 2544 11154
rect 2700 10674 2728 11290
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 1872 10266 1900 10406
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 2516 10062 2544 10542
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2332 9722 2360 9998
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2884 9602 2912 14418
rect 2976 13954 3004 17682
rect 3160 17649 3188 18788
rect 3238 18728 3294 18737
rect 3238 18663 3240 18672
rect 3292 18663 3294 18672
rect 3240 18634 3292 18640
rect 3146 17640 3202 17649
rect 3146 17575 3202 17584
rect 3160 16794 3188 17575
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3068 15638 3096 16526
rect 3252 15978 3280 16526
rect 3240 15972 3292 15978
rect 3240 15914 3292 15920
rect 3056 15632 3108 15638
rect 3056 15574 3108 15580
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3252 14890 3280 15438
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 3146 14648 3202 14657
rect 3146 14583 3202 14592
rect 3160 14074 3188 14583
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 2976 13926 3096 13954
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2976 13462 3004 13806
rect 2964 13456 3016 13462
rect 2964 13398 3016 13404
rect 3068 13308 3096 13926
rect 3146 13696 3202 13705
rect 3146 13631 3202 13640
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 2792 9574 2912 9602
rect 2976 13280 3096 13308
rect 2228 9512 2280 9518
rect 1504 9450 1624 9466
rect 2228 9454 2280 9460
rect 1504 9444 1636 9450
rect 1504 9438 1584 9444
rect 1584 9386 1636 9392
rect 1596 8430 1624 9386
rect 2240 9178 2268 9454
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1492 8016 1544 8022
rect 1492 7958 1544 7964
rect 1504 7546 1532 7958
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1596 6934 1624 8366
rect 2608 8090 2636 8978
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2596 8084 2648 8090
rect 2596 8026 2648 8032
rect 2700 7886 2728 8366
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 2516 7342 2544 7754
rect 2504 7336 2556 7342
rect 2792 7324 2820 9574
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2884 8974 2912 9386
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 8634 2912 8910
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2976 8480 3004 13280
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 3068 10198 3096 10406
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 3160 9994 3188 13631
rect 3148 9988 3200 9994
rect 3148 9930 3200 9936
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3160 8634 3188 8842
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 2884 8452 3004 8480
rect 2884 7585 2912 8452
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2870 7576 2926 7585
rect 2870 7511 2926 7520
rect 2792 7296 2912 7324
rect 2504 7278 2556 7284
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1584 6928 1636 6934
rect 1584 6870 1636 6876
rect 1872 2553 1900 7142
rect 2516 6934 2544 7278
rect 2688 7268 2740 7274
rect 2740 7228 2820 7256
rect 2688 7210 2740 7216
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 1858 2544 1914 2553
rect 1858 2479 1914 2488
rect 2240 480 2268 6802
rect 2792 1601 2820 7228
rect 2884 4321 2912 7296
rect 2976 6458 3004 7890
rect 3252 6730 3280 14826
rect 3344 14498 3372 19858
rect 3436 19514 3464 20159
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3528 18358 3556 22320
rect 3698 21176 3754 21185
rect 3698 21111 3754 21120
rect 3712 21010 3740 21111
rect 3700 21004 3752 21010
rect 3700 20946 3752 20952
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3516 18352 3568 18358
rect 3516 18294 3568 18300
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3344 14470 3464 14498
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3344 9110 3372 10066
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 3344 6254 3372 6734
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 2870 4312 2926 4321
rect 2870 4247 2926 4256
rect 3344 3505 3372 6054
rect 3436 5817 3464 14470
rect 3528 14074 3556 18158
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3528 12753 3556 12854
rect 3514 12744 3570 12753
rect 3514 12679 3570 12688
rect 3514 12608 3570 12617
rect 3514 12543 3570 12552
rect 3528 11694 3556 12543
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3620 11393 3648 18770
rect 3712 18698 3740 19790
rect 3988 19310 4016 22320
rect 4160 19780 4212 19786
rect 4160 19722 4212 19728
rect 3976 19304 4028 19310
rect 4172 19258 4200 19722
rect 4356 19700 4384 22320
rect 3976 19246 4028 19252
rect 4080 19230 4200 19258
rect 4264 19672 4384 19700
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 3700 18692 3752 18698
rect 3700 18634 3752 18640
rect 3804 18290 3832 18906
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3792 18284 3844 18290
rect 3792 18226 3844 18232
rect 3792 17876 3844 17882
rect 3792 17818 3844 17824
rect 3804 17202 3832 17818
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3700 16992 3752 16998
rect 3700 16934 3752 16940
rect 3712 16697 3740 16934
rect 3698 16688 3754 16697
rect 3698 16623 3754 16632
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3712 15638 3740 15914
rect 3700 15632 3752 15638
rect 3700 15574 3752 15580
rect 3712 15094 3740 15574
rect 3700 15088 3752 15094
rect 3700 15030 3752 15036
rect 3712 14414 3740 15030
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3698 12880 3754 12889
rect 3804 12866 3832 16594
rect 3754 12838 3832 12866
rect 3698 12815 3754 12824
rect 3712 11626 3740 12815
rect 3700 11620 3752 11626
rect 3700 11562 3752 11568
rect 3792 11620 3844 11626
rect 3792 11562 3844 11568
rect 3606 11384 3662 11393
rect 3606 11319 3662 11328
rect 3804 10674 3832 11562
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3528 8090 3556 8230
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7177 3556 7686
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3514 7168 3570 7177
rect 3514 7103 3570 7112
rect 3620 6322 3648 7278
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3712 6118 3740 8910
rect 3804 7274 3832 9522
rect 3896 9489 3924 18702
rect 3988 18426 4016 18702
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3988 15706 4016 16934
rect 4080 16833 4108 19230
rect 4264 19174 4292 19672
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4172 18426 4200 19110
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4264 18873 4292 18906
rect 4250 18864 4306 18873
rect 4250 18799 4306 18808
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4816 18465 4844 22320
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4802 18456 4858 18465
rect 4160 18420 4212 18426
rect 4802 18391 4858 18400
rect 4160 18362 4212 18368
rect 4908 18290 4936 18770
rect 4896 18284 4948 18290
rect 4896 18226 4948 18232
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 4172 17338 4200 18158
rect 4816 17762 4844 18158
rect 4252 17740 4304 17746
rect 4816 17734 4936 17762
rect 4252 17682 4304 17688
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4066 16824 4122 16833
rect 4066 16759 4122 16768
rect 4160 16720 4212 16726
rect 4160 16662 4212 16668
rect 4172 16250 4200 16662
rect 4264 16250 4292 17682
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4724 16726 4752 17614
rect 4816 17338 4844 17614
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4172 14618 4200 15438
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4264 14482 4292 16050
rect 4724 15502 4752 16662
rect 4816 16658 4844 17274
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4816 16250 4844 16594
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4908 15910 4936 17734
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4908 15366 4936 15846
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4264 13870 4292 14418
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3988 12986 4016 13738
rect 4724 13462 4752 15302
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4712 13456 4764 13462
rect 4712 13398 4764 13404
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 4068 12368 4120 12374
rect 4066 12336 4068 12345
rect 4120 12336 4122 12345
rect 4066 12271 4122 12280
rect 4172 11898 4200 13330
rect 4264 12850 4292 13330
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4264 12238 4292 12378
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4066 11792 4122 11801
rect 4264 11778 4292 12174
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4066 11727 4122 11736
rect 4172 11750 4292 11778
rect 4080 11694 4108 11727
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4172 11286 4200 11750
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 3974 10840 4030 10849
rect 3974 10775 4030 10784
rect 3988 9994 4016 10775
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 4080 10266 4108 10406
rect 4172 10266 4200 11222
rect 4264 10810 4292 11494
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4724 10742 4752 13262
rect 4816 13258 4844 14758
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4816 11762 4844 12038
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 3882 9480 3938 9489
rect 3882 9415 3938 9424
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 4080 9081 4108 9386
rect 4066 9072 4122 9081
rect 4066 9007 4122 9016
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4080 8537 4108 8842
rect 4066 8528 4122 8537
rect 4066 8463 4122 8472
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3896 7546 3924 7822
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3988 7410 4016 7822
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3896 6934 3924 7278
rect 4172 7206 4200 9998
rect 4264 9382 4292 10542
rect 4356 10062 4384 10678
rect 4816 10554 4844 11154
rect 4908 10810 4936 12718
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4632 10526 4844 10554
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4632 10198 4660 10526
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4632 10062 4660 10134
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4724 9178 4752 10066
rect 4816 9518 4844 10406
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4908 9178 4936 10542
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 4710 9072 4766 9081
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 3884 6928 3936 6934
rect 3884 6870 3936 6876
rect 4264 6798 4292 9046
rect 4710 9007 4766 9016
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4724 7954 4752 9007
rect 4804 8968 4856 8974
rect 4802 8936 4804 8945
rect 4856 8936 4858 8945
rect 4802 8871 4858 8880
rect 4802 8528 4858 8537
rect 4802 8463 4804 8472
rect 4856 8463 4858 8472
rect 4804 8434 4856 8440
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4252 6792 4304 6798
rect 4066 6760 4122 6769
rect 4252 6734 4304 6740
rect 4066 6695 4122 6704
rect 3974 6216 4030 6225
rect 4080 6186 4108 6695
rect 3974 6151 4030 6160
rect 4068 6180 4120 6186
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3988 5914 4016 6151
rect 4068 6122 4120 6128
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3422 5808 3478 5817
rect 3422 5743 3478 5752
rect 4068 5296 4120 5302
rect 4066 5264 4068 5273
rect 4120 5264 4122 5273
rect 4066 5199 4122 5208
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4865 4108 4966
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 4172 3913 4200 6054
rect 4158 3904 4214 3913
rect 4158 3839 4214 3848
rect 3330 3496 3386 3505
rect 3330 3431 3386 3440
rect 4264 2009 4292 6734
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4250 2000 4306 2009
rect 4250 1935 4306 1944
rect 2778 1592 2834 1601
rect 2778 1527 2834 1536
rect 4724 1018 4752 7890
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4816 2961 4844 6870
rect 4908 6118 4936 9114
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 5000 3058 5028 19110
rect 5080 18692 5132 18698
rect 5080 18634 5132 18640
rect 5092 16454 5120 18634
rect 5276 16522 5304 22320
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5552 18601 5580 19246
rect 5538 18592 5594 18601
rect 5538 18527 5594 18536
rect 5644 18290 5672 22320
rect 6104 21162 6132 22320
rect 6104 21134 6224 21162
rect 6092 21004 6144 21010
rect 6092 20946 6144 20952
rect 6104 19514 6132 20946
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 5920 18902 5948 19246
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 6196 18154 6224 21134
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6288 18193 6316 18770
rect 6472 18290 6500 22320
rect 6644 19236 6696 19242
rect 6644 19178 6696 19184
rect 6550 18592 6606 18601
rect 6550 18527 6606 18536
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6274 18184 6330 18193
rect 6092 18148 6144 18154
rect 6092 18090 6144 18096
rect 6184 18148 6236 18154
rect 6274 18119 6330 18128
rect 6184 18090 6236 18096
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5644 17270 5672 17478
rect 5920 17338 5948 17682
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 5632 17264 5684 17270
rect 5632 17206 5684 17212
rect 5448 17060 5500 17066
rect 5448 17002 5500 17008
rect 5460 16794 5488 17002
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5264 16516 5316 16522
rect 5264 16458 5316 16464
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 5092 16046 5120 16390
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 5276 15638 5304 16050
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 5368 15434 5396 15642
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5092 14074 5120 14418
rect 5368 14074 5396 14758
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5092 13938 5120 14010
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5368 12714 5396 13398
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 5092 10010 5120 12582
rect 5264 12300 5316 12306
rect 5316 12260 5396 12288
rect 5264 12242 5316 12248
rect 5368 11762 5396 12260
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5368 11014 5396 11698
rect 5460 11354 5488 15914
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5552 15366 5580 15438
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5736 14498 5764 16458
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5828 14618 5856 14962
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5540 14476 5592 14482
rect 5736 14470 5856 14498
rect 5540 14418 5592 14424
rect 5552 13802 5580 14418
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5552 13326 5580 13738
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5552 12850 5580 13262
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11354 5580 11494
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 5184 10538 5212 10678
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5276 10470 5304 10746
rect 5368 10674 5396 10950
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5092 9982 5212 10010
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5092 9110 5120 9862
rect 5080 9104 5132 9110
rect 5184 9081 5212 9982
rect 5080 9046 5132 9052
rect 5170 9072 5226 9081
rect 5170 9007 5226 9016
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5078 8120 5134 8129
rect 5078 8055 5080 8064
rect 5132 8055 5134 8064
rect 5080 8026 5132 8032
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5092 6798 5120 7278
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5092 6322 5120 6734
rect 5184 6662 5212 8298
rect 5276 6934 5304 10406
rect 5460 9178 5488 11154
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5552 9586 5580 10202
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5356 9104 5408 9110
rect 5354 9072 5356 9081
rect 5408 9072 5410 9081
rect 5736 9042 5764 9318
rect 5354 9007 5410 9016
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 8634 5396 8774
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5552 8537 5580 8570
rect 5538 8528 5594 8537
rect 5538 8463 5594 8472
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5356 8016 5408 8022
rect 5354 7984 5356 7993
rect 5408 7984 5410 7993
rect 5354 7919 5410 7928
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 5368 6254 5396 7142
rect 5552 7018 5580 8230
rect 5644 7954 5672 8434
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5644 7546 5672 7890
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5644 7426 5672 7482
rect 5644 7398 5764 7426
rect 5552 6990 5672 7018
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5552 6458 5580 6802
rect 5644 6662 5672 6990
rect 5736 6798 5764 7398
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5828 3058 5856 14470
rect 6012 14113 6040 17750
rect 5998 14104 6054 14113
rect 5998 14039 6054 14048
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 6012 13326 6040 13874
rect 6104 13530 6132 18090
rect 6182 18048 6238 18057
rect 6182 17983 6238 17992
rect 6196 15706 6224 17983
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5920 12986 5948 13262
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 6196 12850 6224 15642
rect 6380 15473 6408 18226
rect 6366 15464 6422 15473
rect 6366 15399 6422 15408
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5920 11694 5948 12038
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 6012 11354 6040 12582
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 5920 5370 5948 11222
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6012 10130 6040 10610
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6012 9586 6040 10066
rect 6104 9722 6132 12582
rect 6288 11642 6316 13330
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6196 11614 6316 11642
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6012 8974 6040 9522
rect 6196 9042 6224 11614
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 11354 6316 11494
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6380 10674 6408 12786
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6472 10606 6500 11494
rect 6460 10600 6512 10606
rect 6366 10568 6422 10577
rect 6460 10542 6512 10548
rect 6366 10503 6422 10512
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6012 8090 6040 8230
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 6380 3126 6408 10503
rect 6472 10198 6500 10542
rect 6460 10192 6512 10198
rect 6564 10169 6592 18527
rect 6656 13462 6684 19178
rect 6826 19000 6882 19009
rect 6826 18935 6882 18944
rect 6736 18352 6788 18358
rect 6736 18294 6788 18300
rect 6748 17241 6776 18294
rect 6840 18222 6868 18935
rect 6932 18272 6960 22320
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7300 19145 7328 19246
rect 7286 19136 7342 19145
rect 7286 19071 7342 19080
rect 7288 18284 7340 18290
rect 6932 18244 7144 18272
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6840 17814 6868 18158
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6840 17338 6868 17614
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6734 17232 6790 17241
rect 6734 17167 6790 17176
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 13870 6868 14758
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6932 11082 6960 18090
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 7024 17202 7052 18022
rect 7116 17218 7144 18244
rect 7288 18226 7340 18232
rect 7012 17196 7064 17202
rect 7116 17190 7236 17218
rect 7012 17138 7064 17144
rect 7010 17096 7066 17105
rect 7010 17031 7066 17040
rect 7104 17060 7156 17066
rect 7024 11354 7052 17031
rect 7104 17002 7156 17008
rect 7116 14618 7144 17002
rect 7208 16017 7236 17190
rect 7194 16008 7250 16017
rect 7194 15943 7250 15952
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15745 7236 15846
rect 7194 15736 7250 15745
rect 7194 15671 7250 15680
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7116 11694 7144 12378
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6460 10134 6512 10140
rect 6550 10160 6606 10169
rect 6550 10095 6606 10104
rect 6564 10044 6592 10095
rect 6472 10016 6592 10044
rect 6472 8129 6500 10016
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6458 8120 6514 8129
rect 6458 8055 6514 8064
rect 6564 6866 6592 8978
rect 6656 6934 6684 9658
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 4802 2952 4858 2961
rect 4802 2887 4858 2896
rect 6564 1057 6592 6802
rect 6550 1048 6606 1057
rect 2780 1012 2832 1018
rect 2780 954 2832 960
rect 4712 1012 4764 1018
rect 6550 983 6606 992
rect 4712 954 4764 960
rect 2792 649 2820 954
rect 2778 640 2834 649
rect 2778 575 2834 584
rect 6748 480 6776 9318
rect 7208 8974 7236 15506
rect 7300 15162 7328 18226
rect 7392 17105 7420 22320
rect 7564 19780 7616 19786
rect 7564 19722 7616 19728
rect 7576 18766 7604 19722
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7668 18698 7696 19110
rect 7656 18692 7708 18698
rect 7656 18634 7708 18640
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7484 17746 7512 18226
rect 7668 17882 7696 18634
rect 7760 18465 7788 22320
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 7746 18456 7802 18465
rect 7746 18391 7802 18400
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 7472 17604 7524 17610
rect 7472 17546 7524 17552
rect 7378 17096 7434 17105
rect 7378 17031 7434 17040
rect 7484 16726 7512 17546
rect 7576 17202 7604 17818
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 7564 17196 7616 17202
rect 7564 17138 7616 17144
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7392 16590 7420 16662
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7288 13864 7340 13870
rect 7392 13852 7420 16526
rect 7484 16522 7512 16662
rect 7576 16658 7604 17138
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7472 16516 7524 16522
rect 7472 16458 7524 16464
rect 7576 16130 7604 16594
rect 7668 16250 7696 17682
rect 7760 17202 7788 18226
rect 8220 18034 8248 22320
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8312 19378 8340 19654
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8496 18601 8524 19858
rect 8588 19666 8616 22320
rect 8852 19848 8904 19854
rect 8852 19790 8904 19796
rect 8588 19638 8708 19666
rect 8680 19310 8708 19638
rect 8864 19514 8892 19790
rect 8852 19508 8904 19514
rect 8852 19450 8904 19456
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8482 18592 8538 18601
rect 8482 18527 8538 18536
rect 8574 18456 8630 18465
rect 8574 18391 8630 18400
rect 8588 18222 8616 18391
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8668 18148 8720 18154
rect 8668 18090 8720 18096
rect 8680 18057 8708 18090
rect 8666 18048 8722 18057
rect 8220 18006 8524 18034
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8312 17542 8340 17818
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8206 17232 8262 17241
rect 7748 17196 7800 17202
rect 8206 17167 8262 17176
rect 7748 17138 7800 17144
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7576 16114 7696 16130
rect 7760 16114 7788 17138
rect 8220 17134 8248 17167
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8312 16658 8340 17478
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 7576 16108 7708 16114
rect 7576 16102 7656 16108
rect 7656 16050 7708 16056
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 7562 16008 7618 16017
rect 7562 15943 7618 15952
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7340 13824 7420 13852
rect 7288 13806 7340 13812
rect 7300 13326 7328 13806
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7484 10588 7512 15438
rect 7576 14890 7604 15943
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7668 15434 7696 15846
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8114 15600 8170 15609
rect 8114 15535 8116 15544
rect 8168 15535 8170 15544
rect 8116 15506 8168 15512
rect 8220 15502 8248 16050
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8312 15638 8340 15846
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 7656 15428 7708 15434
rect 7656 15370 7708 15376
rect 7840 15428 7892 15434
rect 7840 15370 7892 15376
rect 7852 15162 7880 15370
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7576 14550 7604 14826
rect 7668 14822 7696 15098
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7760 14414 7788 14962
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7576 13870 7604 14214
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7576 13394 7604 13806
rect 7760 13734 7788 14214
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7668 12850 7696 13126
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 8220 12442 8248 14894
rect 8312 14618 8340 14894
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7760 11694 7788 12174
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 8116 11688 8168 11694
rect 8168 11636 8340 11642
rect 8116 11630 8340 11636
rect 8128 11614 8340 11630
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7300 10560 7512 10588
rect 7300 10146 7328 10560
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7484 10266 7512 10406
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7300 10118 7512 10146
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7392 9110 7420 9454
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7196 8968 7248 8974
rect 7300 8945 7328 8978
rect 7196 8910 7248 8916
rect 7286 8936 7342 8945
rect 7286 8871 7342 8880
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6840 7342 6868 8298
rect 7116 8090 7144 8434
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6932 7410 6960 7822
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6840 6798 6868 7278
rect 7116 7274 7144 8026
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 7484 6662 7512 10118
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 9364 7604 10066
rect 7668 9518 7696 10610
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7576 9336 7696 9364
rect 7668 8974 7696 9336
rect 7760 9178 7788 10406
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8220 9178 8248 11154
rect 8312 10470 8340 11614
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8404 9518 8432 15846
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8404 9058 8432 9454
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 8312 9030 8432 9058
rect 7656 8968 7708 8974
rect 7944 8945 7972 8978
rect 7656 8910 7708 8916
rect 7930 8936 7986 8945
rect 7930 8871 7986 8880
rect 7944 8362 7972 8871
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8128 7546 8156 7890
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 2226 0 2282 480
rect 6734 0 6790 480
rect 7576 241 7604 6802
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8312 5914 8340 9030
rect 8496 8480 8524 18006
rect 8666 17983 8722 17992
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8588 16046 8616 17682
rect 8666 17368 8722 17377
rect 8666 17303 8722 17312
rect 8680 17066 8708 17303
rect 8772 17066 8800 18906
rect 8864 18834 8892 19450
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8864 18290 8892 18770
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8956 18222 8984 19110
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 8864 17134 8892 17546
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8668 17060 8720 17066
rect 8668 17002 8720 17008
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 8956 16998 8984 17682
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8588 15434 8616 15982
rect 8576 15428 8628 15434
rect 8576 15370 8628 15376
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8864 14414 8892 14758
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8680 13462 8708 14010
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8668 13456 8720 13462
rect 8668 13398 8720 13404
rect 8680 12850 8708 13398
rect 8864 13258 8892 13738
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8772 12442 8800 12582
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8772 11354 8800 12174
rect 8864 11694 8892 13194
rect 8956 12850 8984 13806
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8956 11558 8984 12038
rect 9048 11694 9076 22320
rect 9508 19802 9536 22320
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 9140 19774 9536 19802
rect 9140 14890 9168 19774
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9404 19440 9456 19446
rect 9404 19382 9456 19388
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9232 18426 9260 19110
rect 9324 18465 9352 19110
rect 9416 18970 9444 19382
rect 9404 18964 9456 18970
rect 9404 18906 9456 18912
rect 9416 18834 9444 18906
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9310 18456 9366 18465
rect 9220 18420 9272 18426
rect 9310 18391 9366 18400
rect 9220 18362 9272 18368
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9232 17814 9260 18022
rect 9508 17882 9536 19654
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9220 17808 9272 17814
rect 9312 17808 9364 17814
rect 9220 17750 9272 17756
rect 9310 17776 9312 17785
rect 9364 17776 9366 17785
rect 9310 17711 9366 17720
rect 9600 17649 9628 19858
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9692 18222 9720 18702
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9692 17678 9720 18158
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9784 17882 9812 18090
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9784 17746 9812 17818
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9680 17672 9732 17678
rect 9586 17640 9642 17649
rect 9680 17614 9732 17620
rect 9586 17575 9642 17584
rect 9586 17368 9642 17377
rect 9586 17303 9588 17312
rect 9640 17303 9642 17312
rect 9588 17274 9640 17280
rect 9496 17264 9548 17270
rect 9496 17206 9548 17212
rect 9220 17060 9272 17066
rect 9220 17002 9272 17008
rect 9232 16153 9260 17002
rect 9508 16998 9536 17206
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9586 16824 9642 16833
rect 9586 16759 9642 16768
rect 9600 16522 9628 16759
rect 9692 16658 9720 17614
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9876 16946 9904 22320
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 9968 19514 9996 19790
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 9968 17066 9996 19450
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9218 16144 9274 16153
rect 9218 16079 9274 16088
rect 9692 16046 9720 16390
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9784 15978 9812 16934
rect 9876 16918 9996 16946
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9876 16046 9904 16594
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9876 15586 9904 15982
rect 9784 15570 9904 15586
rect 9772 15564 9904 15570
rect 9824 15558 9904 15564
rect 9772 15506 9824 15512
rect 9678 15464 9734 15473
rect 9678 15399 9734 15408
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 9140 14550 9168 14826
rect 9692 14770 9720 15399
rect 9968 15162 9996 16918
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9600 14742 9720 14770
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 9600 14498 9628 14742
rect 9678 14648 9734 14657
rect 9784 14618 9812 14758
rect 9678 14583 9680 14592
rect 9732 14583 9734 14592
rect 9772 14612 9824 14618
rect 9680 14554 9732 14560
rect 9772 14554 9824 14560
rect 9600 14470 9720 14498
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9600 13802 9628 13874
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9140 11642 9168 13262
rect 9232 12986 9260 13670
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9310 13424 9366 13433
rect 9310 13359 9366 13368
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9232 11830 9260 12242
rect 9220 11824 9272 11830
rect 9220 11766 9272 11772
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 9048 11354 9076 11630
rect 9140 11614 9260 11642
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9140 11150 9168 11494
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8588 10674 8616 10950
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8576 10464 8628 10470
rect 8680 10452 8708 10950
rect 9140 10792 9168 11086
rect 9232 11014 9260 11614
rect 9324 11082 9352 13359
rect 9416 12850 9444 13466
rect 9692 12986 9720 14470
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9784 14385 9812 14418
rect 9770 14376 9826 14385
rect 9770 14311 9826 14320
rect 9770 14240 9826 14249
rect 9770 14175 9826 14184
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9140 10764 9444 10792
rect 8944 10532 8996 10538
rect 8944 10474 8996 10480
rect 8628 10424 8708 10452
rect 8576 10406 8628 10412
rect 8588 9926 8616 10406
rect 8666 10024 8722 10033
rect 8666 9959 8722 9968
rect 8680 9926 8708 9959
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8588 9722 8616 9862
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8588 9586 8616 9658
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8404 8452 8524 8480
rect 8404 7206 8432 8452
rect 8588 8430 8616 9522
rect 8956 9110 8984 10474
rect 9140 10130 9168 10764
rect 9416 10674 9444 10764
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9324 10266 9352 10610
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 9048 8974 9076 9998
rect 9508 9042 9536 11018
rect 9600 10266 9628 11222
rect 9784 10606 9812 14175
rect 9876 13530 9904 14962
rect 9968 14482 9996 15098
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 10060 13546 10088 19246
rect 10232 18216 10284 18222
rect 10232 18158 10284 18164
rect 10244 16658 10272 18158
rect 10336 17377 10364 22320
rect 10416 19916 10468 19922
rect 10416 19858 10468 19864
rect 10322 17368 10378 17377
rect 10322 17303 10378 17312
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10336 16794 10364 17138
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10336 16590 10364 16730
rect 10324 16584 10376 16590
rect 10428 16572 10456 19858
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10520 17746 10548 19790
rect 10600 18148 10652 18154
rect 10600 18090 10652 18096
rect 10508 17740 10560 17746
rect 10508 17682 10560 17688
rect 10612 17626 10640 18090
rect 10520 17598 10640 17626
rect 10520 16726 10548 17598
rect 10598 17368 10654 17377
rect 10598 17303 10654 17312
rect 10508 16720 10560 16726
rect 10508 16662 10560 16668
rect 10428 16544 10548 16572
rect 10324 16526 10376 16532
rect 10336 15570 10364 16526
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10336 15026 10364 15506
rect 10428 15473 10456 15642
rect 10414 15464 10470 15473
rect 10414 15399 10470 15408
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 10152 13938 10180 14486
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10244 13938 10272 14350
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10336 13870 10364 14962
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10324 13864 10376 13870
rect 10138 13832 10194 13841
rect 10324 13806 10376 13812
rect 10138 13767 10194 13776
rect 10152 13734 10180 13767
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 9864 13524 9916 13530
rect 10060 13518 10272 13546
rect 9864 13466 9916 13472
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10152 12714 10180 13330
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 11286 10088 11494
rect 10152 11393 10180 12242
rect 10138 11384 10194 11393
rect 10138 11319 10194 11328
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9864 11144 9916 11150
rect 10152 11132 10180 11319
rect 9864 11086 9916 11092
rect 10060 11104 10180 11132
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9036 8968 9088 8974
rect 9128 8968 9180 8974
rect 9036 8910 9088 8916
rect 9126 8936 9128 8945
rect 9180 8936 9182 8945
rect 9126 8871 9182 8880
rect 9600 8498 9628 9454
rect 9876 9178 9904 11086
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9864 9172 9916 9178
rect 9864 9114 9916 9120
rect 9968 9042 9996 9318
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8496 7546 8524 8298
rect 8588 8090 8616 8366
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 8090 9260 8230
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9692 7886 9720 8298
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 7206 9076 7278
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9692 6798 9720 7822
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 10060 6186 10088 11104
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10152 9178 10180 10746
rect 10244 9602 10272 13518
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10336 11150 10364 12378
rect 10428 12306 10456 14758
rect 10520 14521 10548 16544
rect 10506 14512 10562 14521
rect 10506 14447 10562 14456
rect 10508 14408 10560 14414
rect 10506 14376 10508 14385
rect 10560 14376 10562 14385
rect 10506 14311 10562 14320
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 11218 10456 11494
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10322 10704 10378 10713
rect 10322 10639 10378 10648
rect 10336 10130 10364 10639
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10244 9574 10364 9602
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10336 9042 10364 9574
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10152 6225 10180 8910
rect 10336 7954 10364 8978
rect 10520 8906 10548 13670
rect 10612 12306 10640 17303
rect 10704 12442 10732 22320
rect 11164 20058 11192 22320
rect 11624 20058 11652 22320
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11612 19916 11664 19922
rect 11612 19858 11664 19864
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 10966 19000 11022 19009
rect 10966 18935 11022 18944
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10796 18222 10824 18566
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 10876 18080 10928 18086
rect 10782 18048 10838 18057
rect 10876 18022 10928 18028
rect 10980 18034 11008 18935
rect 11072 18834 11100 19654
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10782 17983 10838 17992
rect 10796 13734 10824 17983
rect 10888 17202 10916 18022
rect 10980 18006 11100 18034
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 10980 17241 11008 17682
rect 11072 17338 11100 18006
rect 11164 17882 11192 19858
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11244 18284 11296 18290
rect 11244 18226 11296 18232
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11256 17524 11284 18226
rect 11164 17496 11284 17524
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 10966 17232 11022 17241
rect 10876 17196 10928 17202
rect 10966 17167 11022 17176
rect 10876 17138 10928 17144
rect 10888 16794 10916 17138
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 11164 16402 11192 17496
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11624 17338 11652 19858
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11704 19236 11756 19242
rect 11704 19178 11756 19184
rect 11716 18358 11744 19178
rect 11808 19174 11836 19790
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11716 17746 11744 18294
rect 11992 18290 12020 22320
rect 12452 20210 12480 22320
rect 12820 20346 12848 22320
rect 12820 20318 13032 20346
rect 12452 20182 12940 20210
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 12070 18184 12126 18193
rect 12070 18119 12072 18128
rect 12124 18119 12126 18128
rect 12072 18090 12124 18096
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11808 17882 11836 18022
rect 11796 17876 11848 17882
rect 11796 17818 11848 17824
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 11808 17542 11836 17614
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11900 17202 11928 17614
rect 12084 17542 12112 17614
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 12084 17218 12112 17478
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11992 17190 12112 17218
rect 11520 16992 11572 16998
rect 11518 16960 11520 16969
rect 11888 16992 11940 16998
rect 11572 16960 11574 16969
rect 11888 16934 11940 16940
rect 11518 16895 11574 16904
rect 11900 16833 11928 16934
rect 11886 16824 11942 16833
rect 11886 16759 11942 16768
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11072 16374 11192 16402
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10888 15706 10916 15982
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10888 15026 10916 15642
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10888 14074 10916 14758
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10980 13938 11008 14214
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10612 11014 10640 11698
rect 10704 11694 10732 12174
rect 10796 11762 10824 12242
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10782 11656 10838 11665
rect 10782 11591 10838 11600
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10690 10976 10746 10985
rect 10690 10911 10746 10920
rect 10704 9722 10732 10911
rect 10796 10606 10824 11591
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10888 9110 10916 12922
rect 11072 11665 11100 16374
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11256 15638 11284 15846
rect 11244 15632 11296 15638
rect 11244 15574 11296 15580
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11624 14958 11652 15302
rect 11716 15162 11744 15506
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11348 13297 11376 13330
rect 11334 13288 11390 13297
rect 11334 13223 11390 13232
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11058 11656 11114 11665
rect 11058 11591 11114 11600
rect 11164 11370 11192 12174
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11624 11880 11652 14894
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11440 11852 11652 11880
rect 11334 11656 11390 11665
rect 11334 11591 11390 11600
rect 11348 11558 11376 11591
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11072 11342 11284 11370
rect 10966 11112 11022 11121
rect 10966 11047 11022 11056
rect 10980 10606 11008 11047
rect 11072 10810 11100 11342
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 11072 10130 11100 10746
rect 11164 10538 11192 11222
rect 11256 11082 11284 11342
rect 11440 11121 11468 11852
rect 11716 11812 11744 14214
rect 11808 13734 11836 16186
rect 11900 15910 11928 16594
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11900 15502 11928 15846
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11532 11784 11744 11812
rect 11426 11112 11482 11121
rect 11244 11076 11296 11082
rect 11426 11047 11482 11056
rect 11244 11018 11296 11024
rect 11532 10996 11560 11784
rect 11808 11744 11836 13670
rect 11992 12073 12020 17190
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11978 12064 12034 12073
rect 11978 11999 12034 12008
rect 12084 11880 12112 16934
rect 11716 11716 11836 11744
rect 11900 11852 12112 11880
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11624 11257 11652 11562
rect 11610 11248 11666 11257
rect 11610 11183 11666 11192
rect 11624 11150 11652 11183
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11532 10968 11652 10996
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11242 10568 11298 10577
rect 11152 10532 11204 10538
rect 11242 10503 11298 10512
rect 11152 10474 11204 10480
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10704 8090 10732 8230
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10888 7954 10916 9046
rect 10980 8362 11008 9318
rect 11072 8906 11100 10066
rect 11150 10024 11206 10033
rect 11256 9994 11284 10503
rect 11518 10296 11574 10305
rect 11624 10282 11652 10968
rect 11716 10713 11744 11716
rect 11794 11520 11850 11529
rect 11794 11455 11850 11464
rect 11702 10704 11758 10713
rect 11702 10639 11758 10648
rect 11808 10577 11836 11455
rect 11794 10568 11850 10577
rect 11794 10503 11850 10512
rect 11624 10254 11744 10282
rect 11518 10231 11574 10240
rect 11532 10130 11560 10231
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11150 9959 11206 9968
rect 11244 9988 11296 9994
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 11164 6866 11192 9959
rect 11244 9930 11296 9936
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11624 9518 11652 9862
rect 11612 9512 11664 9518
rect 11518 9480 11574 9489
rect 11612 9454 11664 9460
rect 11518 9415 11520 9424
rect 11572 9415 11574 9424
rect 11520 9386 11572 9392
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11612 8288 11664 8294
rect 11716 8276 11744 10254
rect 11900 10033 11928 11852
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11992 11082 12020 11698
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11978 10976 12034 10985
rect 11978 10911 12034 10920
rect 11886 10024 11942 10033
rect 11886 9959 11942 9968
rect 11794 9752 11850 9761
rect 11794 9687 11796 9696
rect 11848 9687 11850 9696
rect 11796 9658 11848 9664
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11808 8838 11836 9386
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11664 8248 11744 8276
rect 11612 8230 11664 8236
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 10138 6216 10194 6225
rect 10048 6180 10100 6186
rect 10138 6151 10194 6160
rect 10048 6122 10100 6128
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11624 5273 11652 8230
rect 11992 7206 12020 10911
rect 12084 7274 12112 11630
rect 12176 8566 12204 19994
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12452 19360 12480 19926
rect 12360 19332 12480 19360
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12268 16726 12296 18294
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 12268 15910 12296 16662
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12268 14414 12296 15846
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12268 13938 12296 14350
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 12268 13190 12296 13874
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12254 13016 12310 13025
rect 12254 12951 12310 12960
rect 12268 12850 12296 12951
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12360 12424 12388 19332
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12452 18630 12480 19110
rect 12622 19000 12678 19009
rect 12622 18935 12678 18944
rect 12636 18766 12664 18935
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12544 18222 12572 18566
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12636 17814 12664 18702
rect 12532 17808 12584 17814
rect 12530 17776 12532 17785
rect 12624 17808 12676 17814
rect 12584 17776 12586 17785
rect 12624 17750 12676 17756
rect 12530 17711 12586 17720
rect 12624 17672 12676 17678
rect 12622 17640 12624 17649
rect 12676 17640 12678 17649
rect 12622 17575 12678 17584
rect 12728 17354 12756 19994
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12820 18766 12848 19178
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12820 18290 12848 18702
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12268 12396 12388 12424
rect 12452 17326 12756 17354
rect 12268 11694 12296 12396
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12360 12073 12388 12242
rect 12452 12209 12480 17326
rect 12532 17264 12584 17270
rect 12530 17232 12532 17241
rect 12820 17252 12848 17818
rect 12584 17232 12586 17241
rect 12530 17167 12586 17176
rect 12728 17224 12848 17252
rect 12728 17105 12756 17224
rect 12714 17096 12770 17105
rect 12912 17082 12940 20182
rect 12714 17031 12770 17040
rect 12820 17054 12940 17082
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12544 15910 12572 15982
rect 12728 15978 12756 16390
rect 12716 15972 12768 15978
rect 12716 15914 12768 15920
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12820 15706 12848 17054
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 16726 12940 16934
rect 12900 16720 12952 16726
rect 12900 16662 12952 16668
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12820 15586 12848 15642
rect 13004 15586 13032 20318
rect 13280 20058 13308 22320
rect 13268 20052 13320 20058
rect 13268 19994 13320 20000
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 12728 15558 12848 15586
rect 12912 15558 13032 15586
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 12544 14618 12572 14826
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12636 14618 12664 14758
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12728 14550 12756 15558
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12820 15162 12848 15438
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12912 15026 12940 15558
rect 12992 15496 13044 15502
rect 13096 15473 13124 18838
rect 13188 18766 13216 19246
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13188 18358 13216 18702
rect 13280 18426 13308 19858
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13372 18970 13400 19790
rect 13556 19174 13584 19790
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13556 18902 13584 19110
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13268 18420 13320 18426
rect 13268 18362 13320 18368
rect 13176 18352 13228 18358
rect 13176 18294 13228 18300
rect 13544 18216 13596 18222
rect 13450 18184 13506 18193
rect 13544 18158 13596 18164
rect 13450 18119 13452 18128
rect 13504 18119 13506 18128
rect 13452 18090 13504 18096
rect 13556 18057 13584 18158
rect 13542 18048 13598 18057
rect 13542 17983 13598 17992
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13188 16998 13216 17478
rect 13176 16992 13228 16998
rect 13176 16934 13228 16940
rect 13280 15502 13308 17682
rect 13358 17640 13414 17649
rect 13358 17575 13414 17584
rect 13372 17542 13400 17575
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13648 17354 13676 22320
rect 14108 19802 14136 22320
rect 14372 20324 14424 20330
rect 14372 20266 14424 20272
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 13924 19774 14136 19802
rect 13924 18630 13952 19774
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14108 19310 14136 19654
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13464 17326 13676 17354
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13372 16522 13400 17138
rect 13360 16516 13412 16522
rect 13360 16458 13412 16464
rect 13268 15496 13320 15502
rect 12992 15438 13044 15444
rect 13082 15464 13138 15473
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 13004 14906 13032 15438
rect 13268 15438 13320 15444
rect 13082 15399 13138 15408
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 12912 14878 13032 14906
rect 12716 14544 12768 14550
rect 12716 14486 12768 14492
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12544 13326 12572 14418
rect 12912 13734 12940 14878
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12438 12200 12494 12209
rect 12438 12135 12494 12144
rect 12346 12064 12402 12073
rect 12346 11999 12402 12008
rect 12452 11898 12480 12135
rect 12544 11898 12572 12378
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12360 10810 12388 11086
rect 12622 10976 12678 10985
rect 12622 10911 12678 10920
rect 12348 10804 12400 10810
rect 12400 10764 12480 10792
rect 12348 10746 12400 10752
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12268 9994 12296 10542
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 12360 9926 12388 10542
rect 12452 10305 12480 10764
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12544 10470 12572 10678
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12438 10296 12494 10305
rect 12438 10231 12494 10240
rect 12636 10198 12664 10911
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12728 9654 12756 13330
rect 12912 13258 12940 13670
rect 13004 13530 13032 14758
rect 13082 14512 13138 14521
rect 13082 14447 13138 14456
rect 13096 14074 13124 14447
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13188 13530 13216 14962
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 13188 12753 13216 12854
rect 13174 12744 13230 12753
rect 13174 12679 13230 12688
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12912 11762 12940 12174
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 13464 11234 13492 17326
rect 13544 16992 13596 16998
rect 13542 16960 13544 16969
rect 13596 16960 13598 16969
rect 13542 16895 13598 16904
rect 13740 16522 13768 17614
rect 13820 17196 13872 17202
rect 14004 17196 14056 17202
rect 13820 17138 13872 17144
rect 13924 17156 14004 17184
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13832 16250 13860 17138
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13648 14278 13676 14962
rect 13740 14890 13768 15846
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13740 14346 13768 14826
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13648 13870 13676 14214
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 12850 13768 13126
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13648 12442 13676 12718
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13648 11694 13676 12378
rect 13832 12345 13860 14894
rect 13924 14600 13952 17156
rect 14004 17138 14056 17144
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 14108 15706 14136 16594
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 13924 14572 14136 14600
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13924 12646 13952 13126
rect 14016 12986 14044 14418
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13818 12336 13874 12345
rect 13818 12271 13874 12280
rect 13832 11744 13860 12271
rect 13832 11716 13952 11744
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13740 11354 13768 11630
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13464 11206 13768 11234
rect 13740 11150 13768 11206
rect 13832 11150 13860 11562
rect 12808 11144 12860 11150
rect 12806 11112 12808 11121
rect 13728 11144 13780 11150
rect 12860 11112 12862 11121
rect 13542 11112 13598 11121
rect 12806 11047 12862 11056
rect 12900 11076 12952 11082
rect 13728 11086 13780 11092
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13542 11047 13598 11056
rect 12900 11018 12952 11024
rect 12912 10674 12940 11018
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 12820 10266 12848 10406
rect 13372 10266 13400 10406
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12176 7886 12204 8502
rect 12268 8498 12296 8774
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12452 8537 12480 8570
rect 12438 8528 12494 8537
rect 12256 8492 12308 8498
rect 12438 8463 12494 8472
rect 12256 8434 12308 8440
rect 12544 8430 12572 9318
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12728 7954 12756 9590
rect 13280 9586 13308 10066
rect 13556 10062 13584 11047
rect 13740 10198 13768 11086
rect 13832 10674 13860 11086
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12820 8090 12848 9318
rect 12912 9178 12940 9318
rect 13096 9178 13124 9522
rect 13648 9518 13676 10066
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 12912 8294 12940 8978
rect 13450 8528 13506 8537
rect 13450 8463 13452 8472
rect 13504 8463 13506 8472
rect 13452 8434 13504 8440
rect 13648 8362 13676 8978
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12912 7886 12940 8230
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 13924 7818 13952 11716
rect 14016 11218 14044 12922
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 14108 10606 14136 14572
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14108 9489 14136 10542
rect 14200 10010 14228 19858
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14292 17921 14320 18634
rect 14278 17912 14334 17921
rect 14278 17847 14334 17856
rect 14384 17746 14412 20266
rect 14568 19242 14596 22320
rect 14936 20330 14964 22320
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 14752 19378 14780 19858
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 14556 19236 14608 19242
rect 14556 19178 14608 19184
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14568 18154 14596 18566
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14554 17776 14610 17785
rect 14372 17740 14424 17746
rect 15028 17746 15056 19858
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15212 17882 15240 19110
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15304 18766 15332 18906
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 14554 17711 14610 17720
rect 15016 17740 15068 17746
rect 14372 17682 14424 17688
rect 14568 17610 14596 17711
rect 15016 17682 15068 17688
rect 14556 17604 14608 17610
rect 14556 17546 14608 17552
rect 14370 17232 14426 17241
rect 14370 17167 14372 17176
rect 14424 17167 14426 17176
rect 15016 17196 15068 17202
rect 14372 17138 14424 17144
rect 15016 17138 15068 17144
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14660 16980 14688 17070
rect 14568 16952 14688 16980
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14278 16688 14334 16697
rect 14384 16674 14412 16730
rect 14568 16674 14596 16952
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 15028 16794 15056 17138
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 14384 16646 14596 16674
rect 15120 16658 15148 17002
rect 15304 16658 15332 18702
rect 15396 17338 15424 22320
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15488 18902 15516 19314
rect 15568 19236 15620 19242
rect 15568 19178 15620 19184
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15488 18426 15516 18838
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15580 18193 15608 19178
rect 15566 18184 15622 18193
rect 15566 18119 15622 18128
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15764 17270 15792 22320
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15948 18426 15976 19110
rect 16040 18834 16068 19858
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15856 17678 15884 18090
rect 16224 17882 16252 22320
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16592 19310 16620 19790
rect 16684 19786 16712 22320
rect 17052 20058 17080 22320
rect 17512 20058 17540 22320
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17880 19990 17908 22320
rect 18340 20058 18368 22320
rect 18800 20058 18828 22320
rect 19168 22250 19196 22320
rect 18892 22222 19196 22250
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 17868 19984 17920 19990
rect 17868 19926 17920 19932
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16776 18358 16804 19858
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17408 19168 17460 19174
rect 17408 19110 17460 19116
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 17328 18426 17356 19110
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 15750 17096 15806 17105
rect 15750 17031 15806 17040
rect 15108 16652 15160 16658
rect 14278 16623 14334 16632
rect 14292 15162 14320 16623
rect 15108 16594 15160 16600
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14476 15570 14504 15982
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 15162 14596 15438
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14752 15026 14780 15098
rect 15212 15026 15240 16458
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15304 15706 15332 16390
rect 15580 16250 15608 16526
rect 15568 16244 15620 16250
rect 15568 16186 15620 16192
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15488 15434 15516 15914
rect 15672 15586 15700 16526
rect 15580 15558 15700 15586
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15580 15162 15608 15558
rect 15764 15450 15792 17031
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 15936 16584 15988 16590
rect 15856 16544 15936 16572
rect 15856 16046 15884 16544
rect 15936 16526 15988 16532
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15672 15422 15792 15450
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 14556 14340 14608 14346
rect 14556 14282 14608 14288
rect 14568 14006 14596 14282
rect 15028 14074 15056 14418
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15120 14074 15148 14214
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 14556 14000 14608 14006
rect 14556 13942 14608 13948
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14292 11898 14320 13126
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14384 11778 14412 13738
rect 14568 13512 14596 13942
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 15028 13512 15056 13738
rect 15200 13728 15252 13734
rect 15198 13696 15200 13705
rect 15292 13728 15344 13734
rect 15252 13696 15254 13705
rect 15292 13670 15344 13676
rect 15198 13631 15254 13640
rect 15304 13530 15332 13670
rect 14568 13484 14872 13512
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14476 12306 14504 13262
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14476 12170 14504 12242
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14568 12102 14596 13262
rect 14844 12782 14872 13484
rect 14936 13484 15056 13512
rect 15292 13524 15344 13530
rect 14936 13190 14964 13484
rect 15292 13466 15344 13472
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 15028 12442 15056 13330
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14292 11750 14412 11778
rect 15028 11762 15056 12106
rect 15016 11756 15068 11762
rect 14292 11098 14320 11750
rect 15016 11698 15068 11704
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14384 11286 14412 11494
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14556 11144 14608 11150
rect 14292 11070 14412 11098
rect 14556 11086 14608 11092
rect 14200 9982 14320 10010
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14200 9722 14228 9862
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14094 9480 14150 9489
rect 14094 9415 14150 9424
rect 13912 7812 13964 7818
rect 13912 7754 13964 7760
rect 14292 7478 14320 9982
rect 14384 7857 14412 11070
rect 14568 10470 14596 11086
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14752 10810 14780 10950
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14844 10606 14872 11018
rect 15028 10810 15056 11562
rect 15120 11354 15148 12650
rect 15212 12442 15240 13398
rect 15488 12889 15516 14758
rect 15672 14618 15700 15422
rect 15856 15026 15884 15982
rect 15934 15600 15990 15609
rect 16040 15570 16068 16662
rect 16316 16561 16344 18022
rect 16500 16998 16528 18022
rect 17420 17882 17448 19110
rect 17500 18896 17552 18902
rect 17500 18838 17552 18844
rect 17512 18290 17540 18838
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17408 17876 17460 17882
rect 17408 17818 17460 17824
rect 17314 17776 17370 17785
rect 17132 17740 17184 17746
rect 17314 17711 17370 17720
rect 17132 17682 17184 17688
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16302 16552 16358 16561
rect 16302 16487 16358 16496
rect 16316 16153 16344 16487
rect 16302 16144 16358 16153
rect 16302 16079 16358 16088
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 15934 15535 15990 15544
rect 16028 15564 16080 15570
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15856 14822 15884 14962
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15948 13802 15976 15535
rect 16028 15506 16080 15512
rect 16224 14929 16252 15574
rect 16408 15502 16436 15846
rect 16500 15570 16528 16934
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16210 14920 16266 14929
rect 16210 14855 16266 14864
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16132 14385 16160 14758
rect 16118 14376 16174 14385
rect 16118 14311 16174 14320
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 16026 13560 16082 13569
rect 15752 13524 15804 13530
rect 16026 13495 16028 13504
rect 15752 13466 15804 13472
rect 16080 13495 16082 13504
rect 16028 13466 16080 13472
rect 15474 12880 15530 12889
rect 15384 12844 15436 12850
rect 15474 12815 15530 12824
rect 15384 12786 15436 12792
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15396 12170 15424 12786
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15396 12073 15424 12106
rect 15382 12064 15438 12073
rect 15382 11999 15438 12008
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15304 11150 15332 11494
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14568 9625 14596 10406
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 15028 10130 15056 10542
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 15120 10062 15148 10746
rect 15212 10282 15240 10950
rect 15396 10674 15424 11999
rect 15488 11529 15516 12815
rect 15764 12374 15792 13466
rect 16132 13326 16160 14311
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15752 12232 15804 12238
rect 15750 12200 15752 12209
rect 15804 12200 15806 12209
rect 15750 12135 15806 12144
rect 15474 11520 15530 11529
rect 15474 11455 15530 11464
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15580 10470 15608 10610
rect 15856 10606 15884 12854
rect 16132 12782 16160 13262
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 15936 12640 15988 12646
rect 16224 12617 16252 14855
rect 16316 14770 16344 15302
rect 16408 14890 16436 15438
rect 16396 14884 16448 14890
rect 16396 14826 16448 14832
rect 16316 14742 16436 14770
rect 16408 14618 16436 14742
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16304 14544 16356 14550
rect 16304 14486 16356 14492
rect 16316 13870 16344 14486
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 15936 12582 15988 12588
rect 16210 12608 16266 12617
rect 15948 11694 15976 12582
rect 16210 12543 16266 12552
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 16132 11626 16160 12174
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16316 11132 16344 13670
rect 16408 13530 16436 13874
rect 16500 13734 16528 14418
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16592 13569 16620 17274
rect 17144 17202 17172 17682
rect 17328 17678 17356 17711
rect 17512 17678 17540 18226
rect 17604 18222 17632 19110
rect 17592 18216 17644 18222
rect 17592 18158 17644 18164
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16868 16114 16896 17070
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16672 15496 16724 15502
rect 17328 15450 17356 17614
rect 17604 17338 17632 18022
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17696 15586 17724 17682
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17788 16726 17816 17138
rect 17880 17066 17908 17682
rect 17972 17542 18000 19790
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18524 19378 18552 19858
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18616 19378 18644 19654
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18248 18970 18276 19314
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18892 18426 18920 22222
rect 18970 22128 19026 22137
rect 18970 22063 19026 22072
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18880 18080 18932 18086
rect 18878 18048 18880 18057
rect 18932 18048 18934 18057
rect 18878 17983 18934 17992
rect 18602 17912 18658 17921
rect 18602 17847 18604 17856
rect 18656 17847 18658 17856
rect 18604 17818 18656 17824
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18050 17232 18106 17241
rect 18050 17167 18106 17176
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 18064 16794 18092 17167
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 17776 16720 17828 16726
rect 17776 16662 17828 16668
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18616 16114 18644 16390
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 18064 15706 18092 15982
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 17512 15570 17724 15586
rect 18708 15586 18736 17682
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18892 17252 18920 17614
rect 18984 17354 19012 22063
rect 19154 21176 19210 21185
rect 19154 21111 19210 21120
rect 19062 19816 19118 19825
rect 19062 19751 19064 19760
rect 19116 19751 19118 19760
rect 19064 19722 19116 19728
rect 19168 19174 19196 21111
rect 19628 20346 19656 22320
rect 19628 20318 19748 20346
rect 19614 20224 19670 20233
rect 19614 20159 19670 20168
rect 19628 20058 19656 20159
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 19168 17814 19196 18226
rect 19156 17808 19208 17814
rect 19156 17750 19208 17756
rect 18984 17326 19196 17354
rect 19260 17338 19288 19246
rect 19352 19242 19380 19790
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19444 18630 19472 19858
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19524 19236 19576 19242
rect 19524 19178 19576 19184
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19352 17649 19380 18294
rect 19536 18222 19564 19178
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 19432 18080 19484 18086
rect 19628 18034 19656 19790
rect 19432 18022 19484 18028
rect 19338 17640 19394 17649
rect 19338 17575 19394 17584
rect 19338 17504 19394 17513
rect 19338 17439 19394 17448
rect 19168 17270 19196 17326
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19156 17264 19208 17270
rect 18892 17224 19012 17252
rect 18788 17060 18840 17066
rect 18788 17002 18840 17008
rect 18800 15706 18828 17002
rect 18878 16552 18934 16561
rect 18878 16487 18934 16496
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 17500 15564 17724 15570
rect 17552 15558 17724 15564
rect 17500 15506 17552 15512
rect 16672 15438 16724 15444
rect 16684 14346 16712 15438
rect 17144 15422 17356 15450
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16578 13560 16634 13569
rect 16396 13524 16448 13530
rect 16578 13495 16634 13504
rect 16396 13466 16448 13472
rect 16394 13424 16450 13433
rect 16394 13359 16450 13368
rect 16408 12782 16436 13359
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16396 12776 16448 12782
rect 16394 12744 16396 12753
rect 16448 12744 16450 12753
rect 16394 12679 16450 12688
rect 16592 11880 16620 12786
rect 16868 12102 16896 14758
rect 16948 14408 17000 14414
rect 16946 14376 16948 14385
rect 17000 14376 17002 14385
rect 16946 14311 17002 14320
rect 17144 13954 17172 15422
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17052 13926 17172 13954
rect 17052 12850 17080 13926
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17052 12646 17080 12786
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16672 11892 16724 11898
rect 16592 11852 16672 11880
rect 16672 11834 16724 11840
rect 16580 11688 16632 11694
rect 16632 11636 16804 11642
rect 16580 11630 16804 11636
rect 16592 11614 16804 11630
rect 17144 11626 17172 13806
rect 17236 12986 17264 13806
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 16040 11104 16344 11132
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15212 10254 15424 10282
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 14554 9616 14610 9625
rect 14554 9551 14556 9560
rect 14608 9551 14610 9560
rect 14556 9522 14608 9528
rect 14568 9491 14596 9522
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 15028 9178 15056 9386
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15028 8906 15056 9114
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 15028 8498 15056 8842
rect 15212 8634 15240 9998
rect 15304 9178 15332 10066
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 15304 8362 15332 8774
rect 15396 8362 15424 10254
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15764 8634 15792 8910
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 16040 8022 16068 11104
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16592 10742 16620 11018
rect 16580 10736 16632 10742
rect 16210 10704 16266 10713
rect 16580 10678 16632 10684
rect 16210 10639 16266 10648
rect 16224 10470 16252 10639
rect 16776 10538 16804 11614
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 16868 11354 16896 11562
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16868 10674 16896 11290
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16960 10606 16988 10950
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16764 10532 16816 10538
rect 16764 10474 16816 10480
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16132 10266 16160 10406
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16224 9722 16252 10066
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16316 9625 16344 9998
rect 16408 9654 16436 10134
rect 16670 9752 16726 9761
rect 16670 9687 16726 9696
rect 16396 9648 16448 9654
rect 16302 9616 16358 9625
rect 16396 9590 16448 9596
rect 16302 9551 16358 9560
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 16316 7954 16344 9551
rect 16684 9382 16712 9687
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16500 9178 16528 9318
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16960 9110 16988 9522
rect 16948 9104 17000 9110
rect 16948 9046 17000 9052
rect 16960 8974 16988 9046
rect 17144 9042 17172 11562
rect 17236 9722 17264 12786
rect 17328 12714 17356 15302
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17420 14550 17448 14758
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 17512 13938 17540 14826
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17498 13152 17554 13161
rect 17498 13087 17554 13096
rect 17512 12850 17540 13087
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17316 12708 17368 12714
rect 17316 12650 17368 12656
rect 17512 12442 17540 12786
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17604 12374 17632 15438
rect 17408 12368 17460 12374
rect 17592 12368 17644 12374
rect 17408 12310 17460 12316
rect 17498 12336 17554 12345
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17328 10198 17356 12242
rect 17420 11558 17448 12310
rect 17696 12345 17724 15558
rect 18604 15564 18656 15570
rect 18708 15558 18828 15586
rect 18604 15506 18656 15512
rect 18512 15428 18564 15434
rect 18512 15370 18564 15376
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17972 15065 18000 15098
rect 17958 15056 18014 15065
rect 17958 14991 18014 15000
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17788 14385 17816 14894
rect 18524 14890 18552 15370
rect 18512 14884 18564 14890
rect 18512 14826 18564 14832
rect 17960 14816 18012 14822
rect 17880 14764 17960 14770
rect 17880 14758 18012 14764
rect 17880 14742 18000 14758
rect 17774 14376 17830 14385
rect 17774 14311 17830 14320
rect 17788 13734 17816 14311
rect 17880 14074 17908 14742
rect 18524 14618 18552 14826
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17788 13394 17816 13670
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 17776 12368 17828 12374
rect 17592 12310 17644 12316
rect 17682 12336 17738 12345
rect 17498 12271 17554 12280
rect 17776 12310 17828 12316
rect 17682 12271 17738 12280
rect 17512 12238 17540 12271
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17684 11824 17736 11830
rect 17684 11766 17736 11772
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17420 10810 17448 11494
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16684 8430 16712 8842
rect 16960 8498 16988 8910
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 17420 8430 17448 9658
rect 17604 9160 17632 11290
rect 17696 11150 17724 11766
rect 17788 11354 17816 12310
rect 17880 11393 17908 13738
rect 17972 12918 18000 14010
rect 18236 14000 18288 14006
rect 18234 13968 18236 13977
rect 18288 13968 18290 13977
rect 18616 13954 18644 15506
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18708 14618 18736 15438
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18800 14482 18828 15558
rect 18892 14498 18920 16487
rect 18984 16454 19012 17224
rect 19156 17206 19208 17212
rect 19352 17202 19380 17439
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19444 16998 19472 18022
rect 19536 18006 19656 18034
rect 19536 17785 19564 18006
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19522 17776 19578 17785
rect 19522 17711 19578 17720
rect 19522 17640 19578 17649
rect 19522 17575 19578 17584
rect 19536 17134 19564 17575
rect 19628 17354 19656 17818
rect 19720 17542 19748 20318
rect 19996 18170 20024 22320
rect 20166 20632 20222 20641
rect 20166 20567 20222 20576
rect 20180 20058 20208 20567
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 19904 18142 20024 18170
rect 19904 17814 19932 18142
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19892 17808 19944 17814
rect 19892 17750 19944 17756
rect 19708 17536 19760 17542
rect 19892 17536 19944 17542
rect 19708 17478 19760 17484
rect 19812 17484 19892 17490
rect 19812 17478 19944 17484
rect 19812 17462 19932 17478
rect 19628 17326 19748 17354
rect 19614 17232 19670 17241
rect 19614 17167 19670 17176
rect 19628 17134 19656 17167
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 19076 15910 19104 16594
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 18984 14618 19012 15846
rect 19076 15570 19104 15846
rect 19064 15564 19116 15570
rect 19064 15506 19116 15512
rect 19168 15434 19196 16934
rect 19524 16788 19576 16794
rect 19628 16776 19656 16934
rect 19576 16748 19656 16776
rect 19524 16730 19576 16736
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19260 15586 19288 16594
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19260 15558 19380 15586
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19156 15428 19208 15434
rect 19156 15370 19208 15376
rect 18972 14612 19024 14618
rect 18972 14554 19024 14560
rect 18788 14476 18840 14482
rect 18892 14470 19012 14498
rect 18788 14418 18840 14424
rect 18880 14340 18932 14346
rect 18880 14282 18932 14288
rect 18234 13903 18290 13912
rect 18524 13926 18644 13954
rect 18234 13696 18290 13705
rect 18234 13631 18290 13640
rect 18248 13394 18276 13631
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 17960 12912 18012 12918
rect 17960 12854 18012 12860
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 18064 12084 18092 12854
rect 17972 12056 18092 12084
rect 17866 11384 17922 11393
rect 17776 11348 17828 11354
rect 17866 11319 17922 11328
rect 17776 11290 17828 11296
rect 17972 11234 18000 12056
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18420 11688 18472 11694
rect 18418 11656 18420 11665
rect 18472 11656 18474 11665
rect 18418 11591 18474 11600
rect 18432 11354 18460 11591
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 17880 11206 18000 11234
rect 17684 11144 17736 11150
rect 17880 11098 17908 11206
rect 17684 11086 17736 11092
rect 17696 10169 17724 11086
rect 17788 11070 17908 11098
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17788 10674 17816 11070
rect 17868 11008 17920 11014
rect 17866 10976 17868 10985
rect 17920 10976 17922 10985
rect 17866 10911 17922 10920
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 17682 10160 17738 10169
rect 17682 10095 17738 10104
rect 17696 9994 17724 10095
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17788 9178 17816 10474
rect 17972 10418 18000 11086
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18524 10810 18552 13926
rect 18604 13728 18656 13734
rect 18604 13670 18656 13676
rect 18786 13696 18842 13705
rect 18616 12850 18644 13670
rect 18786 13631 18842 13640
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18800 11778 18828 13631
rect 18892 12918 18920 14282
rect 18984 13734 19012 14470
rect 19260 14074 19288 15438
rect 19352 14822 19380 15558
rect 19444 15162 19472 15914
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19062 13832 19118 13841
rect 19062 13767 19118 13776
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 18984 12986 19012 13262
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 19076 12918 19104 13767
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 18880 12912 18932 12918
rect 19064 12912 19116 12918
rect 18880 12854 18932 12860
rect 18970 12880 19026 12889
rect 19064 12854 19116 12860
rect 18970 12815 19026 12824
rect 18984 12730 19012 12815
rect 18708 11750 18828 11778
rect 18892 12702 19012 12730
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18708 10606 18736 11750
rect 18892 11642 18920 12702
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 18800 11614 18920 11642
rect 18800 11354 18828 11614
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18892 10810 18920 11494
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18878 10704 18934 10713
rect 18878 10639 18880 10648
rect 18932 10639 18934 10648
rect 18880 10610 18932 10616
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 17880 10390 18000 10418
rect 17776 9172 17828 9178
rect 17604 9132 17724 9160
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 14370 7848 14426 7857
rect 14370 7783 14426 7792
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11992 5302 12020 7142
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 16684 6866 16712 7890
rect 17144 7410 17172 7890
rect 17420 7546 17448 8230
rect 17512 8090 17540 8434
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 11980 5296 12032 5302
rect 11610 5264 11666 5273
rect 11980 5238 12032 5244
rect 11610 5199 11666 5208
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 11164 1986 11192 2926
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11164 1958 11376 1986
rect 11348 480 11376 1958
rect 15856 480 15884 2926
rect 17604 2553 17632 8978
rect 17696 7206 17724 9132
rect 17776 9114 17828 9120
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17590 2544 17646 2553
rect 17590 2479 17646 2488
rect 17788 1601 17816 9114
rect 17880 9110 17908 10390
rect 18156 10266 18184 10542
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18418 10296 18474 10305
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18144 10260 18196 10266
rect 18418 10231 18474 10240
rect 18144 10202 18196 10208
rect 17868 9104 17920 9110
rect 17972 9081 18000 10202
rect 18432 10130 18460 10231
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18515 9846 18552 9862
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18524 9654 18552 9846
rect 18708 9654 18736 9998
rect 18512 9648 18564 9654
rect 18512 9590 18564 9596
rect 18696 9648 18748 9654
rect 18696 9590 18748 9596
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 17868 9046 17920 9052
rect 17958 9072 18014 9081
rect 17958 9007 18014 9016
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17880 8430 17908 8910
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17972 7546 18000 8298
rect 18064 8022 18092 8366
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18340 8090 18368 8298
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18052 8016 18104 8022
rect 18052 7958 18104 7964
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 18064 7002 18092 7346
rect 18432 7274 18460 7414
rect 18420 7268 18472 7274
rect 18420 7210 18472 7216
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 5817 18000 6598
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 17958 5808 18014 5817
rect 17958 5743 18014 5752
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17972 4865 18000 5306
rect 17958 4856 18014 4865
rect 17958 4791 18014 4800
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17774 1592 17830 1601
rect 17774 1527 17830 1536
rect 18708 649 18736 9454
rect 18800 6769 18828 10406
rect 18970 10296 19026 10305
rect 18970 10231 18972 10240
rect 19024 10231 19026 10240
rect 18972 10202 19024 10208
rect 18880 9988 18932 9994
rect 18932 9948 19104 9976
rect 18880 9930 18932 9936
rect 18970 9888 19026 9897
rect 18970 9823 19026 9832
rect 18878 9752 18934 9761
rect 18878 9687 18934 9696
rect 18892 8129 18920 9687
rect 18984 9586 19012 9823
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18878 8120 18934 8129
rect 18878 8055 18934 8064
rect 19076 7478 19104 9948
rect 19168 9489 19196 12038
rect 19260 11898 19288 13670
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19246 11520 19302 11529
rect 19246 11455 19302 11464
rect 19154 9480 19210 9489
rect 19154 9415 19210 9424
rect 19156 8016 19208 8022
rect 19156 7958 19208 7964
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 18786 6760 18842 6769
rect 18786 6695 18842 6704
rect 18892 1057 18920 7414
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 18878 1048 18934 1057
rect 18878 983 18934 992
rect 18694 640 18750 649
rect 18694 575 18750 584
rect 7562 232 7618 241
rect 7562 167 7618 176
rect 11334 0 11390 480
rect 15842 0 15898 480
rect 19076 241 19104 7142
rect 19168 6798 19196 7958
rect 19260 7177 19288 11455
rect 19352 11354 19380 14350
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19444 13190 19472 13806
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19444 12850 19472 13126
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19536 12714 19564 15982
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19628 14618 19656 15302
rect 19720 14890 19748 17326
rect 19812 17202 19840 17462
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19708 14884 19760 14890
rect 19708 14826 19760 14832
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19628 12442 19656 13330
rect 19720 13190 19748 13874
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 19720 12238 19748 13126
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19536 10606 19564 11494
rect 19616 11144 19668 11150
rect 19616 11086 19668 11092
rect 19628 10674 19656 11086
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19432 10464 19484 10470
rect 19628 10452 19656 10610
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19432 10406 19484 10412
rect 19536 10424 19656 10452
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19352 9518 19380 10066
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19444 9450 19472 10406
rect 19536 10169 19564 10424
rect 19616 10192 19668 10198
rect 19522 10160 19578 10169
rect 19616 10134 19668 10140
rect 19522 10095 19578 10104
rect 19536 10062 19564 10095
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19352 9042 19380 9318
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19444 8634 19472 9046
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19536 8090 19564 9318
rect 19628 9110 19656 10134
rect 19720 9654 19748 10542
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19720 8634 19748 9318
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19812 7868 19840 17138
rect 19904 14090 19932 17274
rect 19996 17202 20024 18022
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19996 14278 20024 16594
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19904 14062 20024 14090
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19904 13462 19932 13670
rect 19892 13456 19944 13462
rect 19996 13433 20024 14062
rect 19892 13398 19944 13404
rect 19982 13424 20038 13433
rect 19982 13359 20038 13368
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19996 12442 20024 12582
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19996 10810 20024 11630
rect 20088 11286 20116 19246
rect 20456 18873 20484 22320
rect 20626 21584 20682 21593
rect 20626 21519 20682 21528
rect 20640 20058 20668 21519
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20626 19272 20682 19281
rect 20442 18864 20498 18873
rect 20442 18799 20498 18808
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20180 18290 20208 18566
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20180 17338 20208 18022
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20272 16998 20300 18158
rect 20548 18086 20576 19246
rect 20626 19207 20682 19216
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20534 17504 20590 17513
rect 20534 17439 20590 17448
rect 20548 17134 20576 17439
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20168 15564 20220 15570
rect 20168 15506 20220 15512
rect 20180 13297 20208 15506
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20272 15162 20300 15438
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 20166 13288 20222 13297
rect 20166 13223 20222 13232
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20180 12238 20208 12786
rect 20272 12782 20300 13670
rect 20364 12918 20392 14758
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20352 12912 20404 12918
rect 20352 12854 20404 12860
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20456 12374 20484 13806
rect 20548 13530 20576 15982
rect 20640 15162 20668 19207
rect 20732 19174 20760 22471
rect 20902 22320 20958 22800
rect 21270 22320 21326 22800
rect 21730 22320 21786 22800
rect 22098 22320 22154 22800
rect 22558 22320 22614 22800
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20810 18864 20866 18873
rect 20810 18799 20866 18808
rect 20824 18426 20852 18799
rect 20916 18737 20944 22320
rect 20902 18728 20958 18737
rect 20902 18663 20958 18672
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 21284 17241 21312 22320
rect 21744 19145 21772 22320
rect 22112 19242 22140 22320
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 21730 19136 21786 19145
rect 21730 19071 21786 19080
rect 22190 18184 22246 18193
rect 22572 18170 22600 22320
rect 22246 18142 22600 18170
rect 22190 18119 22246 18128
rect 21270 17232 21326 17241
rect 21270 17167 21326 17176
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20812 15972 20864 15978
rect 20812 15914 20864 15920
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20536 13524 20588 13530
rect 20536 13466 20588 13472
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20548 12850 20576 13126
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20444 12368 20496 12374
rect 20444 12310 20496 12316
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20548 11626 20576 12242
rect 20536 11620 20588 11626
rect 20536 11562 20588 11568
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 20076 11280 20128 11286
rect 20076 11222 20128 11228
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19996 10130 20024 10746
rect 20076 10532 20128 10538
rect 20076 10474 20128 10480
rect 20088 10266 20116 10474
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19904 8838 19932 9522
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19996 8650 20024 10066
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 19904 8622 20024 8650
rect 19904 8294 19932 8622
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 19892 8288 19944 8294
rect 19892 8230 19944 8236
rect 19996 7886 20024 8502
rect 20088 8430 20116 9862
rect 20180 9722 20208 11494
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20180 9518 20208 9658
rect 20272 9654 20300 10202
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20260 9648 20312 9654
rect 20260 9590 20312 9596
rect 20364 9586 20392 9998
rect 20548 9602 20576 11562
rect 20640 11354 20668 14418
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20732 10656 20760 13670
rect 20824 13258 20852 15914
rect 20916 15706 20944 16526
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20994 14104 21050 14113
rect 20994 14039 21050 14048
rect 20812 13252 20864 13258
rect 20812 13194 20864 13200
rect 20904 12708 20956 12714
rect 20904 12650 20956 12656
rect 20916 12442 20944 12650
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20732 10628 20852 10656
rect 20626 10568 20682 10577
rect 20626 10503 20682 10512
rect 20720 10532 20772 10538
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20456 9574 20576 9602
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 19720 7840 19840 7868
rect 19892 7880 19944 7886
rect 19246 7168 19302 7177
rect 19246 7103 19302 7112
rect 19720 6866 19748 7840
rect 19892 7822 19944 7828
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19904 7546 19932 7822
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19168 6322 19196 6734
rect 19260 6458 19288 6802
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19812 5914 19840 7278
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 20088 2961 20116 8230
rect 20180 8090 20208 9318
rect 20364 8362 20392 9522
rect 20352 8356 20404 8362
rect 20352 8298 20404 8304
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20364 7410 20392 8298
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20456 7206 20484 9574
rect 20640 9518 20668 10503
rect 20720 10474 20772 10480
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20548 9178 20576 9318
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20640 9058 20668 9318
rect 20548 9030 20668 9058
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20180 5914 20208 6734
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20364 5710 20392 6394
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20272 5370 20300 5646
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20456 3913 20484 7142
rect 20548 5114 20576 9030
rect 20732 8430 20760 10474
rect 20824 10266 20852 10628
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 21008 8634 21036 14039
rect 21088 12912 21140 12918
rect 21088 12854 21140 12860
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 21100 8537 21128 12854
rect 21364 9648 21416 9654
rect 21364 9590 21416 9596
rect 21086 8528 21142 8537
rect 21086 8463 21142 8472
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20640 6186 20668 6598
rect 20628 6180 20680 6186
rect 20628 6122 20680 6128
rect 20640 5234 20668 6122
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20548 5086 20668 5114
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20548 4321 20576 4966
rect 20534 4312 20590 4321
rect 20534 4247 20590 4256
rect 20442 3904 20498 3913
rect 20442 3839 20498 3848
rect 20640 3505 20668 5086
rect 20626 3496 20682 3505
rect 20626 3431 20682 3440
rect 20074 2952 20130 2961
rect 20074 2887 20130 2896
rect 20444 2916 20496 2922
rect 20444 2858 20496 2864
rect 20456 480 20484 2858
rect 21376 2009 21404 9590
rect 21362 2000 21418 2009
rect 21362 1935 21418 1944
rect 19062 232 19118 241
rect 19062 167 19118 176
rect 20442 0 20498 480
<< via2 >>
rect 3054 22480 3110 22536
rect 1398 19080 1454 19136
rect 1950 19760 2006 19816
rect 1858 18944 1914 19000
rect 1950 18808 2006 18864
rect 1950 18264 2006 18320
rect 1950 17332 2006 17368
rect 1950 17312 1952 17332
rect 1952 17312 2004 17332
rect 2004 17312 2006 17332
rect 2410 19080 2466 19136
rect 2318 17992 2374 18048
rect 1950 16904 2006 16960
rect 1950 16496 2006 16552
rect 1950 15952 2006 16008
rect 1950 15544 2006 15600
rect 1766 14048 1822 14104
rect 2594 18264 2650 18320
rect 2502 17720 2558 17776
rect 2962 22072 3018 22128
rect 2778 21528 2834 21584
rect 2870 20576 2926 20632
rect 2778 19216 2834 19272
rect 20718 22480 20774 22536
rect 3422 20168 3478 20224
rect 3146 19216 3202 19272
rect 2778 17856 2834 17912
rect 2778 16088 2834 16144
rect 2778 15000 2834 15056
rect 2318 13232 2374 13288
rect 3238 18692 3294 18728
rect 3238 18672 3240 18692
rect 3240 18672 3292 18692
rect 3292 18672 3294 18692
rect 3146 17584 3202 17640
rect 3146 14592 3202 14648
rect 3146 13640 3202 13696
rect 2870 7520 2926 7576
rect 1858 2488 1914 2544
rect 3698 21120 3754 21176
rect 2870 4256 2926 4312
rect 3514 12688 3570 12744
rect 3514 12552 3570 12608
rect 3698 16632 3754 16688
rect 3698 12824 3754 12880
rect 3606 11328 3662 11384
rect 3514 7112 3570 7168
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4250 18808 4306 18864
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4802 18400 4858 18456
rect 4066 16768 4122 16824
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4066 12316 4068 12336
rect 4068 12316 4120 12336
rect 4120 12316 4122 12336
rect 4066 12280 4122 12316
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4066 11736 4122 11792
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 3974 10784 4030 10840
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 3882 9424 3938 9480
rect 4066 9016 4122 9072
rect 4066 8472 4122 8528
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4710 9016 4766 9072
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4802 8916 4804 8936
rect 4804 8916 4856 8936
rect 4856 8916 4858 8936
rect 4802 8880 4858 8916
rect 4802 8492 4858 8528
rect 4802 8472 4804 8492
rect 4804 8472 4856 8492
rect 4856 8472 4858 8492
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4066 6704 4122 6760
rect 3974 6160 4030 6216
rect 3422 5752 3478 5808
rect 4066 5244 4068 5264
rect 4068 5244 4120 5264
rect 4120 5244 4122 5264
rect 4066 5208 4122 5244
rect 4066 4800 4122 4856
rect 4158 3848 4214 3904
rect 3330 3440 3386 3496
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 4250 1944 4306 2000
rect 2778 1536 2834 1592
rect 5538 18536 5594 18592
rect 6550 18536 6606 18592
rect 6274 18128 6330 18184
rect 5170 9016 5226 9072
rect 5078 8084 5134 8120
rect 5078 8064 5080 8084
rect 5080 8064 5132 8084
rect 5132 8064 5134 8084
rect 5354 9052 5356 9072
rect 5356 9052 5408 9072
rect 5408 9052 5410 9072
rect 5354 9016 5410 9052
rect 5538 8472 5594 8528
rect 5354 7964 5356 7984
rect 5356 7964 5408 7984
rect 5408 7964 5410 7984
rect 5354 7928 5410 7964
rect 5998 14048 6054 14104
rect 6182 17992 6238 18048
rect 6366 15408 6422 15464
rect 6366 10512 6422 10568
rect 6826 18944 6882 19000
rect 7286 19080 7342 19136
rect 6734 17176 6790 17232
rect 7010 17040 7066 17096
rect 7194 15952 7250 16008
rect 7194 15680 7250 15736
rect 6550 10104 6606 10160
rect 6458 8064 6514 8120
rect 4802 2896 4858 2952
rect 6550 992 6606 1048
rect 2778 584 2834 640
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7746 18400 7802 18456
rect 7378 17040 7434 17096
rect 8482 18536 8538 18592
rect 8574 18400 8630 18456
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 8206 17176 8262 17232
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7562 15952 7618 16008
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 8114 15564 8170 15600
rect 8114 15544 8116 15564
rect 8116 15544 8168 15564
rect 8168 15544 8170 15564
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7286 8880 7342 8936
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7930 8880 7986 8936
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 8666 17992 8722 18048
rect 8666 17312 8722 17368
rect 9310 18400 9366 18456
rect 9310 17756 9312 17776
rect 9312 17756 9364 17776
rect 9364 17756 9366 17776
rect 9310 17720 9366 17756
rect 9586 17584 9642 17640
rect 9586 17332 9642 17368
rect 9586 17312 9588 17332
rect 9588 17312 9640 17332
rect 9640 17312 9642 17332
rect 9586 16768 9642 16824
rect 9218 16088 9274 16144
rect 9678 15408 9734 15464
rect 9678 14612 9734 14648
rect 9678 14592 9680 14612
rect 9680 14592 9732 14612
rect 9732 14592 9734 14612
rect 9310 13368 9366 13424
rect 9770 14320 9826 14376
rect 9770 14184 9826 14240
rect 8666 9968 8722 10024
rect 10322 17312 10378 17368
rect 10598 17312 10654 17368
rect 10414 15408 10470 15464
rect 10138 13776 10194 13832
rect 10138 11328 10194 11384
rect 9126 8916 9128 8936
rect 9128 8916 9180 8936
rect 9180 8916 9182 8936
rect 9126 8880 9182 8916
rect 10506 14456 10562 14512
rect 10506 14356 10508 14376
rect 10508 14356 10560 14376
rect 10560 14356 10562 14376
rect 10506 14320 10562 14356
rect 10322 10648 10378 10704
rect 10966 18944 11022 19000
rect 10782 17992 10838 18048
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 10966 17176 11022 17232
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 12070 18148 12126 18184
rect 12070 18128 12072 18148
rect 12072 18128 12124 18148
rect 12124 18128 12126 18148
rect 11518 16940 11520 16960
rect 11520 16940 11572 16960
rect 11572 16940 11574 16960
rect 11518 16904 11574 16940
rect 11886 16768 11942 16824
rect 10782 11600 10838 11656
rect 10690 10920 10746 10976
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11334 13232 11390 13288
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11058 11600 11114 11656
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11334 11600 11390 11656
rect 10966 11056 11022 11112
rect 11426 11056 11482 11112
rect 11978 12008 12034 12064
rect 11610 11192 11666 11248
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11242 10512 11298 10568
rect 11150 9968 11206 10024
rect 11518 10240 11574 10296
rect 11794 11464 11850 11520
rect 11702 10648 11758 10704
rect 11794 10512 11850 10568
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11518 9444 11574 9480
rect 11518 9424 11520 9444
rect 11520 9424 11572 9444
rect 11572 9424 11574 9444
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11978 10920 12034 10976
rect 11886 9968 11942 10024
rect 11794 9716 11850 9752
rect 11794 9696 11796 9716
rect 11796 9696 11848 9716
rect 11848 9696 11850 9716
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 10138 6160 10194 6216
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 12254 12960 12310 13016
rect 12622 18944 12678 19000
rect 12530 17756 12532 17776
rect 12532 17756 12584 17776
rect 12584 17756 12586 17776
rect 12530 17720 12586 17756
rect 12622 17620 12624 17640
rect 12624 17620 12676 17640
rect 12676 17620 12678 17640
rect 12622 17584 12678 17620
rect 12530 17212 12532 17232
rect 12532 17212 12584 17232
rect 12584 17212 12586 17232
rect 12530 17176 12586 17212
rect 12714 17040 12770 17096
rect 13450 18148 13506 18184
rect 13450 18128 13452 18148
rect 13452 18128 13504 18148
rect 13504 18128 13506 18148
rect 13542 17992 13598 18048
rect 13358 17584 13414 17640
rect 13082 15408 13138 15464
rect 12438 12144 12494 12200
rect 12346 12008 12402 12064
rect 12622 10920 12678 10976
rect 12438 10240 12494 10296
rect 13082 14456 13138 14512
rect 13174 12688 13230 12744
rect 13542 16940 13544 16960
rect 13544 16940 13596 16960
rect 13596 16940 13598 16960
rect 13542 16904 13598 16940
rect 13818 12280 13874 12336
rect 12806 11092 12808 11112
rect 12808 11092 12860 11112
rect 12860 11092 12862 11112
rect 12806 11056 12862 11092
rect 13542 11056 13598 11112
rect 12438 8472 12494 8528
rect 13450 8492 13506 8528
rect 13450 8472 13452 8492
rect 13452 8472 13504 8492
rect 13504 8472 13506 8492
rect 14278 17856 14334 17912
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14554 17720 14610 17776
rect 14370 17196 14426 17232
rect 14370 17176 14372 17196
rect 14372 17176 14424 17196
rect 14424 17176 14426 17196
rect 14278 16632 14334 16688
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 15566 18128 15622 18184
rect 15750 17040 15806 17096
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 15198 13676 15200 13696
rect 15200 13676 15252 13696
rect 15252 13676 15254 13696
rect 15198 13640 15254 13676
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14094 9424 14150 9480
rect 15934 15544 15990 15600
rect 17314 17720 17370 17776
rect 16302 16496 16358 16552
rect 16302 16088 16358 16144
rect 16210 14864 16266 14920
rect 16118 14320 16174 14376
rect 16026 13524 16082 13560
rect 16026 13504 16028 13524
rect 16028 13504 16080 13524
rect 16080 13504 16082 13524
rect 15474 12824 15530 12880
rect 15382 12008 15438 12064
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 15750 12180 15752 12200
rect 15752 12180 15804 12200
rect 15804 12180 15806 12200
rect 15750 12144 15806 12180
rect 15474 11464 15530 11520
rect 16210 12552 16266 12608
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18970 22072 19026 22128
rect 18878 18028 18880 18048
rect 18880 18028 18932 18048
rect 18932 18028 18934 18048
rect 18878 17992 18934 18028
rect 18602 17876 18658 17912
rect 18602 17856 18604 17876
rect 18604 17856 18656 17876
rect 18656 17856 18658 17876
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18050 17176 18106 17232
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 19154 21120 19210 21176
rect 19062 19780 19118 19816
rect 19062 19760 19064 19780
rect 19064 19760 19116 19780
rect 19116 19760 19118 19780
rect 19614 20168 19670 20224
rect 19338 17584 19394 17640
rect 19338 17448 19394 17504
rect 18878 16496 18934 16552
rect 16578 13504 16634 13560
rect 16394 13368 16450 13424
rect 16394 12724 16396 12744
rect 16396 12724 16448 12744
rect 16448 12724 16450 12744
rect 16394 12688 16450 12724
rect 16946 14356 16948 14376
rect 16948 14356 17000 14376
rect 17000 14356 17002 14376
rect 16946 14320 17002 14356
rect 14554 9580 14610 9616
rect 14554 9560 14556 9580
rect 14556 9560 14608 9580
rect 14608 9560 14610 9580
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 16210 10648 16266 10704
rect 16670 9696 16726 9752
rect 16302 9560 16358 9616
rect 17498 13096 17554 13152
rect 17498 12280 17554 12336
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 17958 15000 18014 15056
rect 17774 14320 17830 14376
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 17682 12280 17738 12336
rect 18234 13948 18236 13968
rect 18236 13948 18288 13968
rect 18288 13948 18290 13968
rect 19522 17720 19578 17776
rect 19522 17584 19578 17640
rect 20166 20576 20222 20632
rect 19614 17176 19670 17232
rect 18234 13912 18290 13948
rect 18234 13640 18290 13696
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 17866 11328 17922 11384
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18418 11636 18420 11656
rect 18420 11636 18472 11656
rect 18472 11636 18474 11656
rect 18418 11600 18474 11636
rect 17866 10956 17868 10976
rect 17868 10956 17920 10976
rect 17920 10956 17922 10976
rect 17866 10920 17922 10956
rect 17682 10104 17738 10160
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18786 13640 18842 13696
rect 19062 13776 19118 13832
rect 18970 12824 19026 12880
rect 18878 10668 18934 10704
rect 18878 10648 18880 10668
rect 18880 10648 18932 10668
rect 18932 10648 18934 10668
rect 14370 7792 14426 7848
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 11610 5208 11666 5264
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 17590 2488 17646 2544
rect 18418 10240 18474 10296
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 17958 9016 18014 9072
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 17958 5752 18014 5808
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 17958 4800 18014 4856
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 17774 1536 17830 1592
rect 18970 10260 19026 10296
rect 18970 10240 18972 10260
rect 18972 10240 19024 10260
rect 19024 10240 19026 10260
rect 18970 9832 19026 9888
rect 18878 9696 18934 9752
rect 18878 8064 18934 8120
rect 19246 11464 19302 11520
rect 19154 9424 19210 9480
rect 18786 6704 18842 6760
rect 18878 992 18934 1048
rect 18694 584 18750 640
rect 7562 176 7618 232
rect 19522 10104 19578 10160
rect 19982 13368 20038 13424
rect 20626 21528 20682 21584
rect 20442 18808 20498 18864
rect 20626 19216 20682 19272
rect 20534 17448 20590 17504
rect 20166 13232 20222 13288
rect 20810 18808 20866 18864
rect 20902 18672 20958 18728
rect 21730 19080 21786 19136
rect 22190 18128 22246 18184
rect 21270 17176 21326 17232
rect 20994 14048 21050 14104
rect 20626 10512 20682 10568
rect 19246 7112 19302 7168
rect 21086 8472 21142 8528
rect 20534 4256 20590 4312
rect 20442 3848 20498 3904
rect 20626 3440 20682 3496
rect 20074 2896 20130 2952
rect 21362 1944 21418 2000
rect 19062 176 19118 232
<< metal3 >>
rect 0 22538 480 22568
rect 3049 22538 3115 22541
rect 0 22536 3115 22538
rect 0 22480 3054 22536
rect 3110 22480 3115 22536
rect 0 22478 3115 22480
rect 0 22448 480 22478
rect 3049 22475 3115 22478
rect 20713 22538 20779 22541
rect 22320 22538 22800 22568
rect 20713 22536 22800 22538
rect 20713 22480 20718 22536
rect 20774 22480 22800 22536
rect 20713 22478 22800 22480
rect 20713 22475 20779 22478
rect 22320 22448 22800 22478
rect 0 22130 480 22160
rect 2957 22130 3023 22133
rect 0 22128 3023 22130
rect 0 22072 2962 22128
rect 3018 22072 3023 22128
rect 0 22070 3023 22072
rect 0 22040 480 22070
rect 2957 22067 3023 22070
rect 18965 22130 19031 22133
rect 22320 22130 22800 22160
rect 18965 22128 22800 22130
rect 18965 22072 18970 22128
rect 19026 22072 22800 22128
rect 18965 22070 22800 22072
rect 18965 22067 19031 22070
rect 22320 22040 22800 22070
rect 0 21586 480 21616
rect 2773 21586 2839 21589
rect 0 21584 2839 21586
rect 0 21528 2778 21584
rect 2834 21528 2839 21584
rect 0 21526 2839 21528
rect 0 21496 480 21526
rect 2773 21523 2839 21526
rect 20621 21586 20687 21589
rect 22320 21586 22800 21616
rect 20621 21584 22800 21586
rect 20621 21528 20626 21584
rect 20682 21528 22800 21584
rect 20621 21526 22800 21528
rect 20621 21523 20687 21526
rect 22320 21496 22800 21526
rect 0 21178 480 21208
rect 3693 21178 3759 21181
rect 0 21176 3759 21178
rect 0 21120 3698 21176
rect 3754 21120 3759 21176
rect 0 21118 3759 21120
rect 0 21088 480 21118
rect 3693 21115 3759 21118
rect 19149 21178 19215 21181
rect 22320 21178 22800 21208
rect 19149 21176 22800 21178
rect 19149 21120 19154 21176
rect 19210 21120 22800 21176
rect 19149 21118 22800 21120
rect 19149 21115 19215 21118
rect 22320 21088 22800 21118
rect 0 20634 480 20664
rect 2865 20634 2931 20637
rect 0 20632 2931 20634
rect 0 20576 2870 20632
rect 2926 20576 2931 20632
rect 0 20574 2931 20576
rect 0 20544 480 20574
rect 2865 20571 2931 20574
rect 20161 20634 20227 20637
rect 22320 20634 22800 20664
rect 20161 20632 22800 20634
rect 20161 20576 20166 20632
rect 20222 20576 22800 20632
rect 20161 20574 22800 20576
rect 20161 20571 20227 20574
rect 22320 20544 22800 20574
rect 0 20226 480 20256
rect 3417 20226 3483 20229
rect 0 20224 3483 20226
rect 0 20168 3422 20224
rect 3478 20168 3483 20224
rect 0 20166 3483 20168
rect 0 20136 480 20166
rect 3417 20163 3483 20166
rect 19609 20226 19675 20229
rect 22320 20226 22800 20256
rect 19609 20224 22800 20226
rect 19609 20168 19614 20224
rect 19670 20168 22800 20224
rect 19609 20166 22800 20168
rect 19609 20163 19675 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 0 19818 480 19848
rect 1945 19818 2011 19821
rect 0 19816 2011 19818
rect 0 19760 1950 19816
rect 2006 19760 2011 19816
rect 0 19758 2011 19760
rect 0 19728 480 19758
rect 1945 19755 2011 19758
rect 19057 19818 19123 19821
rect 22320 19818 22800 19848
rect 19057 19816 22800 19818
rect 19057 19760 19062 19816
rect 19118 19760 22800 19816
rect 19057 19758 22800 19760
rect 19057 19755 19123 19758
rect 22320 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 2773 19274 2839 19277
rect 0 19272 2839 19274
rect 0 19216 2778 19272
rect 2834 19216 2839 19272
rect 0 19214 2839 19216
rect 0 19184 480 19214
rect 2773 19211 2839 19214
rect 3141 19274 3207 19277
rect 20621 19274 20687 19277
rect 22320 19274 22800 19304
rect 3141 19272 17050 19274
rect 3141 19216 3146 19272
rect 3202 19216 17050 19272
rect 3141 19214 17050 19216
rect 3141 19211 3207 19214
rect 1393 19138 1459 19141
rect 2405 19138 2471 19141
rect 7281 19138 7347 19141
rect 1393 19136 7347 19138
rect 1393 19080 1398 19136
rect 1454 19080 2410 19136
rect 2466 19080 7286 19136
rect 7342 19080 7347 19136
rect 1393 19078 7347 19080
rect 16990 19138 17050 19214
rect 20621 19272 22800 19274
rect 20621 19216 20626 19272
rect 20682 19216 22800 19272
rect 20621 19214 22800 19216
rect 20621 19211 20687 19214
rect 22320 19184 22800 19214
rect 21725 19138 21791 19141
rect 16990 19136 21791 19138
rect 16990 19080 21730 19136
rect 21786 19080 21791 19136
rect 16990 19078 21791 19080
rect 1393 19075 1459 19078
rect 2405 19075 2471 19078
rect 7281 19075 7347 19078
rect 21725 19075 21791 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 1853 19002 1919 19005
rect 6821 19002 6887 19005
rect 1853 19000 6887 19002
rect 1853 18944 1858 19000
rect 1914 18944 6826 19000
rect 6882 18944 6887 19000
rect 1853 18942 6887 18944
rect 1853 18939 1919 18942
rect 6821 18939 6887 18942
rect 10961 19002 11027 19005
rect 12617 19002 12683 19005
rect 10961 19000 12683 19002
rect 10961 18944 10966 19000
rect 11022 18944 12622 19000
rect 12678 18944 12683 19000
rect 10961 18942 12683 18944
rect 10961 18939 11027 18942
rect 12617 18939 12683 18942
rect 0 18866 480 18896
rect 1945 18866 2011 18869
rect 0 18864 2011 18866
rect 0 18808 1950 18864
rect 2006 18808 2011 18864
rect 0 18806 2011 18808
rect 0 18776 480 18806
rect 1945 18803 2011 18806
rect 4245 18866 4311 18869
rect 20437 18866 20503 18869
rect 4245 18864 20503 18866
rect 4245 18808 4250 18864
rect 4306 18808 20442 18864
rect 20498 18808 20503 18864
rect 4245 18806 20503 18808
rect 4245 18803 4311 18806
rect 20437 18803 20503 18806
rect 20805 18866 20871 18869
rect 22320 18866 22800 18896
rect 20805 18864 22800 18866
rect 20805 18808 20810 18864
rect 20866 18808 22800 18864
rect 20805 18806 22800 18808
rect 20805 18803 20871 18806
rect 22320 18776 22800 18806
rect 3233 18730 3299 18733
rect 20897 18730 20963 18733
rect 3233 18728 20963 18730
rect 3233 18672 3238 18728
rect 3294 18672 20902 18728
rect 20958 18672 20963 18728
rect 3233 18670 20963 18672
rect 3233 18667 3299 18670
rect 20897 18667 20963 18670
rect 5533 18594 5599 18597
rect 6545 18594 6611 18597
rect 8477 18594 8543 18597
rect 5533 18592 8543 18594
rect 5533 18536 5538 18592
rect 5594 18536 6550 18592
rect 6606 18536 8482 18592
rect 8538 18536 8543 18592
rect 5533 18534 8543 18536
rect 5533 18531 5599 18534
rect 6545 18531 6611 18534
rect 8477 18531 8543 18534
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 4797 18460 4863 18461
rect 4797 18456 4844 18460
rect 4908 18458 4914 18460
rect 7741 18458 7807 18461
rect 8334 18458 8340 18460
rect 4797 18400 4802 18456
rect 4797 18396 4844 18400
rect 4908 18398 4954 18458
rect 7741 18456 8340 18458
rect 7741 18400 7746 18456
rect 7802 18400 8340 18456
rect 7741 18398 8340 18400
rect 4908 18396 4914 18398
rect 4797 18395 4863 18396
rect 7741 18395 7807 18398
rect 8334 18396 8340 18398
rect 8404 18396 8410 18460
rect 8569 18458 8635 18461
rect 9305 18458 9371 18461
rect 8569 18456 9371 18458
rect 8569 18400 8574 18456
rect 8630 18400 9310 18456
rect 9366 18400 9371 18456
rect 8569 18398 9371 18400
rect 8569 18395 8635 18398
rect 9305 18395 9371 18398
rect 0 18322 480 18352
rect 1945 18322 2011 18325
rect 0 18320 2011 18322
rect 0 18264 1950 18320
rect 2006 18264 2011 18320
rect 0 18262 2011 18264
rect 0 18232 480 18262
rect 1945 18259 2011 18262
rect 2589 18322 2655 18325
rect 2589 18320 17602 18322
rect 2589 18264 2594 18320
rect 2650 18264 17602 18320
rect 2589 18262 17602 18264
rect 2589 18259 2655 18262
rect 6269 18186 6335 18189
rect 12065 18186 12131 18189
rect 13445 18186 13511 18189
rect 15561 18186 15627 18189
rect 6269 18184 10794 18186
rect 6269 18128 6274 18184
rect 6330 18128 10794 18184
rect 6269 18126 10794 18128
rect 6269 18123 6335 18126
rect 10734 18053 10794 18126
rect 12065 18184 13511 18186
rect 12065 18128 12070 18184
rect 12126 18128 13450 18184
rect 13506 18128 13511 18184
rect 12065 18126 13511 18128
rect 12065 18123 12131 18126
rect 13445 18123 13511 18126
rect 14552 18184 15627 18186
rect 14552 18128 15566 18184
rect 15622 18128 15627 18184
rect 14552 18126 15627 18128
rect 17542 18186 17602 18262
rect 17902 18260 17908 18324
rect 17972 18322 17978 18324
rect 22320 18322 22800 18352
rect 17972 18262 22800 18322
rect 17972 18260 17978 18262
rect 22320 18232 22800 18262
rect 22185 18186 22251 18189
rect 17542 18184 22251 18186
rect 17542 18128 22190 18184
rect 22246 18128 22251 18184
rect 17542 18126 22251 18128
rect 2313 18050 2379 18053
rect 6177 18050 6243 18053
rect 2313 18048 6243 18050
rect 2313 17992 2318 18048
rect 2374 17992 6182 18048
rect 6238 17992 6243 18048
rect 2313 17990 6243 17992
rect 2313 17987 2379 17990
rect 6177 17987 6243 17990
rect 8661 18050 8727 18053
rect 8661 18048 10656 18050
rect 8661 17992 8666 18048
rect 8722 17992 10656 18048
rect 8661 17990 10656 17992
rect 10734 18048 10843 18053
rect 13537 18052 13603 18053
rect 10734 17992 10782 18048
rect 10838 17992 10843 18048
rect 10734 17990 10843 17992
rect 8661 17987 8727 17990
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 2773 17914 2839 17917
rect 0 17912 2839 17914
rect 0 17856 2778 17912
rect 2834 17856 2839 17912
rect 0 17854 2839 17856
rect 0 17824 480 17854
rect 2773 17851 2839 17854
rect 2497 17778 2563 17781
rect 9305 17778 9371 17781
rect 2497 17776 9371 17778
rect 2497 17720 2502 17776
rect 2558 17720 9310 17776
rect 9366 17720 9371 17776
rect 2497 17718 9371 17720
rect 2497 17715 2563 17718
rect 9305 17715 9371 17718
rect 9438 17716 9444 17780
rect 9508 17778 9514 17780
rect 9768 17778 9828 17990
rect 10596 17914 10656 17990
rect 10777 17987 10843 17990
rect 13486 17988 13492 18052
rect 13556 18050 13603 18052
rect 14552 18050 14612 18126
rect 15561 18123 15627 18126
rect 22185 18123 22251 18126
rect 18873 18052 18939 18053
rect 13556 18048 14612 18050
rect 13598 17992 14612 18048
rect 13556 17990 14612 17992
rect 13556 17988 13603 17990
rect 18822 17988 18828 18052
rect 18892 18050 18939 18052
rect 18892 18048 18984 18050
rect 18934 17992 18984 18048
rect 18892 17990 18984 17992
rect 18892 17988 18939 17990
rect 13537 17987 13603 17988
rect 18873 17987 18939 17988
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 14273 17914 14339 17917
rect 10596 17912 14339 17914
rect 10596 17856 14278 17912
rect 14334 17856 14339 17912
rect 10596 17854 14339 17856
rect 14273 17851 14339 17854
rect 18597 17914 18663 17917
rect 22320 17914 22800 17944
rect 18597 17912 22800 17914
rect 18597 17856 18602 17912
rect 18658 17856 22800 17912
rect 18597 17854 22800 17856
rect 18597 17851 18663 17854
rect 22320 17824 22800 17854
rect 9508 17718 9828 17778
rect 12525 17778 12591 17781
rect 14549 17778 14615 17781
rect 12525 17776 14615 17778
rect 12525 17720 12530 17776
rect 12586 17720 14554 17776
rect 14610 17720 14615 17776
rect 12525 17718 14615 17720
rect 9508 17716 9514 17718
rect 12525 17715 12591 17718
rect 14549 17715 14615 17718
rect 17309 17778 17375 17781
rect 19517 17778 19583 17781
rect 17309 17776 19583 17778
rect 17309 17720 17314 17776
rect 17370 17720 19522 17776
rect 19578 17720 19583 17776
rect 17309 17718 19583 17720
rect 17309 17715 17375 17718
rect 19517 17715 19583 17718
rect 3141 17642 3207 17645
rect 9254 17642 9260 17644
rect 3141 17640 9260 17642
rect 3141 17584 3146 17640
rect 3202 17584 9260 17640
rect 3141 17582 9260 17584
rect 3141 17579 3207 17582
rect 9254 17580 9260 17582
rect 9324 17642 9330 17644
rect 9581 17642 9647 17645
rect 9324 17640 9647 17642
rect 9324 17584 9586 17640
rect 9642 17584 9647 17640
rect 9324 17582 9647 17584
rect 9324 17580 9330 17582
rect 9581 17579 9647 17582
rect 12617 17642 12683 17645
rect 13353 17642 13419 17645
rect 12617 17640 13419 17642
rect 12617 17584 12622 17640
rect 12678 17584 13358 17640
rect 13414 17584 13419 17640
rect 12617 17582 13419 17584
rect 12617 17579 12683 17582
rect 13353 17579 13419 17582
rect 19333 17642 19399 17645
rect 19517 17642 19583 17645
rect 19333 17640 19583 17642
rect 19333 17584 19338 17640
rect 19394 17584 19522 17640
rect 19578 17584 19583 17640
rect 19333 17582 19583 17584
rect 19333 17579 19399 17582
rect 19517 17579 19583 17582
rect 19333 17506 19399 17509
rect 20529 17506 20595 17509
rect 19333 17504 20595 17506
rect 19333 17448 19338 17504
rect 19394 17448 20534 17504
rect 20590 17448 20595 17504
rect 19333 17446 20595 17448
rect 19333 17443 19399 17446
rect 20529 17443 20595 17446
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1945 17370 2011 17373
rect 0 17368 2011 17370
rect 0 17312 1950 17368
rect 2006 17312 2011 17368
rect 0 17310 2011 17312
rect 0 17280 480 17310
rect 1945 17307 2011 17310
rect 8661 17370 8727 17373
rect 9581 17370 9647 17373
rect 8661 17368 9647 17370
rect 8661 17312 8666 17368
rect 8722 17312 9586 17368
rect 9642 17312 9647 17368
rect 8661 17310 9647 17312
rect 8661 17307 8727 17310
rect 9581 17307 9647 17310
rect 10317 17370 10383 17373
rect 10593 17370 10659 17373
rect 22320 17370 22800 17400
rect 10317 17368 10659 17370
rect 10317 17312 10322 17368
rect 10378 17312 10598 17368
rect 10654 17312 10659 17368
rect 10317 17310 10659 17312
rect 10317 17307 10383 17310
rect 10593 17307 10659 17310
rect 18646 17310 22800 17370
rect 6729 17234 6795 17237
rect 8201 17234 8267 17237
rect 10961 17234 11027 17237
rect 12525 17234 12591 17237
rect 6729 17232 10840 17234
rect 6729 17176 6734 17232
rect 6790 17176 8206 17232
rect 8262 17176 10840 17232
rect 6729 17174 10840 17176
rect 6729 17171 6795 17174
rect 8201 17171 8267 17174
rect 7005 17098 7071 17101
rect 7373 17098 7439 17101
rect 7005 17096 7439 17098
rect 7005 17040 7010 17096
rect 7066 17040 7378 17096
rect 7434 17040 7439 17096
rect 7005 17038 7439 17040
rect 10780 17098 10840 17174
rect 10961 17232 12591 17234
rect 10961 17176 10966 17232
rect 11022 17176 12530 17232
rect 12586 17176 12591 17232
rect 10961 17174 12591 17176
rect 10961 17171 11027 17174
rect 12525 17171 12591 17174
rect 14365 17234 14431 17237
rect 18045 17234 18111 17237
rect 14365 17232 18111 17234
rect 14365 17176 14370 17232
rect 14426 17176 18050 17232
rect 18106 17176 18111 17232
rect 14365 17174 18111 17176
rect 14365 17171 14431 17174
rect 18045 17171 18111 17174
rect 12709 17098 12775 17101
rect 10780 17096 12775 17098
rect 10780 17040 12714 17096
rect 12770 17040 12775 17096
rect 10780 17038 12775 17040
rect 7005 17035 7071 17038
rect 7373 17035 7439 17038
rect 12709 17035 12775 17038
rect 15745 17098 15811 17101
rect 18646 17098 18706 17310
rect 22320 17280 22800 17310
rect 19609 17234 19675 17237
rect 21265 17234 21331 17237
rect 19609 17232 21331 17234
rect 19609 17176 19614 17232
rect 19670 17176 21270 17232
rect 21326 17176 21331 17232
rect 19609 17174 21331 17176
rect 19609 17171 19675 17174
rect 21265 17171 21331 17174
rect 15745 17096 18706 17098
rect 15745 17040 15750 17096
rect 15806 17040 18706 17096
rect 15745 17038 18706 17040
rect 15745 17035 15811 17038
rect 0 16962 480 16992
rect 1945 16962 2011 16965
rect 0 16960 2011 16962
rect 0 16904 1950 16960
rect 2006 16904 2011 16960
rect 0 16902 2011 16904
rect 0 16872 480 16902
rect 1945 16899 2011 16902
rect 11513 16962 11579 16965
rect 13537 16962 13603 16965
rect 22320 16962 22800 16992
rect 11513 16960 13603 16962
rect 11513 16904 11518 16960
rect 11574 16904 13542 16960
rect 13598 16904 13603 16960
rect 11513 16902 13603 16904
rect 11513 16899 11579 16902
rect 13537 16899 13603 16902
rect 15104 16902 22800 16962
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 3918 16764 3924 16828
rect 3988 16826 3994 16828
rect 4061 16826 4127 16829
rect 3988 16824 4127 16826
rect 3988 16768 4066 16824
rect 4122 16768 4127 16824
rect 3988 16766 4127 16768
rect 3988 16764 3994 16766
rect 4061 16763 4127 16766
rect 9254 16764 9260 16828
rect 9324 16826 9330 16828
rect 9581 16826 9647 16829
rect 11881 16826 11947 16829
rect 9324 16824 9647 16826
rect 9324 16768 9586 16824
rect 9642 16768 9647 16824
rect 9324 16766 9647 16768
rect 9324 16764 9330 16766
rect 9581 16763 9647 16766
rect 11286 16824 11947 16826
rect 11286 16768 11886 16824
rect 11942 16768 11947 16824
rect 11286 16766 11947 16768
rect 3693 16690 3759 16693
rect 11286 16690 11346 16766
rect 11881 16763 11947 16766
rect 3693 16688 11346 16690
rect 3693 16632 3698 16688
rect 3754 16632 11346 16688
rect 3693 16630 11346 16632
rect 14273 16690 14339 16693
rect 15104 16690 15164 16902
rect 22320 16872 22800 16902
rect 14273 16688 15164 16690
rect 14273 16632 14278 16688
rect 14334 16632 15164 16688
rect 14273 16630 15164 16632
rect 3693 16627 3759 16630
rect 14273 16627 14339 16630
rect 0 16554 480 16584
rect 1945 16554 2011 16557
rect 0 16552 2011 16554
rect 0 16496 1950 16552
rect 2006 16496 2011 16552
rect 0 16494 2011 16496
rect 0 16464 480 16494
rect 1945 16491 2011 16494
rect 3918 16492 3924 16556
rect 3988 16554 3994 16556
rect 16297 16554 16363 16557
rect 3988 16552 16363 16554
rect 3988 16496 16302 16552
rect 16358 16496 16363 16552
rect 3988 16494 16363 16496
rect 3988 16492 3994 16494
rect 16297 16491 16363 16494
rect 18873 16554 18939 16557
rect 22320 16554 22800 16584
rect 18873 16552 22800 16554
rect 18873 16496 18878 16552
rect 18934 16496 22800 16552
rect 18873 16494 22800 16496
rect 18873 16491 18939 16494
rect 22320 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 2773 16146 2839 16149
rect 9213 16146 9279 16149
rect 2773 16144 9279 16146
rect 2773 16088 2778 16144
rect 2834 16088 9218 16144
rect 9274 16088 9279 16144
rect 2773 16086 9279 16088
rect 2773 16083 2839 16086
rect 9213 16083 9279 16086
rect 16297 16146 16363 16149
rect 19190 16146 19196 16148
rect 16297 16144 19196 16146
rect 16297 16088 16302 16144
rect 16358 16088 19196 16144
rect 16297 16086 19196 16088
rect 16297 16083 16363 16086
rect 19190 16084 19196 16086
rect 19260 16084 19266 16148
rect 0 16010 480 16040
rect 1945 16010 2011 16013
rect 0 16008 2011 16010
rect 0 15952 1950 16008
rect 2006 15952 2011 16008
rect 0 15950 2011 15952
rect 0 15920 480 15950
rect 1945 15947 2011 15950
rect 7189 16010 7255 16013
rect 7557 16010 7623 16013
rect 7189 16008 7623 16010
rect 7189 15952 7194 16008
rect 7250 15952 7562 16008
rect 7618 15952 7623 16008
rect 7189 15950 7623 15952
rect 7189 15947 7255 15950
rect 7557 15947 7623 15950
rect 19006 15948 19012 16012
rect 19076 16010 19082 16012
rect 22320 16010 22800 16040
rect 19076 15950 22800 16010
rect 19076 15948 19082 15950
rect 22320 15920 22800 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 7189 15738 7255 15741
rect 7189 15736 7482 15738
rect 7189 15680 7194 15736
rect 7250 15680 7482 15736
rect 7189 15678 7482 15680
rect 7189 15675 7255 15678
rect 0 15602 480 15632
rect 1945 15602 2011 15605
rect 0 15600 2011 15602
rect 0 15544 1950 15600
rect 2006 15544 2011 15600
rect 0 15542 2011 15544
rect 7422 15602 7482 15678
rect 8109 15602 8175 15605
rect 7422 15600 8175 15602
rect 7422 15544 8114 15600
rect 8170 15544 8175 15600
rect 7422 15542 8175 15544
rect 0 15512 480 15542
rect 1945 15539 2011 15542
rect 8109 15539 8175 15542
rect 15929 15602 15995 15605
rect 22320 15602 22800 15632
rect 15929 15600 22800 15602
rect 15929 15544 15934 15600
rect 15990 15544 22800 15600
rect 15929 15542 22800 15544
rect 15929 15539 15995 15542
rect 22320 15512 22800 15542
rect 6361 15466 6427 15469
rect 9673 15466 9739 15469
rect 6361 15464 9739 15466
rect 6361 15408 6366 15464
rect 6422 15408 9678 15464
rect 9734 15408 9739 15464
rect 6361 15406 9739 15408
rect 6361 15403 6427 15406
rect 9673 15403 9739 15406
rect 10409 15466 10475 15469
rect 13077 15466 13143 15469
rect 18638 15466 18644 15468
rect 10409 15464 18644 15466
rect 10409 15408 10414 15464
rect 10470 15408 13082 15464
rect 13138 15408 18644 15464
rect 10409 15406 18644 15408
rect 10409 15403 10475 15406
rect 13077 15403 13143 15406
rect 18638 15404 18644 15406
rect 18708 15404 18714 15468
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 480 15088
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14968 480 14998
rect 2773 14995 2839 14998
rect 17953 15058 18019 15061
rect 22320 15058 22800 15088
rect 17953 15056 22800 15058
rect 17953 15000 17958 15056
rect 18014 15000 22800 15056
rect 17953 14998 22800 15000
rect 17953 14995 18019 14998
rect 22320 14968 22800 14998
rect 16205 14922 16271 14925
rect 9676 14920 16271 14922
rect 9676 14864 16210 14920
rect 16266 14864 16271 14920
rect 9676 14862 16271 14864
rect 7808 14720 8128 14721
rect 0 14650 480 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 9676 14653 9736 14862
rect 16205 14859 16271 14862
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 3141 14650 3207 14653
rect 0 14648 3207 14650
rect 0 14592 3146 14648
rect 3202 14592 3207 14648
rect 0 14590 3207 14592
rect 0 14560 480 14590
rect 3141 14587 3207 14590
rect 9673 14648 9739 14653
rect 22320 14650 22800 14680
rect 9673 14592 9678 14648
rect 9734 14592 9739 14648
rect 9673 14587 9739 14592
rect 15104 14590 22800 14650
rect 10501 14514 10567 14517
rect 9630 14512 10567 14514
rect 9630 14456 10506 14512
rect 10562 14456 10567 14512
rect 9630 14454 10567 14456
rect 9630 14242 9690 14454
rect 10501 14451 10567 14454
rect 13077 14514 13143 14517
rect 15104 14514 15164 14590
rect 22320 14560 22800 14590
rect 13077 14512 15164 14514
rect 13077 14456 13082 14512
rect 13138 14456 15164 14512
rect 13077 14454 15164 14456
rect 13077 14451 13143 14454
rect 9765 14378 9831 14381
rect 10501 14378 10567 14381
rect 9765 14376 10567 14378
rect 9765 14320 9770 14376
rect 9826 14320 10506 14376
rect 10562 14320 10567 14376
rect 9765 14318 10567 14320
rect 9765 14315 9831 14318
rect 10501 14315 10567 14318
rect 16113 14378 16179 14381
rect 16941 14378 17007 14381
rect 17769 14378 17835 14381
rect 16113 14376 17835 14378
rect 16113 14320 16118 14376
rect 16174 14320 16946 14376
rect 17002 14320 17774 14376
rect 17830 14320 17835 14376
rect 16113 14318 17835 14320
rect 16113 14315 16179 14318
rect 16941 14315 17007 14318
rect 17769 14315 17835 14318
rect 9765 14242 9831 14245
rect 9630 14240 9831 14242
rect 9630 14184 9770 14240
rect 9826 14184 9831 14240
rect 9630 14182 9831 14184
rect 9765 14179 9831 14182
rect 4376 14176 4696 14177
rect 0 14106 480 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1761 14106 1827 14109
rect 0 14104 1827 14106
rect 0 14048 1766 14104
rect 1822 14048 1827 14104
rect 0 14046 1827 14048
rect 0 14016 480 14046
rect 1761 14043 1827 14046
rect 5993 14106 6059 14109
rect 20989 14106 21055 14109
rect 22320 14106 22800 14136
rect 5993 14104 10058 14106
rect 5993 14048 5998 14104
rect 6054 14048 10058 14104
rect 5993 14046 10058 14048
rect 5993 14043 6059 14046
rect 9998 13834 10058 14046
rect 20989 14104 22800 14106
rect 20989 14048 20994 14104
rect 21050 14048 22800 14104
rect 20989 14046 22800 14048
rect 20989 14043 21055 14046
rect 22320 14016 22800 14046
rect 17902 13908 17908 13972
rect 17972 13970 17978 13972
rect 18229 13970 18295 13973
rect 17972 13968 18295 13970
rect 17972 13912 18234 13968
rect 18290 13912 18295 13968
rect 17972 13910 18295 13912
rect 17972 13908 17978 13910
rect 18229 13907 18295 13910
rect 10133 13834 10199 13837
rect 19057 13834 19123 13837
rect 9998 13832 19123 13834
rect 9998 13776 10138 13832
rect 10194 13776 19062 13832
rect 19118 13776 19123 13832
rect 9998 13774 19123 13776
rect 10133 13771 10199 13774
rect 19057 13771 19123 13774
rect 0 13698 480 13728
rect 3141 13698 3207 13701
rect 0 13696 3207 13698
rect 0 13640 3146 13696
rect 3202 13640 3207 13696
rect 0 13638 3207 13640
rect 0 13608 480 13638
rect 3141 13635 3207 13638
rect 15193 13698 15259 13701
rect 18229 13698 18295 13701
rect 15193 13696 18295 13698
rect 15193 13640 15198 13696
rect 15254 13640 18234 13696
rect 18290 13640 18295 13696
rect 15193 13638 18295 13640
rect 15193 13635 15259 13638
rect 18229 13635 18295 13638
rect 18781 13698 18847 13701
rect 22320 13698 22800 13728
rect 18781 13696 22800 13698
rect 18781 13640 18786 13696
rect 18842 13640 22800 13696
rect 18781 13638 22800 13640
rect 18781 13635 18847 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22320 13608 22800 13638
rect 14672 13567 14992 13568
rect 16021 13562 16087 13565
rect 16573 13562 16639 13565
rect 16021 13560 16639 13562
rect 16021 13504 16026 13560
rect 16082 13504 16578 13560
rect 16634 13504 16639 13560
rect 16021 13502 16639 13504
rect 16021 13499 16087 13502
rect 16573 13499 16639 13502
rect 8334 13364 8340 13428
rect 8404 13426 8410 13428
rect 9305 13426 9371 13429
rect 8404 13424 9371 13426
rect 8404 13368 9310 13424
rect 9366 13368 9371 13424
rect 8404 13366 9371 13368
rect 8404 13364 8410 13366
rect 9305 13363 9371 13366
rect 16389 13426 16455 13429
rect 19977 13426 20043 13429
rect 16389 13424 20043 13426
rect 16389 13368 16394 13424
rect 16450 13368 19982 13424
rect 20038 13368 20043 13424
rect 16389 13366 20043 13368
rect 16389 13363 16455 13366
rect 19977 13363 20043 13366
rect 0 13290 480 13320
rect 2313 13290 2379 13293
rect 0 13288 2379 13290
rect 0 13232 2318 13288
rect 2374 13232 2379 13288
rect 0 13230 2379 13232
rect 0 13200 480 13230
rect 2313 13227 2379 13230
rect 11329 13290 11395 13293
rect 20161 13290 20227 13293
rect 22320 13290 22800 13320
rect 11329 13288 13554 13290
rect 11329 13232 11334 13288
rect 11390 13232 13554 13288
rect 11329 13230 13554 13232
rect 11329 13227 11395 13230
rect 13494 13154 13554 13230
rect 20161 13288 22800 13290
rect 20161 13232 20166 13288
rect 20222 13232 22800 13288
rect 20161 13230 22800 13232
rect 20161 13227 20227 13230
rect 22320 13200 22800 13230
rect 17493 13154 17559 13157
rect 13494 13152 17559 13154
rect 13494 13096 17498 13152
rect 17554 13096 17559 13152
rect 13494 13094 17559 13096
rect 17493 13091 17559 13094
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 12249 13018 12315 13021
rect 12249 13016 16636 13018
rect 12249 12960 12254 13016
rect 12310 12960 16636 13016
rect 12249 12958 16636 12960
rect 12249 12955 12315 12958
rect 3693 12882 3759 12885
rect 15469 12882 15535 12885
rect 3693 12880 15535 12882
rect 3693 12824 3698 12880
rect 3754 12824 15474 12880
rect 15530 12824 15535 12880
rect 3693 12822 15535 12824
rect 3693 12819 3759 12822
rect 15469 12819 15535 12822
rect 0 12746 480 12776
rect 3509 12746 3575 12749
rect 0 12744 3575 12746
rect 0 12688 3514 12744
rect 3570 12688 3575 12744
rect 0 12686 3575 12688
rect 0 12656 480 12686
rect 3509 12683 3575 12686
rect 13169 12746 13235 12749
rect 16389 12746 16455 12749
rect 13169 12744 16455 12746
rect 13169 12688 13174 12744
rect 13230 12688 16394 12744
rect 16450 12688 16455 12744
rect 13169 12686 16455 12688
rect 16576 12746 16636 12958
rect 18965 12884 19031 12885
rect 18965 12882 19012 12884
rect 18920 12880 19012 12882
rect 18920 12824 18970 12880
rect 18920 12822 19012 12824
rect 18965 12820 19012 12822
rect 19076 12820 19082 12884
rect 18965 12819 19031 12820
rect 18822 12746 18828 12748
rect 16576 12686 18828 12746
rect 13169 12683 13235 12686
rect 16389 12683 16455 12686
rect 18822 12684 18828 12686
rect 18892 12746 18898 12748
rect 22320 12746 22800 12776
rect 18892 12686 22800 12746
rect 18892 12684 18898 12686
rect 22320 12656 22800 12686
rect 3509 12610 3575 12613
rect 3918 12610 3924 12612
rect 3509 12608 3924 12610
rect 3509 12552 3514 12608
rect 3570 12552 3924 12608
rect 3509 12550 3924 12552
rect 3509 12547 3575 12550
rect 3918 12548 3924 12550
rect 3988 12548 3994 12612
rect 16205 12610 16271 12613
rect 19006 12610 19012 12612
rect 16205 12608 19012 12610
rect 16205 12552 16210 12608
rect 16266 12552 19012 12608
rect 16205 12550 19012 12552
rect 16205 12547 16271 12550
rect 19006 12548 19012 12550
rect 19076 12548 19082 12612
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 480 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 480 12278
rect 4061 12275 4127 12278
rect 13813 12338 13879 12341
rect 17493 12338 17559 12341
rect 13813 12336 17559 12338
rect 13813 12280 13818 12336
rect 13874 12280 17498 12336
rect 17554 12280 17559 12336
rect 13813 12278 17559 12280
rect 13813 12275 13879 12278
rect 17493 12275 17559 12278
rect 17677 12338 17743 12341
rect 22320 12338 22800 12368
rect 17677 12336 22800 12338
rect 17677 12280 17682 12336
rect 17738 12280 22800 12336
rect 17677 12278 22800 12280
rect 17677 12275 17743 12278
rect 22320 12248 22800 12278
rect 12433 12202 12499 12205
rect 15745 12202 15811 12205
rect 12433 12200 15811 12202
rect 12433 12144 12438 12200
rect 12494 12144 15750 12200
rect 15806 12144 15811 12200
rect 12433 12142 15811 12144
rect 12433 12139 12499 12142
rect 15745 12139 15811 12142
rect 11973 12066 12039 12069
rect 11838 12064 12039 12066
rect 11838 12008 11978 12064
rect 12034 12008 12039 12064
rect 11838 12006 12039 12008
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 0 11794 480 11824
rect 4061 11794 4127 11797
rect 0 11792 4127 11794
rect 0 11736 4066 11792
rect 4122 11736 4127 11792
rect 0 11734 4127 11736
rect 0 11704 480 11734
rect 4061 11731 4127 11734
rect 10777 11658 10843 11661
rect 11053 11658 11119 11661
rect 11329 11658 11395 11661
rect 10777 11656 11395 11658
rect 10777 11600 10782 11656
rect 10838 11600 11058 11656
rect 11114 11600 11334 11656
rect 11390 11600 11395 11656
rect 10777 11598 11395 11600
rect 10777 11595 10843 11598
rect 11053 11595 11119 11598
rect 11329 11595 11395 11598
rect 11838 11525 11898 12006
rect 11973 12003 12039 12006
rect 12341 12066 12407 12069
rect 15377 12066 15443 12069
rect 12341 12064 15443 12066
rect 12341 12008 12346 12064
rect 12402 12008 15382 12064
rect 15438 12008 15443 12064
rect 12341 12006 15443 12008
rect 12341 12003 12407 12006
rect 15377 12003 15443 12006
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 19190 11732 19196 11796
rect 19260 11794 19266 11796
rect 22320 11794 22800 11824
rect 19260 11734 22800 11794
rect 19260 11732 19266 11734
rect 22320 11704 22800 11734
rect 18413 11658 18479 11661
rect 11789 11520 11898 11525
rect 11789 11464 11794 11520
rect 11850 11464 11898 11520
rect 11789 11462 11898 11464
rect 14552 11656 18479 11658
rect 14552 11600 18418 11656
rect 18474 11600 18479 11656
rect 14552 11598 18479 11600
rect 11789 11459 11855 11462
rect 7808 11456 8128 11457
rect 0 11386 480 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 3601 11386 3667 11389
rect 0 11384 3667 11386
rect 0 11328 3606 11384
rect 3662 11328 3667 11384
rect 0 11326 3667 11328
rect 0 11296 480 11326
rect 3601 11323 3667 11326
rect 10133 11386 10199 11389
rect 14552 11386 14612 11598
rect 18413 11595 18479 11598
rect 15469 11522 15535 11525
rect 19241 11522 19307 11525
rect 15469 11520 19307 11522
rect 15469 11464 15474 11520
rect 15530 11464 19246 11520
rect 19302 11464 19307 11520
rect 15469 11462 19307 11464
rect 15469 11459 15535 11462
rect 19241 11459 19307 11462
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 10133 11384 14612 11386
rect 10133 11328 10138 11384
rect 10194 11328 14612 11384
rect 10133 11326 14612 11328
rect 17861 11386 17927 11389
rect 22320 11386 22800 11416
rect 17861 11384 22800 11386
rect 17861 11328 17866 11384
rect 17922 11328 22800 11384
rect 17861 11326 22800 11328
rect 10133 11323 10199 11326
rect 17861 11323 17927 11326
rect 22320 11296 22800 11326
rect 11605 11250 11671 11253
rect 11102 11248 11671 11250
rect 11102 11192 11610 11248
rect 11666 11192 11671 11248
rect 11102 11190 11671 11192
rect 10961 11114 11027 11117
rect 11102 11114 11162 11190
rect 11605 11187 11671 11190
rect 10961 11112 11162 11114
rect 10961 11056 10966 11112
rect 11022 11056 11162 11112
rect 10961 11054 11162 11056
rect 11421 11114 11487 11117
rect 12801 11114 12867 11117
rect 13537 11114 13603 11117
rect 11421 11112 11898 11114
rect 11421 11056 11426 11112
rect 11482 11056 11898 11112
rect 11421 11054 11898 11056
rect 10961 11051 11027 11054
rect 11421 11051 11487 11054
rect 9438 10978 9444 10980
rect 7008 10918 9444 10978
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 3969 10842 4035 10845
rect 0 10840 4035 10842
rect 0 10784 3974 10840
rect 4030 10784 4035 10840
rect 0 10782 4035 10784
rect 0 10752 480 10782
rect 3969 10779 4035 10782
rect 4838 10508 4844 10572
rect 4908 10570 4914 10572
rect 6361 10570 6427 10573
rect 4908 10568 6427 10570
rect 4908 10512 6366 10568
rect 6422 10512 6427 10568
rect 4908 10510 6427 10512
rect 4908 10508 4914 10510
rect 6361 10507 6427 10510
rect 0 10434 480 10464
rect 7008 10434 7068 10918
rect 9438 10916 9444 10918
rect 9508 10978 9514 10980
rect 10685 10978 10751 10981
rect 9508 10976 10751 10978
rect 9508 10920 10690 10976
rect 10746 10920 10751 10976
rect 9508 10918 10751 10920
rect 11838 10978 11898 11054
rect 12801 11112 13603 11114
rect 12801 11056 12806 11112
rect 12862 11056 13542 11112
rect 13598 11056 13603 11112
rect 12801 11054 13603 11056
rect 12801 11051 12867 11054
rect 13537 11051 13603 11054
rect 11973 10978 12039 10981
rect 11838 10976 12039 10978
rect 11838 10920 11978 10976
rect 12034 10920 12039 10976
rect 11838 10918 12039 10920
rect 9508 10916 9514 10918
rect 10685 10915 10751 10918
rect 11973 10915 12039 10918
rect 12617 10978 12683 10981
rect 13486 10978 13492 10980
rect 12617 10976 13492 10978
rect 12617 10920 12622 10976
rect 12678 10920 13492 10976
rect 12617 10918 13492 10920
rect 12617 10915 12683 10918
rect 13486 10916 13492 10918
rect 13556 10978 13562 10980
rect 17861 10978 17927 10981
rect 13556 10976 17927 10978
rect 13556 10920 17866 10976
rect 17922 10920 17927 10976
rect 13556 10918 17927 10920
rect 13556 10916 13562 10918
rect 17861 10915 17927 10918
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 18638 10780 18644 10844
rect 18708 10842 18714 10844
rect 22320 10842 22800 10872
rect 18708 10782 22800 10842
rect 18708 10780 18714 10782
rect 22320 10752 22800 10782
rect 10317 10706 10383 10709
rect 11697 10706 11763 10709
rect 16205 10706 16271 10709
rect 18873 10708 18939 10709
rect 18822 10706 18828 10708
rect 10317 10704 16271 10706
rect 10317 10648 10322 10704
rect 10378 10648 11702 10704
rect 11758 10648 16210 10704
rect 16266 10648 16271 10704
rect 10317 10646 16271 10648
rect 18782 10646 18828 10706
rect 18892 10704 18939 10708
rect 18934 10648 18939 10704
rect 10317 10643 10383 10646
rect 11697 10643 11763 10646
rect 16205 10643 16271 10646
rect 18822 10644 18828 10646
rect 18892 10644 18939 10648
rect 18873 10643 18939 10644
rect 11237 10570 11303 10573
rect 11789 10570 11855 10573
rect 20621 10570 20687 10573
rect 11237 10568 20687 10570
rect 11237 10512 11242 10568
rect 11298 10512 11794 10568
rect 11850 10512 20626 10568
rect 20682 10512 20687 10568
rect 11237 10510 20687 10512
rect 11237 10507 11303 10510
rect 11789 10507 11855 10510
rect 20621 10507 20687 10510
rect 22320 10434 22800 10464
rect 0 10374 7068 10434
rect 17358 10374 22800 10434
rect 0 10344 480 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 11513 10298 11579 10301
rect 12433 10298 12499 10301
rect 11513 10296 12499 10298
rect 11513 10240 11518 10296
rect 11574 10240 12438 10296
rect 12494 10240 12499 10296
rect 11513 10238 12499 10240
rect 11513 10235 11579 10238
rect 12433 10235 12499 10238
rect 6545 10162 6611 10165
rect 17358 10162 17418 10374
rect 22320 10344 22800 10374
rect 18413 10298 18479 10301
rect 18965 10298 19031 10301
rect 18413 10296 19031 10298
rect 18413 10240 18418 10296
rect 18474 10240 18970 10296
rect 19026 10240 19031 10296
rect 18413 10238 19031 10240
rect 18413 10235 18479 10238
rect 18965 10235 19031 10238
rect 6545 10160 17418 10162
rect 6545 10104 6550 10160
rect 6606 10104 17418 10160
rect 6545 10102 17418 10104
rect 17677 10162 17743 10165
rect 19517 10162 19583 10165
rect 17677 10160 19583 10162
rect 17677 10104 17682 10160
rect 17738 10104 19522 10160
rect 19578 10104 19583 10160
rect 17677 10102 19583 10104
rect 6545 10099 6611 10102
rect 17677 10099 17743 10102
rect 19517 10099 19583 10102
rect 0 10026 480 10056
rect 8661 10026 8727 10029
rect 0 10024 8727 10026
rect 0 9968 8666 10024
rect 8722 9968 8727 10024
rect 0 9966 8727 9968
rect 0 9936 480 9966
rect 8661 9963 8727 9966
rect 11145 10026 11211 10029
rect 11881 10026 11947 10029
rect 22320 10026 22800 10056
rect 11145 10024 22800 10026
rect 11145 9968 11150 10024
rect 11206 9968 11886 10024
rect 11942 9968 22800 10024
rect 11145 9966 22800 9968
rect 11145 9963 11211 9966
rect 11881 9963 11947 9966
rect 22320 9936 22800 9966
rect 18822 9828 18828 9892
rect 18892 9890 18898 9892
rect 18965 9890 19031 9893
rect 18892 9888 19031 9890
rect 18892 9832 18970 9888
rect 19026 9832 19031 9888
rect 18892 9830 19031 9832
rect 18892 9828 18898 9830
rect 18965 9827 19031 9830
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 11789 9754 11855 9757
rect 16665 9754 16731 9757
rect 11789 9752 16731 9754
rect 11789 9696 11794 9752
rect 11850 9696 16670 9752
rect 16726 9696 16731 9752
rect 11789 9694 16731 9696
rect 11789 9691 11855 9694
rect 16665 9691 16731 9694
rect 18873 9754 18939 9757
rect 19006 9754 19012 9756
rect 18873 9752 19012 9754
rect 18873 9696 18878 9752
rect 18934 9696 19012 9752
rect 18873 9694 19012 9696
rect 18873 9691 18939 9694
rect 19006 9692 19012 9694
rect 19076 9692 19082 9756
rect 14549 9618 14615 9621
rect 16297 9618 16363 9621
rect 14549 9616 16363 9618
rect 14549 9560 14554 9616
rect 14610 9560 16302 9616
rect 16358 9560 16363 9616
rect 14549 9558 16363 9560
rect 14549 9555 14615 9558
rect 16297 9555 16363 9558
rect 0 9482 480 9512
rect 3877 9482 3943 9485
rect 0 9480 3943 9482
rect 0 9424 3882 9480
rect 3938 9424 3943 9480
rect 0 9422 3943 9424
rect 0 9392 480 9422
rect 3877 9419 3943 9422
rect 11513 9482 11579 9485
rect 14089 9482 14155 9485
rect 11513 9480 14155 9482
rect 11513 9424 11518 9480
rect 11574 9424 14094 9480
rect 14150 9424 14155 9480
rect 11513 9422 14155 9424
rect 11513 9419 11579 9422
rect 14089 9419 14155 9422
rect 19149 9482 19215 9485
rect 22320 9482 22800 9512
rect 19149 9480 22800 9482
rect 19149 9424 19154 9480
rect 19210 9424 22800 9480
rect 19149 9422 22800 9424
rect 19149 9419 19215 9422
rect 22320 9392 22800 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9074 480 9104
rect 4061 9074 4127 9077
rect 0 9072 4127 9074
rect 0 9016 4066 9072
rect 4122 9016 4127 9072
rect 0 9014 4127 9016
rect 0 8984 480 9014
rect 4061 9011 4127 9014
rect 4705 9074 4771 9077
rect 5165 9074 5231 9077
rect 5349 9074 5415 9077
rect 4705 9072 5415 9074
rect 4705 9016 4710 9072
rect 4766 9016 5170 9072
rect 5226 9016 5354 9072
rect 5410 9016 5415 9072
rect 4705 9014 5415 9016
rect 4705 9011 4771 9014
rect 5165 9011 5231 9014
rect 5349 9011 5415 9014
rect 17953 9074 18019 9077
rect 22320 9074 22800 9104
rect 17953 9072 22800 9074
rect 17953 9016 17958 9072
rect 18014 9016 22800 9072
rect 17953 9014 22800 9016
rect 17953 9011 18019 9014
rect 22320 8984 22800 9014
rect 4797 8938 4863 8941
rect 7281 8938 7347 8941
rect 4797 8936 7347 8938
rect 4797 8880 4802 8936
rect 4858 8880 7286 8936
rect 7342 8880 7347 8936
rect 4797 8878 7347 8880
rect 4797 8875 4863 8878
rect 7281 8875 7347 8878
rect 7925 8938 7991 8941
rect 9121 8938 9187 8941
rect 7925 8936 9187 8938
rect 7925 8880 7930 8936
rect 7986 8880 9126 8936
rect 9182 8880 9187 8936
rect 7925 8878 9187 8880
rect 7925 8875 7991 8878
rect 9121 8875 9187 8878
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 0 8530 480 8560
rect 4061 8530 4127 8533
rect 0 8528 4127 8530
rect 0 8472 4066 8528
rect 4122 8472 4127 8528
rect 0 8470 4127 8472
rect 0 8440 480 8470
rect 4061 8467 4127 8470
rect 4797 8530 4863 8533
rect 5533 8530 5599 8533
rect 4797 8528 5599 8530
rect 4797 8472 4802 8528
rect 4858 8472 5538 8528
rect 5594 8472 5599 8528
rect 4797 8470 5599 8472
rect 4797 8467 4863 8470
rect 5533 8467 5599 8470
rect 12433 8530 12499 8533
rect 13445 8530 13511 8533
rect 12433 8528 13511 8530
rect 12433 8472 12438 8528
rect 12494 8472 13450 8528
rect 13506 8472 13511 8528
rect 12433 8470 13511 8472
rect 12433 8467 12499 8470
rect 13445 8467 13511 8470
rect 21081 8530 21147 8533
rect 22320 8530 22800 8560
rect 21081 8528 22800 8530
rect 21081 8472 21086 8528
rect 21142 8472 22800 8528
rect 21081 8470 22800 8472
rect 21081 8467 21147 8470
rect 22320 8440 22800 8470
rect 7808 8192 8128 8193
rect 0 8122 480 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 5073 8122 5139 8125
rect 6453 8122 6519 8125
rect 0 8062 4906 8122
rect 0 8032 480 8062
rect 4846 7986 4906 8062
rect 5073 8120 6519 8122
rect 5073 8064 5078 8120
rect 5134 8064 6458 8120
rect 6514 8064 6519 8120
rect 5073 8062 6519 8064
rect 5073 8059 5139 8062
rect 6453 8059 6519 8062
rect 18873 8122 18939 8125
rect 22320 8122 22800 8152
rect 18873 8120 22800 8122
rect 18873 8064 18878 8120
rect 18934 8064 22800 8120
rect 18873 8062 22800 8064
rect 18873 8059 18939 8062
rect 22320 8032 22800 8062
rect 5349 7986 5415 7989
rect 4846 7984 5415 7986
rect 4846 7928 5354 7984
rect 5410 7928 5415 7984
rect 4846 7926 5415 7928
rect 5349 7923 5415 7926
rect 14365 7850 14431 7853
rect 14365 7848 18706 7850
rect 14365 7792 14370 7848
rect 14426 7792 18706 7848
rect 14365 7790 18706 7792
rect 14365 7787 14431 7790
rect 4376 7648 4696 7649
rect 0 7578 480 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 2865 7578 2931 7581
rect 0 7576 2931 7578
rect 0 7520 2870 7576
rect 2926 7520 2931 7576
rect 0 7518 2931 7520
rect 18646 7578 18706 7790
rect 22320 7578 22800 7608
rect 18646 7518 22800 7578
rect 0 7488 480 7518
rect 2865 7515 2931 7518
rect 22320 7488 22800 7518
rect 0 7170 480 7200
rect 3509 7170 3575 7173
rect 0 7168 3575 7170
rect 0 7112 3514 7168
rect 3570 7112 3575 7168
rect 0 7110 3575 7112
rect 0 7080 480 7110
rect 3509 7107 3575 7110
rect 19241 7170 19307 7173
rect 22320 7170 22800 7200
rect 19241 7168 22800 7170
rect 19241 7112 19246 7168
rect 19302 7112 22800 7168
rect 19241 7110 22800 7112
rect 19241 7107 19307 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 22320 7080 22800 7110
rect 14672 7039 14992 7040
rect 0 6762 480 6792
rect 4061 6762 4127 6765
rect 0 6760 4127 6762
rect 0 6704 4066 6760
rect 4122 6704 4127 6760
rect 0 6702 4127 6704
rect 0 6672 480 6702
rect 4061 6699 4127 6702
rect 18781 6762 18847 6765
rect 22320 6762 22800 6792
rect 18781 6760 22800 6762
rect 18781 6704 18786 6760
rect 18842 6704 22800 6760
rect 18781 6702 22800 6704
rect 18781 6699 18847 6702
rect 22320 6672 22800 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 0 6218 480 6248
rect 3969 6218 4035 6221
rect 0 6216 4035 6218
rect 0 6160 3974 6216
rect 4030 6160 4035 6216
rect 0 6158 4035 6160
rect 0 6128 480 6158
rect 3969 6155 4035 6158
rect 10133 6218 10199 6221
rect 22320 6218 22800 6248
rect 10133 6216 22800 6218
rect 10133 6160 10138 6216
rect 10194 6160 22800 6216
rect 10133 6158 22800 6160
rect 10133 6155 10199 6158
rect 22320 6128 22800 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 3417 5810 3483 5813
rect 0 5808 3483 5810
rect 0 5752 3422 5808
rect 3478 5752 3483 5808
rect 0 5750 3483 5752
rect 0 5720 480 5750
rect 3417 5747 3483 5750
rect 17953 5810 18019 5813
rect 22320 5810 22800 5840
rect 17953 5808 22800 5810
rect 17953 5752 17958 5808
rect 18014 5752 22800 5808
rect 17953 5750 22800 5752
rect 17953 5747 18019 5750
rect 22320 5720 22800 5750
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 480 5296
rect 4061 5266 4127 5269
rect 0 5264 4127 5266
rect 0 5208 4066 5264
rect 4122 5208 4127 5264
rect 0 5206 4127 5208
rect 0 5176 480 5206
rect 4061 5203 4127 5206
rect 11605 5266 11671 5269
rect 22320 5266 22800 5296
rect 11605 5264 22800 5266
rect 11605 5208 11610 5264
rect 11666 5208 22800 5264
rect 11605 5206 22800 5208
rect 11605 5203 11671 5206
rect 22320 5176 22800 5206
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 4061 4858 4127 4861
rect 0 4856 4127 4858
rect 0 4800 4066 4856
rect 4122 4800 4127 4856
rect 0 4798 4127 4800
rect 0 4768 480 4798
rect 4061 4795 4127 4798
rect 17953 4858 18019 4861
rect 22320 4858 22800 4888
rect 17953 4856 22800 4858
rect 17953 4800 17958 4856
rect 18014 4800 22800 4856
rect 17953 4798 22800 4800
rect 17953 4795 18019 4798
rect 22320 4768 22800 4798
rect 4376 4384 4696 4385
rect 0 4314 480 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 2865 4314 2931 4317
rect 0 4312 2931 4314
rect 0 4256 2870 4312
rect 2926 4256 2931 4312
rect 0 4254 2931 4256
rect 0 4224 480 4254
rect 2865 4251 2931 4254
rect 20529 4314 20595 4317
rect 22320 4314 22800 4344
rect 20529 4312 22800 4314
rect 20529 4256 20534 4312
rect 20590 4256 22800 4312
rect 20529 4254 22800 4256
rect 20529 4251 20595 4254
rect 22320 4224 22800 4254
rect 0 3906 480 3936
rect 4153 3906 4219 3909
rect 0 3904 4219 3906
rect 0 3848 4158 3904
rect 4214 3848 4219 3904
rect 0 3846 4219 3848
rect 0 3816 480 3846
rect 4153 3843 4219 3846
rect 20437 3906 20503 3909
rect 22320 3906 22800 3936
rect 20437 3904 22800 3906
rect 20437 3848 20442 3904
rect 20498 3848 22800 3904
rect 20437 3846 22800 3848
rect 20437 3843 20503 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22320 3816 22800 3846
rect 14672 3775 14992 3776
rect 0 3498 480 3528
rect 3325 3498 3391 3501
rect 0 3496 3391 3498
rect 0 3440 3330 3496
rect 3386 3440 3391 3496
rect 0 3438 3391 3440
rect 0 3408 480 3438
rect 3325 3435 3391 3438
rect 20621 3498 20687 3501
rect 22320 3498 22800 3528
rect 20621 3496 22800 3498
rect 20621 3440 20626 3496
rect 20682 3440 22800 3496
rect 20621 3438 22800 3440
rect 20621 3435 20687 3438
rect 22320 3408 22800 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 0 2954 480 2984
rect 4797 2954 4863 2957
rect 0 2952 4863 2954
rect 0 2896 4802 2952
rect 4858 2896 4863 2952
rect 0 2894 4863 2896
rect 0 2864 480 2894
rect 4797 2891 4863 2894
rect 20069 2954 20135 2957
rect 22320 2954 22800 2984
rect 20069 2952 22800 2954
rect 20069 2896 20074 2952
rect 20130 2896 22800 2952
rect 20069 2894 22800 2896
rect 20069 2891 20135 2894
rect 22320 2864 22800 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 480 2576
rect 1853 2546 1919 2549
rect 0 2544 1919 2546
rect 0 2488 1858 2544
rect 1914 2488 1919 2544
rect 0 2486 1919 2488
rect 0 2456 480 2486
rect 1853 2483 1919 2486
rect 17585 2546 17651 2549
rect 22320 2546 22800 2576
rect 17585 2544 22800 2546
rect 17585 2488 17590 2544
rect 17646 2488 22800 2544
rect 17585 2486 22800 2488
rect 17585 2483 17651 2486
rect 22320 2456 22800 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 480 2032
rect 4245 2002 4311 2005
rect 0 2000 4311 2002
rect 0 1944 4250 2000
rect 4306 1944 4311 2000
rect 0 1942 4311 1944
rect 0 1912 480 1942
rect 4245 1939 4311 1942
rect 21357 2002 21423 2005
rect 22320 2002 22800 2032
rect 21357 2000 22800 2002
rect 21357 1944 21362 2000
rect 21418 1944 22800 2000
rect 21357 1942 22800 1944
rect 21357 1939 21423 1942
rect 22320 1912 22800 1942
rect 0 1594 480 1624
rect 2773 1594 2839 1597
rect 0 1592 2839 1594
rect 0 1536 2778 1592
rect 2834 1536 2839 1592
rect 0 1534 2839 1536
rect 0 1504 480 1534
rect 2773 1531 2839 1534
rect 17769 1594 17835 1597
rect 22320 1594 22800 1624
rect 17769 1592 22800 1594
rect 17769 1536 17774 1592
rect 17830 1536 22800 1592
rect 17769 1534 22800 1536
rect 17769 1531 17835 1534
rect 22320 1504 22800 1534
rect 0 1050 480 1080
rect 6545 1050 6611 1053
rect 0 1048 6611 1050
rect 0 992 6550 1048
rect 6606 992 6611 1048
rect 0 990 6611 992
rect 0 960 480 990
rect 6545 987 6611 990
rect 18873 1050 18939 1053
rect 22320 1050 22800 1080
rect 18873 1048 22800 1050
rect 18873 992 18878 1048
rect 18934 992 22800 1048
rect 18873 990 22800 992
rect 18873 987 18939 990
rect 22320 960 22800 990
rect 0 642 480 672
rect 2773 642 2839 645
rect 0 640 2839 642
rect 0 584 2778 640
rect 2834 584 2839 640
rect 0 582 2839 584
rect 0 552 480 582
rect 2773 579 2839 582
rect 18689 642 18755 645
rect 22320 642 22800 672
rect 18689 640 22800 642
rect 18689 584 18694 640
rect 18750 584 22800 640
rect 18689 582 22800 584
rect 18689 579 18755 582
rect 22320 552 22800 582
rect 0 234 480 264
rect 7557 234 7623 237
rect 0 232 7623 234
rect 0 176 7562 232
rect 7618 176 7623 232
rect 0 174 7623 176
rect 0 144 480 174
rect 7557 171 7623 174
rect 19057 234 19123 237
rect 22320 234 22800 264
rect 19057 232 22800 234
rect 19057 176 19062 232
rect 19118 176 22800 232
rect 19057 174 22800 176
rect 19057 171 19123 174
rect 22320 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 4844 18456 4908 18460
rect 4844 18400 4858 18456
rect 4858 18400 4908 18456
rect 4844 18396 4908 18400
rect 8340 18396 8404 18460
rect 17908 18260 17972 18324
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 9444 17716 9508 17780
rect 13492 18048 13556 18052
rect 13492 17992 13542 18048
rect 13542 17992 13556 18048
rect 13492 17988 13556 17992
rect 18828 18048 18892 18052
rect 18828 17992 18878 18048
rect 18878 17992 18892 18048
rect 18828 17988 18892 17992
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 9260 17580 9324 17644
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 3924 16764 3988 16828
rect 9260 16764 9324 16828
rect 3924 16492 3988 16556
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 19196 16084 19260 16148
rect 19012 15948 19076 16012
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 18644 15404 18708 15468
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 17908 13908 17972 13972
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 8340 13364 8404 13428
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 19012 12880 19076 12884
rect 19012 12824 19026 12880
rect 19026 12824 19076 12880
rect 19012 12820 19076 12824
rect 18828 12684 18892 12748
rect 3924 12548 3988 12612
rect 19012 12548 19076 12612
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 19196 11732 19260 11796
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 4844 10508 4908 10572
rect 9444 10916 9508 10980
rect 13492 10916 13556 10980
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 18644 10780 18708 10844
rect 18828 10704 18892 10708
rect 18828 10648 18878 10704
rect 18878 10648 18892 10704
rect 18828 10644 18892 10648
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 18828 9828 18892 9892
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 19012 9692 19076 9756
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 4843 18460 4909 18461
rect 4843 18396 4844 18460
rect 4908 18396 4909 18460
rect 4843 18395 4909 18396
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 3923 16828 3989 16829
rect 3923 16764 3924 16828
rect 3988 16764 3989 16828
rect 3923 16763 3989 16764
rect 3926 16557 3986 16763
rect 3923 16556 3989 16557
rect 3923 16492 3924 16556
rect 3988 16492 3989 16556
rect 3923 16491 3989 16492
rect 3926 12613 3986 16491
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 3923 12612 3989 12613
rect 3923 12548 3924 12612
rect 3988 12548 3989 12612
rect 3923 12547 3989 12548
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4846 10573 4906 18395
rect 7808 17984 8128 19008
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 8339 18460 8405 18461
rect 8339 18396 8340 18460
rect 8404 18396 8405 18460
rect 8339 18395 8405 18396
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 8342 13429 8402 18395
rect 9443 17780 9509 17781
rect 9443 17716 9444 17780
rect 9508 17716 9509 17780
rect 9443 17715 9509 17716
rect 9259 17644 9325 17645
rect 9259 17580 9260 17644
rect 9324 17580 9325 17644
rect 9259 17579 9325 17580
rect 9262 16829 9322 17579
rect 9259 16828 9325 16829
rect 9259 16764 9260 16828
rect 9324 16764 9325 16828
rect 9259 16763 9325 16764
rect 8339 13428 8405 13429
rect 8339 13364 8340 13428
rect 8404 13364 8405 13428
rect 8339 13363 8405 13364
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 4843 10572 4909 10573
rect 4843 10508 4844 10572
rect 4908 10508 4909 10572
rect 4843 10507 4909 10508
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 10368 8128 11392
rect 9446 10981 9506 17715
rect 11240 17440 11560 18464
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 13491 18052 13557 18053
rect 13491 17988 13492 18052
rect 13556 17988 13557 18052
rect 13491 17987 13557 17988
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 9443 10980 9509 10981
rect 9443 10916 9444 10980
rect 9508 10916 9509 10980
rect 9443 10915 9509 10916
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 10912 11560 11936
rect 13494 10981 13554 17987
rect 14672 17984 14992 19008
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 17907 18324 17973 18325
rect 17907 18260 17908 18324
rect 17972 18260 17973 18324
rect 17907 18259 17973 18260
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 17910 13973 17970 18259
rect 18104 17440 18424 18464
rect 18827 18052 18893 18053
rect 18827 17988 18828 18052
rect 18892 17988 18893 18052
rect 18827 17987 18893 17988
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18643 15468 18709 15469
rect 18643 15404 18644 15468
rect 18708 15404 18709 15468
rect 18643 15403 18709 15404
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 17907 13972 17973 13973
rect 17907 13908 17908 13972
rect 17972 13908 17973 13972
rect 17907 13907 17973 13908
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 13491 10980 13557 10981
rect 13491 10916 13492 10980
rect 13556 10916 13557 10980
rect 13491 10915 13557 10916
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18646 10845 18706 15403
rect 18830 12749 18890 17987
rect 19195 16148 19261 16149
rect 19195 16084 19196 16148
rect 19260 16084 19261 16148
rect 19195 16083 19261 16084
rect 19011 16012 19077 16013
rect 19011 15948 19012 16012
rect 19076 15948 19077 16012
rect 19011 15947 19077 15948
rect 19014 12885 19074 15947
rect 19011 12884 19077 12885
rect 19011 12820 19012 12884
rect 19076 12820 19077 12884
rect 19011 12819 19077 12820
rect 18827 12748 18893 12749
rect 18827 12684 18828 12748
rect 18892 12684 18893 12748
rect 18827 12683 18893 12684
rect 19011 12612 19077 12613
rect 19011 12548 19012 12612
rect 19076 12548 19077 12612
rect 19011 12547 19077 12548
rect 18643 10844 18709 10845
rect 18643 10780 18644 10844
rect 18708 10780 18709 10844
rect 18643 10779 18709 10780
rect 18827 10708 18893 10709
rect 18827 10644 18828 10708
rect 18892 10644 18893 10708
rect 18827 10643 18893 10644
rect 18830 9893 18890 10643
rect 18827 9892 18893 9893
rect 18827 9828 18828 9892
rect 18892 9828 18893 9892
rect 18827 9827 18893 9828
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 19014 9757 19074 12547
rect 19198 11797 19258 16083
rect 19195 11796 19261 11797
rect 19195 11732 19196 11796
rect 19260 11732 19261 11796
rect 19195 11731 19261 11732
rect 19011 9756 19077 9757
rect 19011 9692 19012 9756
rect 19076 9692 19077 9756
rect 19011 9691 19077 9692
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606256979
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606256979
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4692 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1606256979
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1606256979
transform 1 0 5612 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606256979
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1606256979
transform 1 0 5244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_55
timestamp 1606256979
transform 1 0 6164 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606256979
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1606256979
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606256979
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1606256979
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1606256979
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1606256979
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1606256979
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1606256979
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1606256979
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1606256979
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1606256979
transform 1 0 15180 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1606256979
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_147
timestamp 1606256979
transform 1 0 14628 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1606256979
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1606256979
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1606256979
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1606256979
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1606256979
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1606256979
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1606256979
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1606256979
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1606256979
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1606256979
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606256979
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606256979
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606256979
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1606256979
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1606256979
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1606256979
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1606256979
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1606256979
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1606256979
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1606256979
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1606256979
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1606256979
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1606256979
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1606256979
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606256979
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606256979
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606256979
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606256979
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606256979
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1606256979
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1606256979
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1606256979
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1606256979
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1606256979
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1606256979
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1606256979
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1606256979
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1606256979
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1606256979
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1606256979
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606256979
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606256979
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606256979
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1606256979
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1606256979
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1606256979
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1606256979
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1606256979
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1606256979
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1606256979
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1606256979
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1606256979
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1606256979
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1606256979
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606256979
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606256979
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606256979
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606256979
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606256979
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606256979
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606256979
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1606256979
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1606256979
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1606256979
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1606256979
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1606256979
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1606256979
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1606256979
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1606256979
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1606256979
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 20056 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_196
timestamp 1606256979
transform 1 0 19136 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1606256979
transform 1 0 20884 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1606256979
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1606256979
transform 1 0 2944 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606256979
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1606256979
transform 1 0 2484 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_19
timestamp 1606256979
transform 1 0 2852 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606256979
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_29
timestamp 1606256979
transform 1 0 3772 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_41
timestamp 1606256979
transform 1 0 4876 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1606256979
transform 1 0 4968 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1606256979
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1606256979
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606256979
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606256979
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1606256979
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1606256979
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1606256979
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1606256979
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1606256979
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1606256979
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1606256979
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1606256979
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1606256979
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1606256979
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1606256979
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1606256979
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1606256979
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1606256979
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1606256979
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1606256979
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1606256979
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 19320 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19780 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1606256979
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_202
timestamp 1606256979
transform 1 0 19688 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_196
timestamp 1606256979
transform 1 0 19136 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1606256979
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606256979
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606256979
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_214
timestamp 1606256979
transform 1 0 20792 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 1564 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3312 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1606256979
transform 1 0 4140 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_21
timestamp 1606256979
transform 1 0 3036 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606256979
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_32
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6164 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1606256979
transform 1 0 5152 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_42
timestamp 1606256979
transform 1 0 4968 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 1606256979
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1606256979
transform 1 0 7176 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_64
timestamp 1606256979
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_75
timestamp 1606256979
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1606256979
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1606256979
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1606256979
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1606256979
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1606256979
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1606256979
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_166
timestamp 1606256979
transform 1 0 16376 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16652 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_8_185
timestamp 1606256979
transform 1 0 18124 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 19136 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1606256979
transform 1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606256979
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1606256979
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_218
timestamp 1606256979
transform 1 0 21160 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2484 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1606256979
transform 1 0 1472 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_13
timestamp 1606256979
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606256979
transform 1 0 4508 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_31
timestamp 1606256979
transform 1 0 3956 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1606256979
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4968 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1606256979
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_62
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6900 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8556 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1606256979
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_90
timestamp 1606256979
transform 1 0 9384 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_102
timestamp 1606256979
transform 1 0 10488 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_114
timestamp 1606256979
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1606256979
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1606256979
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_159
timestamp 1606256979
transform 1 0 15732 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_165
timestamp 1606256979
transform 1 0 16284 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_175
timestamp 1606256979
transform 1 0 17204 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 19872 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19136 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1606256979
transform 1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_202
timestamp 1606256979
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_213
timestamp 1606256979
transform 1 0 20700 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1606256979
transform 1 0 21252 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2576 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_15
timestamp 1606256979
transform 1 0 2484 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_25
timestamp 1606256979
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp 1606256979
transform 1 0 4876 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 5704 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 1606256979
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7820 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_10_66
timestamp 1606256979
transform 1 0 7176 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_72
timestamp 1606256979
transform 1 0 7728 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9936 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1606256979
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_93
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12328 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1606256979
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_117
timestamp 1606256979
transform 1 0 11868 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_121
timestamp 1606256979
transform 1 0 12236 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_131
timestamp 1606256979
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_143
timestamp 1606256979
transform 1 0 14260 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606256979
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_166
timestamp 1606256979
transform 1 0 16376 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16836 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_170
timestamp 1606256979
transform 1 0 16744 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_187
timestamp 1606256979
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 19412 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_10_208
timestamp 1606256979
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606256979
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606256979
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1472 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_20
timestamp 1606256979
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4324 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 3128 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_31
timestamp 1606256979
transform 1 0 3956 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1606256979
transform 1 0 5336 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_44
timestamp 1606256979
transform 1 0 5152 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_55
timestamp 1606256979
transform 1 0 6164 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_62
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8556 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7544 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_79
timestamp 1606256979
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10212 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_97
timestamp 1606256979
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11224 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_108
timestamp 1606256979
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 1606256979
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_139
timestamp 1606256979
transform 1 0 13892 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1606256979
transform 1 0 15732 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 14720 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_147
timestamp 1606256979
transform 1 0 14628 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_157
timestamp 1606256979
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 18032 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16928 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_168
timestamp 1606256979
transform 1 0 16560 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1606256979
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 19688 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1606256979
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 20700 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_211
timestamp 1606256979
transform 1 0 20516 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_217
timestamp 1606256979
transform 1 0 21068 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1472 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1606256979
transform 1 0 2208 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_10
timestamp 1606256979
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1606256979
transform 1 0 4416 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_21
timestamp 1606256979
transform 1 0 3036 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1606256979
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1606256979
transform 1 0 5428 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_45
timestamp 1606256979
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_56
timestamp 1606256979
transform 1 0 6256 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1606256979
transform 1 0 7084 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8096 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_64
timestamp 1606256979
transform 1 0 6992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_74
timestamp 1606256979
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1606256979
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1606256979
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_102
timestamp 1606256979
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11868 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10764 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_114
timestamp 1606256979
transform 1 0 11592 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 13524 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1606256979
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 16284 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1606256979
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1606256979
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 18216 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_12_174
timestamp 1606256979
transform 1 0 17112 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19872 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_202
timestamp 1606256979
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606256979
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1606256979
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_218
timestamp 1606256979
transform 1 0 21160 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1606256979
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1606256979
transform 1 0 1840 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1748 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_17
timestamp 1606256979
transform 1 0 2668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1606256979
transform 1 0 2300 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606256979
transform 1 0 2852 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2668 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606256979
transform 1 0 3496 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1606256979
transform 1 0 4324 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_33
timestamp 1606256979
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_23
timestamp 1606256979
transform 1 0 3220 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1606256979
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1606256979
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5428 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1606256979
transform 1 0 5336 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_left_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5060 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_44
timestamp 1606256979
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_55
timestamp 1606256979
transform 1 0 6164 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_62
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 1606256979
transform 1 0 5336 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606256979
transform 1 0 7452 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7912 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7544 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_14_63
timestamp 1606256979
transform 1 0 6900 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp 1606256979
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9936 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_86
timestamp 1606256979
transform 1 0 9016 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_94
timestamp 1606256979
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606256979
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_102
timestamp 1606256979
transform 1 0 10488 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 11224 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_112
timestamp 1606256979
transform 1 0 11408 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1606256979
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_126
timestamp 1606256979
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1606256979
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12880 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606256979
transform 1 0 13432 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1606256979
transform 1 0 14076 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_137
timestamp 1606256979
transform 1 0 13708 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_143
timestamp 1606256979
transform 1 0 14260 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_137
timestamp 1606256979
transform 1 0 13708 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 14168 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606256979
transform 1 0 14352 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 14812 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16284 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1606256979
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_165
timestamp 1606256979
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1606256979
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1606256979
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606256979
transform 1 0 17940 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1606256979
transform 1 0 16468 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 18124 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_176
timestamp 1606256979
transform 1 0 17296 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1606256979
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_184
timestamp 1606256979
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_181
timestamp 1606256979
transform 1 0 17756 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_187
timestamp 1606256979
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 19688 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 20148 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 19136 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 18492 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_194
timestamp 1606256979
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_205
timestamp 1606256979
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_198
timestamp 1606256979
transform 1 0 19320 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_216
timestamp 1606256979
transform 1 0 20976 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1606256979
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606256979
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606256979
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1606256979
transform 1 0 2668 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1606256979
transform 1 0 1656 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_15
timestamp 1606256979
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1606256979
transform 1 0 4876 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1606256979
transform 1 0 3864 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_26
timestamp 1606256979
transform 1 0 3496 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_39
timestamp 1606256979
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_50
timestamp 1606256979
transform 1 0 5704 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_58
timestamp 1606256979
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8648 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1606256979
transform 1 0 7268 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 8280 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1606256979
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_76
timestamp 1606256979
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_81
timestamp 1606256979
transform 1 0 8556 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10672 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9660 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_91
timestamp 1606256979
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_102
timestamp 1606256979
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606256979
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1606256979
transform 1 0 13616 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_132
timestamp 1606256979
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1606256979
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1606256979
transform 1 0 14904 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16100 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 14628 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1606256979
transform 1 0 15732 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_172
timestamp 1606256979
transform 1 0 16928 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1606256979
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1606256979
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1606256979
transform 1 0 19412 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1606256979
transform 1 0 18400 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1606256979
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_208
timestamp 1606256979
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 20424 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_216
timestamp 1606256979
transform 1 0 20976 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1472 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1606256979
transform 1 0 2944 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_28
timestamp 1606256979
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6716 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5704 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_48
timestamp 1606256979
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1606256979
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_70
timestamp 1606256979
transform 1 0 7544 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_78
timestamp 1606256979
transform 1 0 8280 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10396 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606256979
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12236 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 11960 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_110
timestamp 1606256979
transform 1 0 11224 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13248 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 14260 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_130
timestamp 1606256979
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1606256979
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606256979
transform 1 0 14720 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_146
timestamp 1606256979
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1606256979
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606256979
transform 1 0 18308 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16928 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1606256979
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_181
timestamp 1606256979
transform 1 0 17756 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19964 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1606256979
transform 1 0 18860 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_191
timestamp 1606256979
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_202
timestamp 1606256979
transform 1 0 19688 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606256979
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_211
timestamp 1606256979
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_218
timestamp 1606256979
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2116 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_20
timestamp 1606256979
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4140 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1606256979
transform 1 0 3128 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_31
timestamp 1606256979
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_42
timestamp 1606256979
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_53
timestamp 1606256979
transform 1 0 5980 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1606256979
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 8188 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7176 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_75
timestamp 1606256979
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10028 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1606256979
transform 1 0 9660 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11040 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_106
timestamp 1606256979
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1606256979
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1606256979
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_123
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13064 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1606256979
transform 1 0 12972 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 16008 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1606256979
transform 1 0 14720 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_146
timestamp 1606256979
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_157
timestamp 1606256979
transform 1 0 15548 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_161
timestamp 1606256979
transform 1 0 15916 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606256979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_178
timestamp 1606256979
transform 1 0 17480 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1606256979
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1606256979
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606256979
transform 1 0 18400 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1606256979
transform 1 0 18952 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1606256979
transform 1 0 19964 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_192
timestamp 1606256979
transform 1 0 18768 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1606256979
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_214
timestamp 1606256979
transform 1 0 20792 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 1564 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4416 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_21
timestamp 1606256979
transform 1 0 3036 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1606256979
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6072 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1606256979
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7728 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_70
timestamp 1606256979
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10212 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1606256979
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_93
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11224 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_108
timestamp 1606256979
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12880 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_126
timestamp 1606256979
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_144
timestamp 1606256979
transform 1 0 14352 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606256979
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1606256979
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1606256979
transform 1 0 16100 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 16468 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_183
timestamp 1606256979
transform 1 0 17940 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1606256979
transform 1 0 18584 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1606256979
transform 1 0 19596 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1606256979
transform 1 0 18492 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_199
timestamp 1606256979
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1606256979
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606256979
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1606256979
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_218
timestamp 1606256979
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_9
timestamp 1606256979
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1606256979
transform 1 0 1472 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606256979
transform 1 0 1564 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_13
timestamp 1606256979
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2116 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_17
timestamp 1606256979
transform 1 0 2668 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2484 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606256979
transform 1 0 4232 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1606256979
transform 1 0 4692 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1606256979
transform 1 0 4416 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_31
timestamp 1606256979
transform 1 0 3956 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1606256979
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1606256979
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5428 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1606256979
transform 1 0 6440 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1606256979
transform 1 0 5704 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_48
timestamp 1606256979
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606256979
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_45
timestamp 1606256979
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_56
timestamp 1606256979
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7452 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1606256979
transform 1 0 8188 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1606256979
transform 1 0 7176 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_75
timestamp 1606256979
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_67
timestamp 1606256979
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_93
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606256979
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1606256979
transform 1 0 8924 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1606256979
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_86
timestamp 1606256979
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 9660 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606256979
transform 1 0 9200 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_100
timestamp 1606256979
transform 1 0 10304 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1606256979
transform 1 0 9936 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_left_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10396 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10028 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11500 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1606256979
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_123
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 14260 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12972 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13800 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13248 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 12696 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_129
timestamp 1606256979
transform 1 0 12972 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_141
timestamp 1606256979
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606256979
transform 1 0 14628 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16284 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1606256979
transform 1 0 15916 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_159
timestamp 1606256979
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1606256979
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1606256979
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 17940 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1606256979
transform 1 0 16928 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18216 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606256979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1606256979
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1606256979
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1606256979
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_181
timestamp 1606256979
transform 1 0 17756 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1606256979
transform 1 0 19964 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 18952 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1606256979
transform 1 0 19596 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_192
timestamp 1606256979
transform 1 0 18768 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 1606256979
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_199
timestamp 1606256979
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606256979
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_214
timestamp 1606256979
transform 1 0 20792 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1606256979
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606256979
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606256979
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606256979
transform 1 0 2392 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606256979
transform 1 0 2944 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1656 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1606256979
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_18
timestamp 1606256979
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 3680 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_24
timestamp 1606256979
transform 1 0 3312 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5336 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_44
timestamp 1606256979
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_55
timestamp 1606256979
transform 1 0 6164 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7268 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_66
timestamp 1606256979
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_83
timestamp 1606256979
transform 1 0 8740 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9660 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10488 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1606256979
transform 1 0 8832 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 11316 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1606256979
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606256979
transform 1 0 12788 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 13340 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_131
timestamp 1606256979
transform 1 0 13156 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1606256979
transform 1 0 16008 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1606256979
transform 1 0 14996 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1606256979
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_160
timestamp 1606256979
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606256979
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 17204 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606256979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_171
timestamp 1606256979
transform 1 0 16836 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1606256979
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 18584 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 20240 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1606256979
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1606256979
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_217
timestamp 1606256979
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606256979
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 2576 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_11
timestamp 1606256979
transform 1 0 2116 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_15
timestamp 1606256979
transform 1 0 2484 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4416 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_25
timestamp 1606256979
transform 1 0 3404 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6072 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1606256979
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1606256979
transform 1 0 7728 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_70
timestamp 1606256979
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_81
timestamp 1606256979
transform 1 0 8556 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606256979
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1606256979
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_102
timestamp 1606256979
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1606256979
transform 1 0 10764 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12236 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11224 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_108
timestamp 1606256979
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_119
timestamp 1606256979
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1606256979
transform 1 0 14168 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 13892 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_137
timestamp 1606256979
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1606256979
transform 1 0 15364 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15916 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1606256979
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_154
timestamp 1606256979
transform 1 0 15272 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_159
timestamp 1606256979
transform 1 0 15732 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 16928 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_170
timestamp 1606256979
transform 1 0 16744 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1606256979
transform 1 0 19596 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 18584 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1606256979
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_199
timestamp 1606256979
transform 1 0 19412 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606256979
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1606256979
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1606256979
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1606256979
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2208 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1472 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1606256979
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_10
timestamp 1606256979
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4416 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_28
timestamp 1606256979
transform 1 0 3680 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606256979
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_45
timestamp 1606256979
transform 1 0 5244 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1606256979
transform 1 0 6348 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8372 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 7820 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1606256979
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_76
timestamp 1606256979
transform 1 0 8096 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1606256979
transform 1 0 9384 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10396 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_88
timestamp 1606256979
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_99
timestamp 1606256979
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606256979
transform 1 0 11776 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12604 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606256979
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_110
timestamp 1606256979
transform 1 0 11224 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1606256979
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1606256979
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606256979
transform 1 0 14076 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_134
timestamp 1606256979
transform 1 0 13432 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_140
timestamp 1606256979
transform 1 0 13984 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_145
timestamp 1606256979
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16008 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1606256979
transform 1 0 14628 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 15732 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_156
timestamp 1606256979
transform 1 0 15456 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18032 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606256979
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_178
timestamp 1606256979
transform 1 0 17480 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1606256979
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1606256979
transform 1 0 19688 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1606256979
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606256979
transform 1 0 20700 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_211
timestamp 1606256979
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_217
timestamp 1606256979
transform 1 0 21068 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606256979
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1606256979
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_11
timestamp 1606256979
transform 1 0 2116 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1606256979
transform 1 0 3496 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606256979
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_23
timestamp 1606256979
transform 1 0 3220 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1606256979
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1606256979
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 5060 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_52
timestamp 1606256979
transform 1 0 5888 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606256979
transform 1 0 7084 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1606256979
transform 1 0 7544 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_64
timestamp 1606256979
transform 1 0 6992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_68
timestamp 1606256979
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_79
timestamp 1606256979
transform 1 0 8372 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606256979
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1606256979
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12328 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11316 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_109
timestamp 1606256979
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_120
timestamp 1606256979
transform 1 0 12144 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13340 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1606256979
transform 1 0 14076 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_131
timestamp 1606256979
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_139
timestamp 1606256979
transform 1 0 13892 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606256979
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15732 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606256979
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1606256979
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1606256979
transform 1 0 15548 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1606256979
transform 1 0 17756 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 16744 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_168
timestamp 1606256979
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_179
timestamp 1606256979
transform 1 0 17572 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19780 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1606256979
transform 1 0 18768 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_190
timestamp 1606256979
transform 1 0 18584 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_201
timestamp 1606256979
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606256979
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1606256979
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606256979
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606256979
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606256979
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2576 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1606256979
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_11
timestamp 1606256979
transform 1 0 2116 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1606256979
transform 1 0 2484 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 4324 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_32
timestamp 1606256979
transform 1 0 4048 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606256979
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 5336 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_44
timestamp 1606256979
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_49
timestamp 1606256979
transform 1 0 5612 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1606256979
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1606256979
transform 1 0 7912 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6900 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_72
timestamp 1606256979
transform 1 0 7728 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_83
timestamp 1606256979
transform 1 0 8740 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10028 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9016 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_95
timestamp 1606256979
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12512 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606256979
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1606256979
transform 1 0 11500 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_123
timestamp 1606256979
transform 1 0 12420 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 14168 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_140
timestamp 1606256979
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15824 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_158
timestamp 1606256979
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606256979
transform 1 0 17480 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18032 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606256979
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_176
timestamp 1606256979
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1606256979
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18860 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_190
timestamp 1606256979
transform 1 0 18584 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 20516 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1606256979
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_217
timestamp 1606256979
transform 1 0 21068 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1606256979
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1606256979
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606256979
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606256979
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_17
timestamp 1606256979
transform 1 0 2668 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1606256979
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_15
timestamp 1606256979
transform 1 0 2484 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1606256979
transform 1 0 2116 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2576 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1606256979
transform 1 0 2300 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4048 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4600 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 3588 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606256979
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_25
timestamp 1606256979
transform 1 0 3404 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_25
timestamp 1606256979
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_36
timestamp 1606256979
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 6072 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606256979
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_48
timestamp 1606256979
transform 1 0 5520 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_54
timestamp 1606256979
transform 1 0 6072 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1606256979
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7728 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1606256979
transform 1 0 7820 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_70
timestamp 1606256979
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_71
timestamp 1606256979
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_82
timestamp 1606256979
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8832 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9660 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606256979
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1606256979
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_102
timestamp 1606256979
transform 1 0 10488 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_90
timestamp 1606256979
transform 1 0 9384 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_102
timestamp 1606256979
transform 1 0 10488 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1606256979
transform 1 0 10764 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11316 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11224 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606256979
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_110
timestamp 1606256979
transform 1 0 11224 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1606256979
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_119
timestamp 1606256979
transform 1 0 12052 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_123
timestamp 1606256979
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13892 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12972 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12880 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1606256979
transform 1 0 14076 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1606256979
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_138
timestamp 1606256979
transform 1 0 13800 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_127
timestamp 1606256979
transform 1 0 12788 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1606256979
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_148
timestamp 1606256979
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1606256979
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606256979
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14904 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1606256979
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_162
timestamp 1606256979
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_156
timestamp 1606256979
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1606256979
transform 1 0 16100 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1606256979
transform 1 0 15640 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1606256979
transform 1 0 16192 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 18216 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 16468 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1606256979
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 16928 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606256979
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_183
timestamp 1606256979
transform 1 0 17940 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_168
timestamp 1606256979
transform 1 0 16560 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1606256979
transform 1 0 17480 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1606256979
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606256979
transform 1 0 20056 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19872 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1606256979
transform 1 0 19044 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_202
timestamp 1606256979
transform 1 0 19688 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1606256979
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_204
timestamp 1606256979
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1606256979
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1606256979
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606256979
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1606256979
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_218
timestamp 1606256979
transform 1 0 21160 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606256979
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1606256979
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1606256979
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1606256979
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606256979
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606256979
transform 1 0 2300 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606256979
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1606256979
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1606256979
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_17
timestamp 1606256979
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606256979
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_23
timestamp 1606256979
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_41
timestamp 1606256979
transform 1 0 4876 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5612 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 7268 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_left_track_1.prog_clk
timestamp 1606256979
transform 1 0 8280 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_65
timestamp 1606256979
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_76
timestamp 1606256979
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606256979
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1606256979
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1606256979
transform 1 0 12328 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11316 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1606256979
transform 1 0 11132 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_120
timestamp 1606256979
transform 1 0 12144 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606256979
transform 1 0 13984 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14444 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12880 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_126
timestamp 1606256979
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1606256979
transform 1 0 13708 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_143
timestamp 1606256979
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1606256979
transform 1 0 16284 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1606256979
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606256979
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1606256979
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1606256979
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1606256979
transform 1 0 17848 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16836 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_169
timestamp 1606256979
transform 1 0 16652 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_180
timestamp 1606256979
transform 1 0 17664 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_186
timestamp 1606256979
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606256979
transform 1 0 18400 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18952 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_192
timestamp 1606256979
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606256979
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606256979
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_210
timestamp 1606256979
transform 1 0 20424 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606256979
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606256979
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1606256979
transform 1 0 2300 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1606256979
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2852 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606256979
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1606256979
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1606256979
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1606256979
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 4600 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_25
timestamp 1606256979
transform 1 0 3404 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_37
timestamp 1606256979
transform 1 0 4508 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606256979
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1606256979
transform 1 0 5152 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_56
timestamp 1606256979
transform 1 0 6256 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_60
timestamp 1606256979
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1606256979
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1606256979
transform 1 0 8188 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6992 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_73
timestamp 1606256979
transform 1 0 7820 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10120 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 9200 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_86
timestamp 1606256979
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_94
timestamp 1606256979
transform 1 0 9752 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1606256979
transform 1 0 11776 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1606256979
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606256979
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1606256979
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1606256979
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 14260 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12880 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_126
timestamp 1606256979
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_137
timestamp 1606256979
transform 1 0 13708 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15916 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_159
timestamp 1606256979
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606256979
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16928 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606256979
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_170
timestamp 1606256979
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1606256979
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18584 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1606256979
transform 1 0 19596 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_188
timestamp 1606256979
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_199
timestamp 1606256979
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606256979
transform 1 0 20608 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606256979
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1606256979
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_216
timestamp 1606256979
transform 1 0 20976 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1606256979
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1606256979
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606256979
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1606256979
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_11
timestamp 1606256979
transform 1 0 2116 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_19
timestamp 1606256979
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606256979
transform 1 0 3036 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606256979
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606256979
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_25
timestamp 1606256979
transform 1 0 3404 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_36
timestamp 1606256979
transform 1 0 4416 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1606256979
transform 1 0 5428 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 6256 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_44
timestamp 1606256979
transform 1 0 5152 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_51
timestamp 1606256979
transform 1 0 5796 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_55
timestamp 1606256979
transform 1 0 6164 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_62
timestamp 1606256979
transform 1 0 6808 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1606256979
transform 1 0 7176 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7728 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_70
timestamp 1606256979
transform 1 0 7544 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606256979
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1606256979
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11408 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12144 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_30_109
timestamp 1606256979
transform 1 0 11132 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_118
timestamp 1606256979
transform 1 0 11960 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13156 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_129
timestamp 1606256979
transform 1 0 12972 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15456 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606256979
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_147
timestamp 1606256979
transform 1 0 14628 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1606256979
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 17112 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_172
timestamp 1606256979
transform 1 0 16928 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18768 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1606256979
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_208
timestamp 1606256979
transform 1 0 20240 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606256979
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606256979
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606256979
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606256979
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1606256979
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1606256979
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606256979
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1606256979
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1606256979
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_17
timestamp 1606256979
transform 1 0 2668 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1606256979
transform 1 0 3220 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3772 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_27
timestamp 1606256979
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_41
timestamp 1606256979
transform 1 0 4876 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1606256979
transform 1 0 5888 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606256979
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_49
timestamp 1606256979
transform 1 0 5612 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_56
timestamp 1606256979
transform 1 0 6256 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1606256979
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_62
timestamp 1606256979
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7176 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_82
timestamp 1606256979
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1606256979
transform 1 0 9844 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10396 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8832 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_93
timestamp 1606256979
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_98
timestamp 1606256979
transform 1 0 10120 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606256979
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_117
timestamp 1606256979
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1606256979
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14076 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1606256979
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1606256979
transform 1 0 14812 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15824 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_147
timestamp 1606256979
transform 1 0 14628 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_158
timestamp 1606256979
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_166
timestamp 1606256979
transform 1 0 16376 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16928 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606256979
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1606256979
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606256979
transform 1 0 18768 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606256979
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19228 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_190
timestamp 1606256979
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_195
timestamp 1606256979
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1606256979
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606256979
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606256979
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1606256979
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1606256979
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1606256979
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1606256979
transform 1 0 2392 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1606256979
transform 1 0 1840 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606256979
transform 1 0 2944 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606256979
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1606256979
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1606256979
transform 1 0 1748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_12
timestamp 1606256979
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_18
timestamp 1606256979
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606256979
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_24
timestamp 1606256979
transform 1 0 3312 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1606256979
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1606256979
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606256979
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1606256979
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1606256979
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8280 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606256979
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_75
timestamp 1606256979
transform 1 0 8004 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9844 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606256979
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1606256979
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_94
timestamp 1606256979
transform 1 0 9752 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_104
timestamp 1606256979
transform 1 0 10672 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10948 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606256979
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_116
timestamp 1606256979
transform 1 0 11776 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_125
timestamp 1606256979
transform 1 0 12604 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606256979
transform 1 0 14168 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12880 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_137
timestamp 1606256979
transform 1 0 13708 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1606256979
transform 1 0 14076 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606256979
transform 1 0 14720 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1606256979
transform 1 0 16376 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1606256979
transform 1 0 15824 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606256979
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_146
timestamp 1606256979
transform 1 0 14536 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_152
timestamp 1606256979
transform 1 0 15088 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1606256979
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_164
timestamp 1606256979
transform 1 0 16192 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606256979
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606256979
transform 1 0 17480 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1606256979
transform 1 0 16928 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606256979
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_170
timestamp 1606256979
transform 1 0 16744 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_176
timestamp 1606256979
transform 1 0 17296 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_182
timestamp 1606256979
transform 1 0 17848 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606256979
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606256979
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606256979
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp 1606256979
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1606256979
transform 1 0 19228 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1606256979
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606256979
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606256979
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606256979
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1606256979
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1606256979
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606256979
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 202 22320 258 22800 6 SC_IN_TOP
port 0 nsew default input
rlabel metal2 s 22558 22320 22614 22800 6 SC_OUT_TOP
port 1 nsew default tristate
rlabel metal2 s 4342 22320 4398 22800 6 Test_en_N_out
port 2 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 Test_en_S_in
port 3 nsew default input
rlabel metal2 s 2226 0 2282 480 6 ccff_head
port 4 nsew default input
rlabel metal2 s 6734 0 6790 480 6 ccff_tail
port 5 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[0]
port 6 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[10]
port 7 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[11]
port 8 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[12]
port 9 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[13]
port 10 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[14]
port 11 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[15]
port 12 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[16]
port 13 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[17]
port 14 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[18]
port 15 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[19]
port 16 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[1]
port 17 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[2]
port 18 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[3]
port 19 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[4]
port 20 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[5]
port 21 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[6]
port 22 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[7]
port 23 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[8]
port 24 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[9]
port 25 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[0]
port 26 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[10]
port 27 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[11]
port 28 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[12]
port 29 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[13]
port 30 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[14]
port 31 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[15]
port 32 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 33 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[17]
port 34 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 35 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[19]
port 36 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[1]
port 37 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[2]
port 38 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[4]
port 40 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[5]
port 41 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[6]
port 42 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[7]
port 43 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[8]
port 44 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[9]
port 45 nsew default tristate
rlabel metal3 s 22320 4224 22800 4344 6 chanx_right_in[0]
port 46 nsew default input
rlabel metal3 s 22320 8984 22800 9104 6 chanx_right_in[10]
port 47 nsew default input
rlabel metal3 s 22320 9392 22800 9512 6 chanx_right_in[11]
port 48 nsew default input
rlabel metal3 s 22320 9936 22800 10056 6 chanx_right_in[12]
port 49 nsew default input
rlabel metal3 s 22320 10344 22800 10464 6 chanx_right_in[13]
port 50 nsew default input
rlabel metal3 s 22320 10752 22800 10872 6 chanx_right_in[14]
port 51 nsew default input
rlabel metal3 s 22320 11296 22800 11416 6 chanx_right_in[15]
port 52 nsew default input
rlabel metal3 s 22320 11704 22800 11824 6 chanx_right_in[16]
port 53 nsew default input
rlabel metal3 s 22320 12248 22800 12368 6 chanx_right_in[17]
port 54 nsew default input
rlabel metal3 s 22320 12656 22800 12776 6 chanx_right_in[18]
port 55 nsew default input
rlabel metal3 s 22320 13200 22800 13320 6 chanx_right_in[19]
port 56 nsew default input
rlabel metal3 s 22320 4768 22800 4888 6 chanx_right_in[1]
port 57 nsew default input
rlabel metal3 s 22320 5176 22800 5296 6 chanx_right_in[2]
port 58 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 chanx_right_in[3]
port 59 nsew default input
rlabel metal3 s 22320 6128 22800 6248 6 chanx_right_in[4]
port 60 nsew default input
rlabel metal3 s 22320 6672 22800 6792 6 chanx_right_in[5]
port 61 nsew default input
rlabel metal3 s 22320 7080 22800 7200 6 chanx_right_in[6]
port 62 nsew default input
rlabel metal3 s 22320 7488 22800 7608 6 chanx_right_in[7]
port 63 nsew default input
rlabel metal3 s 22320 8032 22800 8152 6 chanx_right_in[8]
port 64 nsew default input
rlabel metal3 s 22320 8440 22800 8560 6 chanx_right_in[9]
port 65 nsew default input
rlabel metal3 s 22320 13608 22800 13728 6 chanx_right_out[0]
port 66 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[10]
port 67 nsew default tristate
rlabel metal3 s 22320 18776 22800 18896 6 chanx_right_out[11]
port 68 nsew default tristate
rlabel metal3 s 22320 19184 22800 19304 6 chanx_right_out[12]
port 69 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 chanx_right_out[13]
port 70 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[14]
port 71 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 chanx_right_out[15]
port 72 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[16]
port 73 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[17]
port 74 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 chanx_right_out[18]
port 75 nsew default tristate
rlabel metal3 s 22320 22448 22800 22568 6 chanx_right_out[19]
port 76 nsew default tristate
rlabel metal3 s 22320 14016 22800 14136 6 chanx_right_out[1]
port 77 nsew default tristate
rlabel metal3 s 22320 14560 22800 14680 6 chanx_right_out[2]
port 78 nsew default tristate
rlabel metal3 s 22320 14968 22800 15088 6 chanx_right_out[3]
port 79 nsew default tristate
rlabel metal3 s 22320 15512 22800 15632 6 chanx_right_out[4]
port 80 nsew default tristate
rlabel metal3 s 22320 15920 22800 16040 6 chanx_right_out[5]
port 81 nsew default tristate
rlabel metal3 s 22320 16464 22800 16584 6 chanx_right_out[6]
port 82 nsew default tristate
rlabel metal3 s 22320 16872 22800 16992 6 chanx_right_out[7]
port 83 nsew default tristate
rlabel metal3 s 22320 17280 22800 17400 6 chanx_right_out[8]
port 84 nsew default tristate
rlabel metal3 s 22320 17824 22800 17944 6 chanx_right_out[9]
port 85 nsew default tristate
rlabel metal2 s 5630 22320 5686 22800 6 chany_top_in[0]
port 86 nsew default input
rlabel metal2 s 9862 22320 9918 22800 6 chany_top_in[10]
port 87 nsew default input
rlabel metal2 s 10322 22320 10378 22800 6 chany_top_in[11]
port 88 nsew default input
rlabel metal2 s 10690 22320 10746 22800 6 chany_top_in[12]
port 89 nsew default input
rlabel metal2 s 11150 22320 11206 22800 6 chany_top_in[13]
port 90 nsew default input
rlabel metal2 s 11610 22320 11666 22800 6 chany_top_in[14]
port 91 nsew default input
rlabel metal2 s 11978 22320 12034 22800 6 chany_top_in[15]
port 92 nsew default input
rlabel metal2 s 12438 22320 12494 22800 6 chany_top_in[16]
port 93 nsew default input
rlabel metal2 s 12806 22320 12862 22800 6 chany_top_in[17]
port 94 nsew default input
rlabel metal2 s 13266 22320 13322 22800 6 chany_top_in[18]
port 95 nsew default input
rlabel metal2 s 13634 22320 13690 22800 6 chany_top_in[19]
port 96 nsew default input
rlabel metal2 s 6090 22320 6146 22800 6 chany_top_in[1]
port 97 nsew default input
rlabel metal2 s 6458 22320 6514 22800 6 chany_top_in[2]
port 98 nsew default input
rlabel metal2 s 6918 22320 6974 22800 6 chany_top_in[3]
port 99 nsew default input
rlabel metal2 s 7378 22320 7434 22800 6 chany_top_in[4]
port 100 nsew default input
rlabel metal2 s 7746 22320 7802 22800 6 chany_top_in[5]
port 101 nsew default input
rlabel metal2 s 8206 22320 8262 22800 6 chany_top_in[6]
port 102 nsew default input
rlabel metal2 s 8574 22320 8630 22800 6 chany_top_in[7]
port 103 nsew default input
rlabel metal2 s 9034 22320 9090 22800 6 chany_top_in[8]
port 104 nsew default input
rlabel metal2 s 9494 22320 9550 22800 6 chany_top_in[9]
port 105 nsew default input
rlabel metal2 s 14094 22320 14150 22800 6 chany_top_out[0]
port 106 nsew default tristate
rlabel metal2 s 18326 22320 18382 22800 6 chany_top_out[10]
port 107 nsew default tristate
rlabel metal2 s 18786 22320 18842 22800 6 chany_top_out[11]
port 108 nsew default tristate
rlabel metal2 s 19154 22320 19210 22800 6 chany_top_out[12]
port 109 nsew default tristate
rlabel metal2 s 19614 22320 19670 22800 6 chany_top_out[13]
port 110 nsew default tristate
rlabel metal2 s 19982 22320 20038 22800 6 chany_top_out[14]
port 111 nsew default tristate
rlabel metal2 s 20442 22320 20498 22800 6 chany_top_out[15]
port 112 nsew default tristate
rlabel metal2 s 20902 22320 20958 22800 6 chany_top_out[16]
port 113 nsew default tristate
rlabel metal2 s 21270 22320 21326 22800 6 chany_top_out[17]
port 114 nsew default tristate
rlabel metal2 s 21730 22320 21786 22800 6 chany_top_out[18]
port 115 nsew default tristate
rlabel metal2 s 22098 22320 22154 22800 6 chany_top_out[19]
port 116 nsew default tristate
rlabel metal2 s 14554 22320 14610 22800 6 chany_top_out[1]
port 117 nsew default tristate
rlabel metal2 s 14922 22320 14978 22800 6 chany_top_out[2]
port 118 nsew default tristate
rlabel metal2 s 15382 22320 15438 22800 6 chany_top_out[3]
port 119 nsew default tristate
rlabel metal2 s 15750 22320 15806 22800 6 chany_top_out[4]
port 120 nsew default tristate
rlabel metal2 s 16210 22320 16266 22800 6 chany_top_out[5]
port 121 nsew default tristate
rlabel metal2 s 16670 22320 16726 22800 6 chany_top_out[6]
port 122 nsew default tristate
rlabel metal2 s 17038 22320 17094 22800 6 chany_top_out[7]
port 123 nsew default tristate
rlabel metal2 s 17498 22320 17554 22800 6 chany_top_out[8]
port 124 nsew default tristate
rlabel metal2 s 17866 22320 17922 22800 6 chany_top_out[9]
port 125 nsew default tristate
rlabel metal2 s 4802 22320 4858 22800 6 clk_3_N_out
port 126 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 clk_3_S_in
port 127 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_11_
port 128 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_13_
port 129 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_15_
port 130 nsew default input
rlabel metal3 s 0 3816 480 3936 6 left_bottom_grid_pin_17_
port 131 nsew default input
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_1_
port 132 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_3_
port 133 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_5_
port 134 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_7_
port 135 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_9_
port 136 nsew default input
rlabel metal2 s 3974 22320 4030 22800 6 prog_clk_0_N_in
port 137 nsew default input
rlabel metal2 s 5262 22320 5318 22800 6 prog_clk_3_N_out
port 138 nsew default tristate
rlabel metal2 s 11334 0 11390 480 6 prog_clk_3_S_in
port 139 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_11_
port 140 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_13_
port 141 nsew default input
rlabel metal3 s 22320 3408 22800 3528 6 right_bottom_grid_pin_15_
port 142 nsew default input
rlabel metal3 s 22320 3816 22800 3936 6 right_bottom_grid_pin_17_
port 143 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_1_
port 144 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_3_
port 145 nsew default input
rlabel metal3 s 22320 960 22800 1080 6 right_bottom_grid_pin_5_
port 146 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_7_
port 147 nsew default input
rlabel metal3 s 22320 1912 22800 2032 6 right_bottom_grid_pin_9_
port 148 nsew default input
rlabel metal2 s 570 22320 626 22800 6 top_left_grid_pin_42_
port 149 nsew default input
rlabel metal2 s 1030 22320 1086 22800 6 top_left_grid_pin_43_
port 150 nsew default input
rlabel metal2 s 1398 22320 1454 22800 6 top_left_grid_pin_44_
port 151 nsew default input
rlabel metal2 s 1858 22320 1914 22800 6 top_left_grid_pin_45_
port 152 nsew default input
rlabel metal2 s 2226 22320 2282 22800 6 top_left_grid_pin_46_
port 153 nsew default input
rlabel metal2 s 2686 22320 2742 22800 6 top_left_grid_pin_47_
port 154 nsew default input
rlabel metal2 s 3146 22320 3202 22800 6 top_left_grid_pin_48_
port 155 nsew default input
rlabel metal2 s 3514 22320 3570 22800 6 top_left_grid_pin_49_
port 156 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 157 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 158 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
