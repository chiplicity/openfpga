* NGSPICE file created from grid_clb.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxbp_1 abstract view
.subckt sky130_fd_sc_hd__dfxbp_1 D Q Q_N CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__sdfxbp_1 abstract view
.subckt sky130_fd_sc_hd__sdfxbp_1 D Q Q_N SCD SCE CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

.subckt grid_clb Test_en bottom_width_0_height_0__pin_16_ bottom_width_0_height_0__pin_17_
+ bottom_width_0_height_0__pin_18_ bottom_width_0_height_0__pin_19_ bottom_width_0_height_0__pin_20_
+ bottom_width_0_height_0__pin_21_ bottom_width_0_height_0__pin_22_ bottom_width_0_height_0__pin_23_
+ bottom_width_0_height_0__pin_24_ bottom_width_0_height_0__pin_25_ bottom_width_0_height_0__pin_26_
+ bottom_width_0_height_0__pin_27_ bottom_width_0_height_0__pin_28_ bottom_width_0_height_0__pin_29_
+ bottom_width_0_height_0__pin_30_ bottom_width_0_height_0__pin_31_ bottom_width_0_height_0__pin_42_lower
+ bottom_width_0_height_0__pin_42_upper bottom_width_0_height_0__pin_43_lower bottom_width_0_height_0__pin_43_upper
+ bottom_width_0_height_0__pin_44_lower bottom_width_0_height_0__pin_44_upper bottom_width_0_height_0__pin_45_lower
+ bottom_width_0_height_0__pin_45_upper bottom_width_0_height_0__pin_46_lower bottom_width_0_height_0__pin_46_upper
+ bottom_width_0_height_0__pin_47_lower bottom_width_0_height_0__pin_47_upper bottom_width_0_height_0__pin_48_lower
+ bottom_width_0_height_0__pin_48_upper bottom_width_0_height_0__pin_49_lower bottom_width_0_height_0__pin_49_upper
+ bottom_width_0_height_0__pin_50_ bottom_width_0_height_0__pin_51_ ccff_head ccff_tail
+ clk left_width_0_height_0__pin_52_ prog_clk right_width_0_height_0__pin_0_ right_width_0_height_0__pin_10_
+ right_width_0_height_0__pin_11_ right_width_0_height_0__pin_12_ right_width_0_height_0__pin_13_
+ right_width_0_height_0__pin_14_ right_width_0_height_0__pin_15_ right_width_0_height_0__pin_1_
+ right_width_0_height_0__pin_2_ right_width_0_height_0__pin_34_lower right_width_0_height_0__pin_34_upper
+ right_width_0_height_0__pin_35_lower right_width_0_height_0__pin_35_upper right_width_0_height_0__pin_36_lower
+ right_width_0_height_0__pin_36_upper right_width_0_height_0__pin_37_lower right_width_0_height_0__pin_37_upper
+ right_width_0_height_0__pin_38_lower right_width_0_height_0__pin_38_upper right_width_0_height_0__pin_39_lower
+ right_width_0_height_0__pin_39_upper right_width_0_height_0__pin_3_ right_width_0_height_0__pin_40_lower
+ right_width_0_height_0__pin_40_upper right_width_0_height_0__pin_41_lower right_width_0_height_0__pin_41_upper
+ right_width_0_height_0__pin_4_ right_width_0_height_0__pin_5_ right_width_0_height_0__pin_6_
+ right_width_0_height_0__pin_7_ right_width_0_height_0__pin_8_ right_width_0_height_0__pin_9_
+ top_width_0_height_0__pin_32_ top_width_0_height_0__pin_33_ VPWR VGND
XFILLER_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _62_/HI
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _36_/HI
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_43_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_41_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_66_ bottom_width_0_height_0__pin_44_lower bottom_width_0_height_0__pin_44_upper
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ right_width_0_height_0__pin_0_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_49_ _49_/HI _49_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
+ ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _35_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ right_width_0_height_0__pin_8_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_5_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_65_ bottom_width_0_height_0__pin_43_lower bottom_width_0_height_0__pin_43_upper
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ bottom_width_0_height_0__pin_31_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ bottom_width_0_height_0__pin_18_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_48_ _48_/HI _48_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_52_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ccff_tail
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_5_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_64_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_64_ bottom_width_0_height_0__pin_42_lower bottom_width_0_height_0__pin_42_upper
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_64_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XFILLER_55_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _61_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ bottom_width_0_height_0__pin_17_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_47_ _47_/HI _47_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ right_width_0_height_0__pin_5_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _48_/HI
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_49_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_80_ right_width_0_height_0__pin_41_lower right_width_0_height_0__pin_41_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_63_ _63_/HI _63_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ bottom_width_0_height_0__pin_16_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_46_ _46_/HI _46_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _47_/HI ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _56_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _63_/HI ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ bottom_width_0_height_0__pin_27_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_53_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_62_ _62_/HI _62_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _57_/HI
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_36_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_45_ _45_/HI _45_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_46_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _55_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ right_width_0_height_0__pin_2_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_clk_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_16_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ right_width_0_height_0__pin_3_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ bottom_width_0_height_0__pin_30_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_61_ _61_/HI _61_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_44_ _44_/HI _44_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_64_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _45_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XFILLER_43_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_0_0_clk_A clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_60_ _60_/HI _60_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ bottom_width_0_height_0__pin_24_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_43_ _43_/HI _43_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_60_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _40_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _38_/HI
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _37_/HI
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_42_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_42_ _42_/HI _42_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
+ ccff_head ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ bottom_width_0_height_0__pin_19_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ right_width_0_height_0__pin_6_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ bottom_width_0_height_0__pin_21_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_41_ _41_/HI _41_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_42_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__64__A bottom_width_0_height_0__pin_42_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_45_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__72__A bottom_width_0_height_0__pin_50_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ right_width_0_height_0__pin_15_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ bottom_width_0_height_0__pin_50_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ right_width_0_height_0__pin_5_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__67__A bottom_width_0_height_0__pin_45_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_40_ _40_/HI _40_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__80__A right_width_0_height_0__pin_41_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__75__A right_width_0_height_0__pin_36_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XFILLER_24_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _60_/HI
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_39_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_50_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ right_width_0_height_0__pin_4_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ bottom_width_0_height_0__pin_18_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _49_/HI
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_48_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_16_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _43_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__78__A right_width_0_height_0__pin_39_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ top_width_0_height_0__pin_33_ Test_en clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _57_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ bottom_width_0_height_0__pin_22_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_50_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ right_width_0_height_0__pin_12_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_64_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ bottom_width_0_height_0__pin_50_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_42_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _52_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ bottom_width_0_height_0__pin_21_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _35_/HI ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _40_/HI
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_45_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_46_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ bottom_width_0_height_0__pin_20_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_1_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ right_width_0_height_0__pin_9_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _51_/HI ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_79_ right_width_0_height_0__pin_40_lower right_width_0_height_0__pin_40_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _41_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_44_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ right_width_0_height_0__pin_3_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _63_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _46_/HI
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _58_/HI
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_36_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ bottom_width_0_height_0__pin_31_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_78_ right_width_0_height_0__pin_39_lower right_width_0_height_0__pin_39_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_51_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ right_width_0_height_0__pin_7_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XFILLER_21_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _36_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ right_width_0_height_0__pin_6_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_44_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_77_ right_width_0_height_0__pin_38_lower right_width_0_height_0__pin_38_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ right_width_0_height_0__pin_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_76_ right_width_0_height_0__pin_37_lower right_width_0_height_0__pin_37_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ bottom_width_0_height_0__pin_28_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_59_ _59_/HI _59_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _61_/HI
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_38_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_75_ right_width_0_height_0__pin_36_lower right_width_0_height_0__pin_36_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ bottom_width_0_height_0__pin_23_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _51_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_58_ _58_/HI _58_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ right_width_0_height_0__pin_10_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_52_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ bottom_width_0_height_0__pin_25_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_74_ right_width_0_height_0__pin_35_lower right_width_0_height_0__pin_35_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _53_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_1_0_clk clkbuf_0_clk/X clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_57_ _57_/HI _57_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ right_width_0_height_0__pin_9_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_40_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_4_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ bottom_width_0_height_0__pin_19_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_73_ right_width_0_height_0__pin_34_lower right_width_0_height_0__pin_34_upper VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_14_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_64_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_56_ _56_/HI _56_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ right_width_0_height_0__pin_8_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_39_ _39_/HI _39_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_52_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _52_/HI
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_35_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0_clk clkbuf_0_clk/X clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_43_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _41_/HI
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_44_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ bottom_width_0_height_0__pin_22_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _54_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__70__A bottom_width_0_height_0__pin_48_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_72_ bottom_width_0_height_0__pin_50_ bottom_width_0_height_0__pin_51_ VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__65__A bottom_width_0_height_0__pin_43_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ bottom_width_0_height_0__pin_26_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_55_ _55_/HI _55_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_38_ _38_/HI _38_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__73__A right_width_0_height_0__pin_34_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__68__A bottom_width_0_height_0__pin_46_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _34_/HI
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_53_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_71_ bottom_width_0_height_0__pin_49_lower bottom_width_0_height_0__pin_49_upper
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ bottom_width_0_height_0__pin_16_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _39_/HI ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ bottom_width_0_height_0__pin_25_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_54_ _54_/HI _54_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _58_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _37_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__76__A right_width_0_height_0__pin_37_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_37_ _37_/HI _37_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _55_/HI ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__79__A right_width_0_height_0__pin_40_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_70_ bottom_width_0_height_0__pin_48_lower bottom_width_0_height_0__pin_48_upper
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ bottom_width_0_height_0__pin_24_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_53_ _53_/HI _53_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _32_/HI
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_41_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_36_ _36_/HI _36_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _62_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _32_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ right_width_0_height_0__pin_13_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _39_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_52_ _52_/HI _52_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_35_ _35_/HI _35_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ right_width_0_height_0__pin_7_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _34_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ right_width_0_height_0__pin_11_ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XFILLER_41_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_55_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ top_width_0_height_0__pin_33_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_51_ _51_/HI _51_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_1_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_34_ _34_/HI _34_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ right_width_0_height_0__pin_10_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_4_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_50_ _50_/HI _50_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _38_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _44_/HI
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_47_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_33_ _33_/HI _33_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_45_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _48_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ right_width_0_height_0__pin_4_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_32_ _32_/HI _32_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_60_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _42_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _59_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _53_/HI
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_34_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ bottom_width_0_height_0__pin_27_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ right_width_0_height_0__pin_14_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_49_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__CLK
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_45_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ right_width_0_height_0__pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ right_width_0_height_0__pin_13_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _46_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _42_/HI
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _54_/HI
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ bottom_width_0_height_0__pin_29_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4__A
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ right_width_0_height_0__pin_12_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ bottom_width_0_height_0__pin_23_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A0
+ _50_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_51_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _33_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XFILLER_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_ top_width_0_height_0__pin_32_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _33_/HI
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ right_width_0_height_0__pin_40_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ bottom_width_0_height_0__pin_30_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _43_/HI ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ bottom_width_0_height_0__pin_26_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
+ _59_/HI ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ top_width_0_height_0__pin_32_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _60_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ bottom_width_0_height_0__pin_29_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0__A
+ bottom_width_0_height_0__pin_20_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_41_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5__A
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_15_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_61_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
+ bottom_width_0_height_0__pin_28_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_61_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_1_1_0_clk_A clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__71__A bottom_width_0_height_0__pin_49_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_10_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ bottom_width_0_height_0__pin_50_ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ Test_en clkbuf_1_1_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__66__A bottom_width_0_height_0__pin_44_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_ _56_/HI
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ right_width_0_height_0__pin_37_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A0
+ _47_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_14_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_69_ bottom_width_0_height_0__pin_47_lower bottom_width_0_height_0__pin_47_upper
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_ _45_/HI
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ bottom_width_0_height_0__pin_46_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A0
+ _49_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__74__A right_width_0_height_0__pin_35_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_0.sky130_fd_sc_hd__sdfxbp_1_0_/Q_N
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 Test_en
+ clkbuf_1_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__sdfxbp_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__69__A bottom_width_0_height_0__pin_47_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
+ bottom_width_0_height_0__pin_17_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_16__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__77__A right_width_0_height_0__pin_38_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_13_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_6__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_68_ bottom_width_0_height_0__pin_46_lower bottom_width_0_height_0__pin_46_upper
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ right_width_0_height_0__pin_15_ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__or2_1
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_4__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
+ right_width_0_height_0__pin_2_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_3_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A0
+ _44_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
+ right_width_0_height_0__pin_11_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9__D
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_9_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/S
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A1 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_fabric_out_1.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCE
+ Test_en VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7__D
+ ltile_clb_mode_0.ltile_clb_fle_4.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_md_fle_mp_fab_md_ff_1.sky130_fd_sc_hd__sdfxbp_1_0__SCD
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_5__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_12_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A1
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_7_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_67_ bottom_width_0_height_0__pin_45_lower bottom_width_0_height_0__pin_45_upper
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/A0 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxbp_1_1__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.mux_fabric_out_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
+ right_width_0_height_0__pin_1_ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1__S
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5__A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6__A
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_34_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0__S
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__S
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_15__D
+ ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l2_in_0__A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.mux_fabric_out_0.mux_l1_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_ _50_/HI
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l1_in_0_/X ccff_tail
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.mux_ff_0_D_0.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_3.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
+ right_width_0_height_0__pin_14_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_/X
+ ltile_clb_mode_0.ltile_clb_fle_1.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A0
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/A1
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_5.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_11__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8__D
+ ltile_clb_mode_0.ltile_clb_fle_7.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1__A0
+ ltile_clb_mode_0.ltile_clb_fle_2.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_/A0
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.sky130_fd_sc_hd__dfxbp_1_8_/Q_N
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_ltile_clb_mode_0.ltile_clb_fle_0.ltile_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
+ prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A0
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/A1
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_/X
+ ltile_clb_mode_0.ltile_clb_fle_6.ltile_fabric_0.ltile_clb_frac_logic_0.ltile_clb_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
.ends

