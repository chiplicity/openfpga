* NGSPICE file created from sb_3__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt sb_3__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ bottom_right_grid_pin_13_ bottom_right_grid_pin_15_
+ bottom_right_grid_pin_1_ bottom_right_grid_pin_3_ bottom_right_grid_pin_5_ bottom_right_grid_pin_7_
+ bottom_right_grid_pin_9_ chanx_left_in[0] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_out[0] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4]
+ chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chany_bottom_in[0]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] data_in enable left_bottom_grid_pin_12_
+ left_top_grid_pin_11_ left_top_grid_pin_13_ left_top_grid_pin_15_ left_top_grid_pin_1_
+ left_top_grid_pin_3_ left_top_grid_pin_5_ left_top_grid_pin_7_ left_top_grid_pin_9_
+ vpwr vgnd
XFILLER_22_166 vgnd vpwr scs8hd_decap_12
XFILLER_22_144 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_111 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_166 vpwr vgnd scs8hd_fill_2
XFILLER_3_34 vpwr vgnd scs8hd_fill_2
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _225_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_21 vpwr vgnd scs8hd_fill_2
XFILLER_12_43 vpwr vgnd scs8hd_fill_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XANTENNA__108__B enable vgnd vpwr scs8hd_diode_2
XFILLER_5_162 vgnd vpwr scs8hd_decap_4
XANTENNA__124__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _190_/A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_53 vgnd vpwr scs8hd_decap_4
XFILLER_23_42 vpwr vgnd scs8hd_fill_2
X_131_ _135_/A _130_/X _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_165 vgnd vpwr scs8hd_decap_8
XFILLER_2_154 vpwr vgnd scs8hd_fill_2
XFILLER_2_110 vgnd vpwr scs8hd_decap_3
XANTENNA__110__C _100_/X vgnd vpwr scs8hd_diode_2
XANTENNA__119__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_22 vgnd vpwr scs8hd_decap_3
XFILLER_9_88 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _173_/Y mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_34_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
X_114_ _163_/B _130_/B vgnd vpwr scs8hd_buf_1
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
XFILLER_39_19 vpwr vgnd scs8hd_fill_2
XFILLER_29_74 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _223_/HI _194_/Y mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_87 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__116__B _115_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__132__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_53 vgnd vpwr scs8hd_decap_8
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _187_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XANTENNA__127__A _127_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_120 vpwr vgnd scs8hd_fill_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vgnd vpwr scs8hd_decap_12
XFILLER_22_178 vgnd vpwr scs8hd_decap_12
XFILLER_9_105 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_3_79 vpwr vgnd scs8hd_fill_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XFILLER_3_13 vgnd vpwr scs8hd_decap_4
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_10_104 vpwr vgnd scs8hd_fill_2
XFILLER_10_137 vpwr vgnd scs8hd_fill_2
XFILLER_12_88 vgnd vpwr scs8hd_decap_4
XANTENNA__230__A _230_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.tap_buf4_0_.scs8hd_inv_1 mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _206_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XANTENNA__124__B _124_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _173_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__140__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_23_21 vgnd vpwr scs8hd_decap_4
X_130_ _130_/A _130_/B _130_/C _169_/A _130_/X vgnd vpwr scs8hd_or4_4
XFILLER_2_122 vpwr vgnd scs8hd_fill_2
XANTENNA__110__D _110_/D vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__119__B _118_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__135__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_5.tap_buf4_0_.scs8hd_inv_1 mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _232_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_76 vpwr vgnd scs8hd_fill_2
XFILLER_7_214 vgnd vpwr scs8hd_fill_1
XFILLER_7_225 vpwr vgnd scs8hd_fill_2
XFILLER_7_236 vgnd vpwr scs8hd_decap_8
X_113_ address[2] _163_/B vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
XFILLER_15_7 vgnd vpwr scs8hd_fill_1
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_20_66 vgnd vpwr scs8hd_decap_4
XFILLER_29_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_53 vgnd vpwr scs8hd_decap_8
XFILLER_29_42 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_13 vpwr vgnd scs8hd_fill_2
XFILLER_6_24 vpwr vgnd scs8hd_fill_2
XFILLER_6_35 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _193_/A mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
Xmem_left_track_5.LATCH_1_.latch data_in _194_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_77 vpwr vgnd scs8hd_fill_2
XFILLER_15_88 vpwr vgnd scs8hd_fill_2
XFILLER_31_98 vgnd vpwr scs8hd_decap_12
XANTENNA__233__A _233_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_253 vpwr vgnd scs8hd_fill_2
XFILLER_31_135 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _175_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__127__B _127_/B vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_257 vgnd vpwr scs8hd_decap_12
XFILLER_30_190 vgnd vpwr scs8hd_decap_12
XFILLER_26_10 vpwr vgnd scs8hd_fill_2
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_87 vgnd vpwr scs8hd_decap_4
XFILLER_26_43 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _235_/A vgnd vpwr scs8hd_inv_1
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A address[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _197_/Y mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_175 vgnd vpwr scs8hd_decap_6
XFILLER_5_197 vpwr vgnd scs8hd_fill_2
XANTENNA__140__B _143_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XFILLER_3_3 vgnd vpwr scs8hd_fill_1
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
XANTENNA__241__A _241_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XANTENNA__135__B _135_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XFILLER_18_88 vpwr vgnd scs8hd_fill_2
X_112_ _128_/A _110_/X _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__236__A _236_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_248 vpwr vgnd scs8hd_fill_2
XANTENNA__146__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_270 vgnd vpwr scs8hd_decap_4
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_20_12 vpwr vgnd scs8hd_fill_2
XFILLER_20_23 vgnd vpwr scs8hd_decap_6
XFILLER_29_98 vgnd vpwr scs8hd_decap_12
XFILLER_28_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_6 vgnd vpwr scs8hd_decap_4
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_130 vgnd vpwr scs8hd_decap_12
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XFILLER_15_23 vpwr vgnd scs8hd_fill_2
XFILLER_15_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_31_22 vpwr vgnd scs8hd_fill_2
XFILLER_31_11 vpwr vgnd scs8hd_fill_2
XFILLER_0_265 vpwr vgnd scs8hd_fill_2
XFILLER_0_243 vgnd vpwr scs8hd_decap_4
XFILLER_16_133 vgnd vpwr scs8hd_decap_8
XFILLER_16_144 vgnd vpwr scs8hd_decap_8
XFILLER_31_147 vgnd vpwr scs8hd_decap_12
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _143_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_66 vpwr vgnd scs8hd_fill_2
XFILLER_26_55 vgnd vpwr scs8hd_decap_8
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__138__B _166_/D vgnd vpwr scs8hd_diode_2
XFILLER_8_184 vpwr vgnd scs8hd_fill_2
XANTENNA__154__A _170_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_15_ mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_68 vgnd vpwr scs8hd_fill_1
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XFILLER_38_7 vgnd vpwr scs8hd_decap_12
Xmem_left_track_15.LATCH_0_.latch data_in _205_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_132 vgnd vpwr scs8hd_decap_4
XFILLER_5_143 vpwr vgnd scs8hd_fill_2
XANTENNA__140__C _139_/X vgnd vpwr scs8hd_diode_2
XANTENNA__149__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _188_/A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_220 vgnd vpwr scs8hd_decap_12
XFILLER_23_78 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_102 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_14 vpwr vgnd scs8hd_fill_2
XFILLER_9_36 vpwr vgnd scs8hd_fill_2
X_188_ _188_/A _188_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__151__B _149_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_18_23 vpwr vgnd scs8hd_fill_2
XFILLER_18_56 vgnd vpwr scs8hd_fill_1
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
X_111_ _127_/A _110_/X _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
XANTENNA__146__B _130_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_1_92 vpwr vgnd scs8hd_fill_2
XFILLER_20_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_263 vpwr vgnd scs8hd_fill_2
XFILLER_3_252 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_142 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_0_200 vpwr vgnd scs8hd_fill_2
XFILLER_31_159 vgnd vpwr scs8hd_decap_12
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__143__C _139_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _222_/HI _192_/Y mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_3
XFILLER_22_104 vpwr vgnd scs8hd_fill_2
XFILLER_7_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _207_/Y vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in _190_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XFILLER_13_115 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_38 vgnd vpwr scs8hd_decap_4
XANTENNA__154__B _156_/B vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _110_/D vgnd vpwr scs8hd_diode_2
XFILLER_12_25 vpwr vgnd scs8hd_fill_2
XFILLER_12_47 vpwr vgnd scs8hd_fill_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_166 vgnd vpwr scs8hd_fill_1
XANTENNA__140__D _103_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _130_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_4_81 vgnd vpwr scs8hd_decap_4
XFILLER_23_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_57 vgnd vpwr scs8hd_fill_1
Xmux_left_track_13.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_13_ mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A _187_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_180 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_202 vgnd vpwr scs8hd_decap_12
XFILLER_18_46 vpwr vgnd scs8hd_fill_2
XFILLER_18_68 vpwr vgnd scs8hd_fill_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _118_/A _143_/B _100_/X _110_/D _110_/X vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _186_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_202 vgnd vpwr scs8hd_decap_12
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
XFILLER_7_217 vgnd vpwr scs8hd_fill_1
X_239_ _239_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__146__C _139_/X vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _161_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XFILLER_1_71 vpwr vgnd scs8hd_fill_2
XFILLER_29_34 vgnd vpwr scs8hd_decap_4
XFILLER_29_12 vpwr vgnd scs8hd_fill_2
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
XFILLER_3_275 vpwr vgnd scs8hd_fill_2
XFILLER_13_7 vgnd vpwr scs8hd_decap_3
XFILLER_19_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__157__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_0_212 vgnd vpwr scs8hd_decap_3
XFILLER_24_190 vgnd vpwr scs8hd_decap_12
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_157 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _172_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__143__D _109_/A vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A _169_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _191_/A mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_26_35 vgnd vpwr scs8hd_decap_8
XFILLER_13_149 vgnd vpwr scs8hd_decap_6
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_171 vgnd vpwr scs8hd_decap_12
XFILLER_9_109 vgnd vpwr scs8hd_decap_3
XANTENNA__170__B _169_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_131 vgnd vpwr scs8hd_decap_4
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XFILLER_10_108 vpwr vgnd scs8hd_fill_2
XFILLER_10_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
XANTENNA__149__C _139_/X vgnd vpwr scs8hd_diode_2
XANTENNA__165__B _165_/B vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_36 vgnd vpwr scs8hd_decap_4
Xmux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _195_/Y mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_2_126 vpwr vgnd scs8hd_fill_2
X_186_ _186_/A _186_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_11.LATCH_0_.latch data_in _201_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XFILLER_11_214 vgnd vpwr scs8hd_decap_12
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd
+ vpwr scs8hd_diode_2
X_238_ _238_/A chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA__146__D _103_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_11.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_11_ mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_169_ _169_/A _169_/B _169_/C _169_/Y vgnd vpwr scs8hd_nor3_4
Xmem_bottom_track_7.LATCH_0_.latch data_in _179_/A _120_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_46 vgnd vpwr scs8hd_decap_4
XFILLER_28_166 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_17 vgnd vpwr scs8hd_decap_4
XFILLER_6_28 vgnd vpwr scs8hd_decap_3
XFILLER_6_39 vgnd vpwr scs8hd_decap_4
XFILLER_3_243 vgnd vpwr scs8hd_fill_1
XFILLER_19_166 vgnd vpwr scs8hd_decap_12
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XANTENNA__157__C _139_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_257 vgnd vpwr scs8hd_decap_4
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_169 vgnd vpwr scs8hd_decap_12
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _169_/B vgnd vpwr scs8hd_diode_2
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_60 vgnd vpwr scs8hd_fill_1
XFILLER_12_150 vgnd vpwr scs8hd_decap_3
XFILLER_8_165 vgnd vpwr scs8hd_decap_8
XANTENNA__170__C _170_/C vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_113 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__149__D _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XFILLER_14_212 vpwr vgnd scs8hd_fill_2
X_185_ _185_/A _185_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_92 vgnd vpwr scs8hd_fill_1
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_226 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _186_/A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_237_ _237_/A chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
X_168_ _169_/A _169_/B _170_/C _168_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_3
X_099_ address[4] address[5] _130_/C vgnd vpwr scs8hd_or2_4
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_49 vpwr vgnd scs8hd_fill_2
XFILLER_28_178 vgnd vpwr scs8hd_decap_12
XANTENNA__097__A address[3] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_15.LATCH_0_.latch data_in _187_/A _136_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_71 vpwr vgnd scs8hd_fill_2
XFILLER_10_93 vpwr vgnd scs8hd_fill_2
XFILLER_19_178 vgnd vpwr scs8hd_decap_4
XANTENNA__157__D _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_159 vgnd vpwr scs8hd_decap_12
XFILLER_15_38 vpwr vgnd scs8hd_fill_2
XFILLER_0_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
XFILLER_16_104 vgnd vpwr scs8hd_decap_3
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_5.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__168__C _170_/C vgnd vpwr scs8hd_diode_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_19 vpwr vgnd scs8hd_fill_2
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_188 vgnd vpwr scs8hd_decap_4
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _217_/HI _190_/Y mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_147 vgnd vpwr scs8hd_decap_4
XFILLER_5_169 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _241_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XFILLER_2_139 vgnd vpwr scs8hd_decap_4
XFILLER_2_106 vpwr vgnd scs8hd_fill_2
XFILLER_9_18 vpwr vgnd scs8hd_fill_2
X_184_ _184_/A _184_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_71 vgnd vpwr scs8hd_decap_4
XFILLER_1_172 vpwr vgnd scs8hd_fill_2
XFILLER_9_261 vgnd vpwr scs8hd_decap_12
XFILLER_20_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vpwr vgnd scs8hd_fill_2
XFILLER_11_238 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_098_ address[2] _143_/B vgnd vpwr scs8hd_buf_1
X_236_ _236_/A chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_10_271 vgnd vpwr scs8hd_decap_4
X_167_ _166_/X _169_/B vgnd vpwr scs8hd_buf_1
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _206_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XFILLER_3_212 vpwr vgnd scs8hd_fill_2
XFILLER_3_267 vgnd vpwr scs8hd_decap_8
XFILLER_10_61 vpwr vgnd scs8hd_fill_2
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XFILLER_18_190 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_3.LATCH_0_.latch data_in _175_/A _112_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_116 vpwr vgnd scs8hd_fill_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_93 vpwr vgnd scs8hd_fill_2
XFILLER_21_71 vpwr vgnd scs8hd_fill_2
XFILLER_39_208 vgnd vpwr scs8hd_decap_12
XFILLER_22_108 vgnd vpwr scs8hd_decap_12
XPHY_2 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _189_/A mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_160 vpwr vgnd scs8hd_fill_2
XFILLER_15_171 vgnd vpwr scs8hd_decap_12
XFILLER_30_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_73 vpwr vgnd scs8hd_fill_2
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_21_196 vgnd vpwr scs8hd_decap_12
XFILLER_13_119 vgnd vpwr scs8hd_decap_3
XFILLER_16_71 vgnd vpwr scs8hd_decap_4
XFILLER_16_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_123 vpwr vgnd scs8hd_fill_2
XFILLER_8_145 vgnd vpwr scs8hd_decap_8
XFILLER_12_163 vgnd vpwr scs8hd_decap_8
XFILLER_12_174 vgnd vpwr scs8hd_decap_8
XFILLER_12_185 vgnd vpwr scs8hd_decap_8
XFILLER_12_196 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_15.INVTX1_1_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_81 vgnd vpwr scs8hd_decap_12
XFILLER_27_70 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _234_/A vgnd vpwr scs8hd_inv_1
XFILLER_4_85 vgnd vpwr scs8hd_fill_1
XFILLER_4_52 vgnd vpwr scs8hd_fill_1
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_23_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _175_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_9_ mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_183_ _183_/A _183_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_195 vpwr vgnd scs8hd_fill_2
XFILLER_1_184 vpwr vgnd scs8hd_fill_2
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XFILLER_9_273 vgnd vpwr scs8hd_decap_4
XFILLER_20_239 vgnd vpwr scs8hd_decap_12
XFILLER_1_6 vpwr vgnd scs8hd_fill_2
XFILLER_24_93 vgnd vpwr scs8hd_decap_12
XFILLER_24_71 vpwr vgnd scs8hd_fill_2
X_235_ _235_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
Xmux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _193_/Y mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_097_ address[3] _118_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_166_ address[3] address[2] address[4] _166_/D _166_/X vgnd vpwr scs8hd_or4_4
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
XFILLER_1_31 vpwr vgnd scs8hd_fill_2
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_1_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_38 vgnd vpwr scs8hd_fill_1
XFILLER_29_16 vpwr vgnd scs8hd_fill_2
XFILLER_3_235 vgnd vpwr scs8hd_decap_8
XFILLER_10_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
XFILLER_19_93 vpwr vgnd scs8hd_fill_2
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
X_149_ address[3] _130_/B _139_/X _109_/A _149_/X vgnd vpwr scs8hd_or4_4
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_106 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _237_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_227 vgnd vpwr scs8hd_decap_8
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_track_11.LATCH_0_.latch data_in _183_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_52 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _177_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_102 vpwr vgnd scs8hd_fill_2
XFILLER_12_142 vgnd vpwr scs8hd_decap_8
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_135 vgnd vpwr scs8hd_fill_1
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_5_138 vpwr vgnd scs8hd_fill_2
XFILLER_27_93 vgnd vpwr scs8hd_decap_12
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_20 vgnd vpwr scs8hd_decap_4
XFILLER_4_182 vpwr vgnd scs8hd_fill_2
XFILLER_4_64 vpwr vgnd scs8hd_fill_2
XFILLER_14_204 vgnd vpwr scs8hd_decap_8
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_182_ _182_/A _182_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_40 vpwr vgnd scs8hd_fill_2
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_13_95 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_13.INVTX1_1_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__100__A _130_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_230 vgnd vpwr scs8hd_decap_12
X_234_ _234_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
X_165_ _169_/C _165_/B _165_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XFILLER_34_7 vgnd vpwr scs8hd_decap_8
X_096_ _095_/Y _127_/A vgnd vpwr scs8hd_buf_1
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
XFILLER_1_10 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_7_ mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_15.LATCH_1_.latch data_in _204_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_41 vgnd vpwr scs8hd_decap_3
XFILLER_19_126 vpwr vgnd scs8hd_fill_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _184_/A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_148_ _133_/A _148_/B _148_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd vpwr
+ scs8hd_diode_2
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
XFILLER_25_3 vpwr vgnd scs8hd_fill_2
XFILLER_25_118 vgnd vpwr scs8hd_decap_4
XFILLER_15_19 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_29 vgnd vpwr scs8hd_decap_12
XFILLER_31_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_239 vpwr vgnd scs8hd_fill_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_154 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_110 vpwr vgnd scs8hd_fill_2
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XFILLER_16_51 vgnd vpwr scs8hd_decap_6
XFILLER_16_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _188_/Y mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_43 vgnd vpwr scs8hd_decap_3
XFILLER_4_150 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
X_181_ _181_/A _181_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_9_242 vpwr vgnd scs8hd_fill_2
XFILLER_34_18 vgnd vpwr scs8hd_decap_12
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
X_233_ _233_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_24_84 vgnd vpwr scs8hd_decap_8
X_164_ _170_/C _165_/B _164_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
X_095_ address[0] _095_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_88 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _127_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_29_29 vgnd vpwr scs8hd_decap_3
XFILLER_28_105 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_11.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_259 vpwr vgnd scs8hd_fill_2
XFILLER_3_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
X_147_ _135_/A _148_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_270 vgnd vpwr scs8hd_decap_4
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_5_ mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_141 vgnd vpwr scs8hd_decap_12
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_30 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_30_166 vgnd vpwr scs8hd_decap_12
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
XFILLER_7_65 vpwr vgnd scs8hd_fill_2
XFILLER_7_87 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _206_/A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _187_/A mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_62 vgnd vpwr scs8hd_decap_4
XFILLER_17_269 vgnd vpwr scs8hd_decap_8
XFILLER_4_88 vpwr vgnd scs8hd_fill_2
XANTENNA__114__A _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _208_/HI vgnd vpwr
+ scs8hd_diode_2
X_180_ _180_/A _180_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_53 vgnd vpwr scs8hd_decap_6
XFILLER_1_176 vgnd vpwr scs8hd_decap_4
XFILLER_1_154 vgnd vpwr scs8hd_decap_3
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
X_232_ _232_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_6_224 vgnd vpwr scs8hd_decap_8
XFILLER_6_235 vgnd vpwr scs8hd_decap_8
XFILLER_6_246 vgnd vpwr scs8hd_decap_12
X_163_ _163_/A _163_/B _163_/C _109_/A _165_/B vgnd vpwr scs8hd_or4_4
XFILLER_1_23 vpwr vgnd scs8hd_fill_2
XANTENNA__111__B _110_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_117 vgnd vpwr scs8hd_decap_12
XFILLER_3_216 vpwr vgnd scs8hd_fill_2
XFILLER_10_10 vpwr vgnd scs8hd_fill_2
XFILLER_10_65 vgnd vpwr scs8hd_decap_4
XFILLER_19_41 vgnd vpwr scs8hd_fill_1
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
X_146_ address[3] _130_/B _139_/X _103_/A _148_/B vgnd vpwr scs8hd_or4_4
XANTENNA__122__A _163_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _191_/Y mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_208 vpwr vgnd scs8hd_fill_2
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_11.LATCH_1_.latch data_in _200_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_97 vpwr vgnd scs8hd_fill_2
XFILLER_21_75 vgnd vpwr scs8hd_decap_3
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_30_178 vgnd vpwr scs8hd_decap_12
XANTENNA__117__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_33 vpwr vgnd scs8hd_fill_2
XFILLER_7_77 vgnd vpwr scs8hd_fill_1
X_129_ _095_/Y _135_/A vgnd vpwr scs8hd_buf_1
XFILLER_21_123 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _180_/A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_7.LATCH_1_.latch data_in _178_/A _119_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_30 vgnd vpwr scs8hd_fill_1
XFILLER_8_127 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_3_ mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_27_74 vgnd vpwr scs8hd_decap_4
Xmem_left_track_7.LATCH_0_.latch data_in _197_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__130__A _130_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_251 vgnd vpwr scs8hd_decap_12
XFILLER_1_199 vpwr vgnd scs8hd_fill_2
XFILLER_1_111 vpwr vgnd scs8hd_fill_2
XFILLER_8_3 vpwr vgnd scs8hd_fill_2
XANTENNA__125__A _128_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_231_ _231_/A chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_24_53 vgnd vpwr scs8hd_decap_3
XFILLER_10_243 vgnd vpwr scs8hd_fill_1
X_162_ _169_/C _161_/B _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_258 vgnd vpwr scs8hd_decap_12
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_129 vgnd vpwr scs8hd_decap_12
XFILLER_10_88 vpwr vgnd scs8hd_fill_2
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vgnd vpwr scs8hd_decap_4
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_19_75 vgnd vpwr scs8hd_decap_3
XFILLER_19_97 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
X_145_ _133_/A _143_/X _145_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_7 vgnd vpwr scs8hd_decap_8
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _220_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_154 vgnd vpwr scs8hd_decap_12
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XANTENNA__117__B _115_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_56 vpwr vgnd scs8hd_fill_2
XANTENNA__133__A _133_/A vgnd vpwr scs8hd_diode_2
X_128_ _128_/A _127_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_135 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _182_/A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_12_135 vgnd vpwr scs8hd_decap_4
XFILLER_16_21 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_6
XFILLER_8_106 vpwr vgnd scs8hd_fill_2
XFILLER_20_190 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_15.LATCH_1_.latch data_in _186_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__128__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XFILLER_5_109 vpwr vgnd scs8hd_fill_2
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XFILLER_4_24 vgnd vpwr scs8hd_fill_1
XFILLER_4_131 vgnd vpwr scs8hd_decap_4
XFILLER_4_142 vgnd vpwr scs8hd_decap_8
XFILLER_4_68 vgnd vpwr scs8hd_decap_4
XFILLER_4_186 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_1_ mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__130__B _130_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_208 vgnd vpwr scs8hd_decap_12
XFILLER_22_263 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _186_/Y mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_77 vpwr vgnd scs8hd_fill_2
XFILLER_13_88 vgnd vpwr scs8hd_decap_4
XFILLER_13_99 vgnd vpwr scs8hd_fill_1
XANTENNA__231__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__125__B _124_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vpwr vgnd scs8hd_fill_2
XANTENNA__141__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_171 vgnd vpwr scs8hd_decap_12
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
X_230_ _230_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_8
XFILLER_24_21 vpwr vgnd scs8hd_fill_2
X_161_ _170_/C _161_/B _161_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XANTENNA__136__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XFILLER_3_229 vgnd vpwr scs8hd_decap_4
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
X_144_ _135_/A _143_/X _144_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_6 vpwr vgnd scs8hd_fill_2
XFILLER_18_130 vpwr vgnd scs8hd_fill_2
XFILLER_18_141 vgnd vpwr scs8hd_decap_12
XFILLER_24_166 vgnd vpwr scs8hd_decap_12
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__133__B _130_/X vgnd vpwr scs8hd_diode_2
X_127_ _127_/A _127_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _243_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_147 vgnd vpwr scs8hd_decap_12
XFILLER_21_114 vgnd vpwr scs8hd_decap_8
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_125 vgnd vpwr scs8hd_fill_1
XFILLER_16_77 vpwr vgnd scs8hd_fill_2
XFILLER_16_88 vpwr vgnd scs8hd_fill_2
XFILLER_16_99 vgnd vpwr scs8hd_decap_3
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA__234__A _234_/A vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_191 vpwr vgnd scs8hd_fill_2
XANTENNA__128__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_162 vpwr vgnd scs8hd_fill_2
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_32 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_3.LATCH_1_.latch data_in _174_/A _111_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_165 vpwr vgnd scs8hd_fill_2
XANTENNA__130__C _130_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _163_/C vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _204_/A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_23 vpwr vgnd scs8hd_fill_2
XFILLER_1_135 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _185_/A mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
XANTENNA__141__B _142_/B vgnd vpwr scs8hd_diode_2
Xmem_left_track_3.LATCH_0_.latch data_in _193_/A _148_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
X_160_ _163_/A _163_/B _163_/C _103_/A _161_/B vgnd vpwr scs8hd_or4_4
XANTENNA__242__A _242_/A vgnd vpwr scs8hd_diode_2
XANTENNA__136__B _135_/B vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _095_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_46 vpwr vgnd scs8hd_fill_2
XFILLER_19_22 vpwr vgnd scs8hd_fill_2
XFILLER_19_33 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__237__A _237_/A vgnd vpwr scs8hd_diode_2
X_143_ _118_/A _143_/B _139_/X _109_/A _143_/X vgnd vpwr scs8hd_or4_4
XFILLER_2_274 vgnd vpwr scs8hd_fill_1
XFILLER_2_241 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _189_/Y mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__147__A _135_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_24_178 vgnd vpwr scs8hd_decap_12
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_45 vpwr vgnd scs8hd_fill_2
XFILLER_21_23 vgnd vpwr scs8hd_fill_1
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vpwr vgnd scs8hd_fill_2
XFILLER_15_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_145 vpwr vgnd scs8hd_fill_2
XFILLER_15_156 vpwr vgnd scs8hd_fill_2
XFILLER_15_167 vpwr vgnd scs8hd_fill_2
XFILLER_7_69 vpwr vgnd scs8hd_fill_2
X_126_ _130_/A _143_/B _100_/X _110_/D _127_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_21_159 vgnd vpwr scs8hd_decap_12
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_119 vpwr vgnd scs8hd_fill_2
XFILLER_12_115 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__144__B _143_/X vgnd vpwr scs8hd_diode_2
XFILLER_11_170 vpwr vgnd scs8hd_fill_2
XANTENNA__160__A _163_/A vgnd vpwr scs8hd_diode_2
X_109_ _109_/A _110_/D vgnd vpwr scs8hd_buf_1
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_66 vgnd vpwr scs8hd_fill_1
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _178_/A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_48 vpwr vgnd scs8hd_fill_2
XFILLER_4_199 vgnd vpwr scs8hd_decap_12
XANTENNA__130__D _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_11.LATCH_1_.latch data_in _182_/A _127_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _177_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_24_67 vpwr vgnd scs8hd_fill_2
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_206 vgnd vpwr scs8hd_decap_8
XFILLER_10_213 vgnd vpwr scs8hd_fill_1
XFILLER_6_3 vgnd vpwr scs8hd_fill_1
XFILLER_1_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_11 vgnd vpwr scs8hd_decap_12
XFILLER_27_121 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _207_/A mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
X_142_ _133_/A _142_/B _142_/Y vgnd vpwr scs8hd_nor2_4
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.tap_buf4_0_.scs8hd_inv_1 mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _227_/A vgnd vpwr scs8hd_inv_1
XANTENNA__147__B _148_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_12
XANTENNA__163__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_113 vpwr vgnd scs8hd_fill_2
XFILLER_30_105 vgnd vpwr scs8hd_decap_12
X_125_ _128_/A _124_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_37 vpwr vgnd scs8hd_fill_2
XFILLER_30_7 vpwr vgnd scs8hd_fill_2
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA__158__A _170_/C vgnd vpwr scs8hd_diode_2
XFILLER_16_57 vgnd vpwr scs8hd_fill_1
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _179_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_7.tap_buf4_0_.scs8hd_inv_1 mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _231_/A vgnd vpwr scs8hd_inv_1
X_108_ address[1] enable _109_/A vgnd vpwr scs8hd_nand2_4
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_7_197 vpwr vgnd scs8hd_fill_2
XFILLER_11_182 vgnd vpwr scs8hd_fill_1
XANTENNA__160__B _163_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vpwr vgnd scs8hd_fill_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _183_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_208 vgnd vpwr scs8hd_decap_12
XFILLER_4_27 vpwr vgnd scs8hd_fill_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XANTENNA__171__A _110_/D vgnd vpwr scs8hd_diode_2
XFILLER_13_36 vpwr vgnd scs8hd_fill_2
XFILLER_1_159 vpwr vgnd scs8hd_fill_2
XFILLER_1_115 vpwr vgnd scs8hd_fill_2
XFILLER_8_7 vpwr vgnd scs8hd_fill_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _209_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_204 vpwr vgnd scs8hd_fill_2
XFILLER_9_215 vpwr vgnd scs8hd_fill_2
XFILLER_9_226 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__166__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_5_92 vpwr vgnd scs8hd_fill_2
XFILLER_39_196 vgnd vpwr scs8hd_decap_12
XFILLER_24_13 vpwr vgnd scs8hd_fill_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_247 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _184_/Y mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _181_/A mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_35_23 vgnd vpwr scs8hd_decap_12
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
X_141_ _135_/A _142_/B _141_/Y vgnd vpwr scs8hd_nor2_4
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
XFILLER_18_166 vgnd vpwr scs8hd_decap_12
XANTENNA__163__B _163_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _221_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_60 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_117 vgnd vpwr scs8hd_decap_12
X_124_ _127_/A _124_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_7 vgnd vpwr scs8hd_fill_1
XFILLER_11_91 vpwr vgnd scs8hd_fill_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
XANTENNA__158__B _158_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_180 vgnd vpwr scs8hd_decap_12
XFILLER_16_25 vpwr vgnd scs8hd_fill_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XFILLER_12_139 vgnd vpwr scs8hd_fill_1
X_107_ _128_/A _104_/X _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_132 vpwr vgnd scs8hd_fill_2
XFILLER_7_143 vgnd vpwr scs8hd_decap_4
XFILLER_14_3 vpwr vgnd scs8hd_fill_2
XANTENNA__160__C _163_/C vgnd vpwr scs8hd_diode_2
XANTENNA__169__A _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vgnd vpwr scs8hd_decap_4
XFILLER_25_220 vgnd vpwr scs8hd_decap_12
XFILLER_4_113 vgnd vpwr scs8hd_decap_3
XFILLER_4_102 vpwr vgnd scs8hd_fill_2
XFILLER_4_135 vgnd vpwr scs8hd_fill_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XANTENNA__171__B _169_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_9_249 vgnd vpwr scs8hd_decap_12
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XANTENNA__166__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_8_271 vgnd vpwr scs8hd_decap_4
XANTENNA__182__A _182_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_71 vpwr vgnd scs8hd_fill_2
Xmux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _202_/A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_24_25 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XFILLER_10_259 vgnd vpwr scs8hd_decap_12
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_252 vpwr vgnd scs8hd_fill_2
XFILLER_5_263 vpwr vgnd scs8hd_fill_2
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _183_/A mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_35_35 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vgnd vpwr scs8hd_decap_12
X_140_ _118_/A _143_/B _139_/X _103_/A _142_/B vgnd vpwr scs8hd_or4_4
XFILLER_18_134 vgnd vpwr scs8hd_decap_4
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XFILLER_25_90 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_178 vgnd vpwr scs8hd_decap_12
XANTENNA__163__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_72 vgnd vpwr scs8hd_fill_1
XFILLER_21_26 vpwr vgnd scs8hd_fill_2
XFILLER_30_129 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _221_/HI _206_/Y mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_123_ _130_/A _143_/B _100_/X _169_/A _124_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_7 vgnd vpwr scs8hd_fill_1
XFILLER_14_192 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _187_/Y mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
X_106_ address[0] _128_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_166 vgnd vpwr scs8hd_decap_4
XANTENNA__160__D _103_/A vgnd vpwr scs8hd_diode_2
XANTENNA__169__B _169_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_71 vpwr vgnd scs8hd_fill_2
XFILLER_27_36 vgnd vpwr scs8hd_decap_6
XFILLER_25_232 vgnd vpwr scs8hd_decap_12
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XANTENNA__095__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_4_169 vgnd vpwr scs8hd_decap_4
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XANTENNA__171__C _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_22_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_1_139 vpwr vgnd scs8hd_fill_2
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XFILLER_0_161 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _176_/A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__166__C address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_231 vgnd vpwr scs8hd_fill_1
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XFILLER_5_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_7.LATCH_1_.latch data_in _196_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_135 vgnd vpwr scs8hd_decap_12
XFILLER_19_26 vpwr vgnd scs8hd_fill_2
XFILLER_19_37 vgnd vpwr scs8hd_decap_4
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_35_47 vgnd vpwr scs8hd_decap_12
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_201 vpwr vgnd scs8hd_fill_2
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_26_190 vgnd vpwr scs8hd_decap_12
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__163__D _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_84 vgnd vpwr scs8hd_decap_3
XFILLER_24_105 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _216_/HI _180_/Y mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_21_49 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__098__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_105 vpwr vgnd scs8hd_fill_2
XFILLER_23_171 vgnd vpwr scs8hd_decap_12
XFILLER_7_18 vpwr vgnd scs8hd_fill_2
XFILLER_15_138 vgnd vpwr scs8hd_decap_4
XFILLER_15_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_122_ _163_/A _130_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _205_/A mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XFILLER_20_152 vgnd vpwr scs8hd_fill_1
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd
+ vpwr scs8hd_diode_2
X_105_ _127_/A _104_/X _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_112 vpwr vgnd scs8hd_fill_2
XFILLER_11_174 vgnd vpwr scs8hd_decap_8
XANTENNA__169__C _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_27_15 vpwr vgnd scs8hd_fill_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_107 vpwr vgnd scs8hd_fill_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_91 vgnd vpwr scs8hd_fill_1
XANTENNA__166__D _166_/D vgnd vpwr scs8hd_diode_2
XFILLER_24_49 vpwr vgnd scs8hd_fill_2
XFILLER_10_239 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_71 vpwr vgnd scs8hd_fill_2
XFILLER_5_210 vpwr vgnd scs8hd_fill_2
XFILLER_39_7 vpwr vgnd scs8hd_fill_2
XFILLER_27_147 vgnd vpwr scs8hd_decap_12
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_224 vgnd vpwr scs8hd_decap_8
XFILLER_18_125 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_41 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _209_/HI _182_/Y mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _179_/A mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_117 vgnd vpwr scs8hd_decap_3
X_121_ address[3] _163_/A vgnd vpwr scs8hd_inv_8
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
XFILLER_16_17 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_0_.latch data_in _207_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_104_ _118_/A _143_/B _100_/X _169_/A _104_/X vgnd vpwr scs8hd_or4_4
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_153 vpwr vgnd scs8hd_fill_2
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_21_7 vgnd vpwr scs8hd_decap_3
XFILLER_8_84 vpwr vgnd scs8hd_fill_2
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_138 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_171 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_3
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_1_119 vgnd vpwr scs8hd_decap_3
XFILLER_9_208 vgnd vpwr scs8hd_decap_4
XFILLER_9_219 vgnd vpwr scs8hd_decap_4
XFILLER_0_196 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_241 vgnd vpwr scs8hd_decap_12
XFILLER_5_96 vpwr vgnd scs8hd_fill_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_17 vpwr vgnd scs8hd_fill_2
XFILLER_30_93 vgnd vpwr scs8hd_decap_12
XFILLER_30_71 vgnd vpwr scs8hd_decap_12
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_27_159 vgnd vpwr scs8hd_decap_12
XFILLER_2_258 vgnd vpwr scs8hd_decap_12
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_25_71 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _200_/A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_64 vpwr vgnd scs8hd_fill_2
XFILLER_24_129 vgnd vpwr scs8hd_decap_12
Xmem_left_track_3.LATCH_1_.latch data_in _192_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
X_120_ _128_/A _118_/X _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_73 vpwr vgnd scs8hd_fill_2
XFILLER_11_95 vpwr vgnd scs8hd_fill_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_29 vpwr vgnd scs8hd_fill_2
XFILLER_20_154 vgnd vpwr scs8hd_decap_12
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_7_136 vpwr vgnd scs8hd_fill_2
XFILLER_11_187 vpwr vgnd scs8hd_fill_2
XFILLER_11_198 vpwr vgnd scs8hd_fill_2
X_103_ _103_/A _169_/A vgnd vpwr scs8hd_buf_1
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _220_/HI _204_/Y mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_63 vpwr vgnd scs8hd_fill_2
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_106 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _185_/Y mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_213 vgnd vpwr scs8hd_fill_1
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_60 vgnd vpwr scs8hd_fill_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_94 vpwr vgnd scs8hd_fill_2
XFILLER_22_227 vgnd vpwr scs8hd_decap_12
XFILLER_13_19 vpwr vgnd scs8hd_fill_2
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_0_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_253 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_75 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_15.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_15_ mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_135 vgnd vpwr scs8hd_decap_12
XFILLER_24_29 vpwr vgnd scs8hd_fill_2
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
XFILLER_14_40 vpwr vgnd scs8hd_fill_2
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
XFILLER_30_83 vgnd vpwr scs8hd_decap_8
XFILLER_5_234 vgnd vpwr scs8hd_decap_8
XFILLER_5_245 vgnd vpwr scs8hd_decap_3
XFILLER_5_256 vgnd vpwr scs8hd_decap_4
XFILLER_5_267 vgnd vpwr scs8hd_decap_8
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XFILLER_27_105 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _174_/A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_25_94 vgnd vpwr scs8hd_decap_12
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_10 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
XFILLER_17_182 vgnd vpwr scs8hd_fill_1
XFILLER_32_141 vgnd vpwr scs8hd_decap_12
XFILLER_21_19 vgnd vpwr scs8hd_decap_4
XFILLER_23_196 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_152 vgnd vpwr scs8hd_fill_1
X_179_ _179_/A _179_/Y vgnd vpwr scs8hd_inv_8
XFILLER_32_18 vgnd vpwr scs8hd_decap_12
XFILLER_20_166 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _215_/HI _178_/Y mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_104 vpwr vgnd scs8hd_fill_2
XFILLER_22_84 vpwr vgnd scs8hd_fill_2
XFILLER_22_62 vgnd vpwr scs8hd_decap_3
X_102_ address[1] _101_/Y _103_/A vgnd vpwr scs8hd_or2_4
Xmux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _203_/A mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_4_118 vpwr vgnd scs8hd_fill_2
XFILLER_17_73 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_195 vpwr vgnd scs8hd_fill_2
XANTENNA__104__A _118_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_239 vgnd vpwr scs8hd_decap_12
Xmem_left_track_13.LATCH_0_.latch data_in _203_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_165 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_0_.latch data_in _181_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _179_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_209 vgnd vpwr scs8hd_decap_4
Xmux_left_track_11.tap_buf4_0_.scs8hd_inv_1 mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _207_/Y mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _183_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_27_117 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_13.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_13_ mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_7 vpwr vgnd scs8hd_fill_2
XFILLER_2_205 vgnd vpwr scs8hd_decap_8
XFILLER_18_106 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_40 vpwr vgnd scs8hd_fill_2
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__112__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_260 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.tap_buf4_0_.scs8hd_inv_1 mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _233_/A vgnd vpwr scs8hd_inv_1
XFILLER_15_109 vpwr vgnd scs8hd_fill_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__107__A _128_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vgnd vpwr scs8hd_decap_3
XFILLER_20_178 vgnd vpwr scs8hd_decap_12
X_101_ enable _101_/Y vgnd vpwr scs8hd_inv_8
XFILLER_7_116 vgnd vpwr scs8hd_decap_4
XFILLER_11_134 vpwr vgnd scs8hd_fill_2
XFILLER_7_149 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _177_/A mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_43 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _181_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_19 vpwr vgnd scs8hd_fill_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _185_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_152 vpwr vgnd scs8hd_fill_2
XFILLER_3_141 vpwr vgnd scs8hd_fill_2
XANTENNA__104__B _143_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _128_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _198_/A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _236_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_251 vgnd vpwr scs8hd_decap_12
XFILLER_5_22 vgnd vpwr scs8hd_fill_1
XANTENNA__115__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_159 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _181_/Y mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_40_19 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_0_.latch data_in _189_/A _142_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_214 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_89 vgnd vpwr scs8hd_decap_3
XANTENNA__112__B _110_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
XFILLER_23_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_65 vpwr vgnd scs8hd_fill_2
XFILLER_11_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_11.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_177_ _177_/A _177_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__107__B _104_/X vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _130_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _222_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XFILLER_20_113 vgnd vpwr scs8hd_decap_8
XFILLER_20_124 vgnd vpwr scs8hd_decap_12
XFILLER_28_202 vgnd vpwr scs8hd_decap_12
X_100_ _130_/C _100_/X vgnd vpwr scs8hd_buf_1
XFILLER_11_157 vpwr vgnd scs8hd_fill_2
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XFILLER_8_22 vgnd vpwr scs8hd_decap_4
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
X_229_ _229_/A chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_6_161 vgnd vpwr scs8hd_decap_6
XFILLER_8_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_205 vgnd vpwr scs8hd_decap_8
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_30 vgnd vpwr scs8hd_decap_12
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XANTENNA__104__C _100_/X vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _118_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XFILLER_38_19 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _219_/HI _202_/Y mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_156 vgnd vpwr scs8hd_fill_1
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
XFILLER_28_63 vgnd vpwr scs8hd_decap_12
XFILLER_28_52 vgnd vpwr scs8hd_decap_8
XFILLER_28_41 vgnd vpwr scs8hd_decap_8
XFILLER_8_201 vgnd vpwr scs8hd_decap_12
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XANTENNA__115__B _130_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_34 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _183_/Y mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__131__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_54 vgnd vpwr scs8hd_decap_6
XFILLER_14_65 vgnd vpwr scs8hd_decap_4
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_171 vgnd vpwr scs8hd_decap_12
XANTENNA__126__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.LATCH_0_.latch data_in _177_/A _117_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_141 vgnd vpwr scs8hd_decap_12
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_18_119 vgnd vpwr scs8hd_decap_4
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XFILLER_25_75 vpwr vgnd scs8hd_fill_2
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_68 vpwr vgnd scs8hd_fill_2
XFILLER_2_46 vgnd vpwr scs8hd_decap_3
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XFILLER_2_6 vpwr vgnd scs8hd_fill_2
XFILLER_11_77 vgnd vpwr scs8hd_fill_1
XFILLER_11_99 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _172_/A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_176_ _176_/A _176_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__B _143_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_20_136 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_22_43 vpwr vgnd scs8hd_fill_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_269 vgnd vpwr scs8hd_decap_8
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_67 vpwr vgnd scs8hd_fill_2
XANTENNA__118__B _130_/B vgnd vpwr scs8hd_diode_2
X_228_ _228_/A chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_195 vgnd vpwr scs8hd_decap_6
XANTENNA__134__A _130_/A vgnd vpwr scs8hd_diode_2
X_159_ _169_/C _158_/B _159_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XFILLER_17_32 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_42 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_98 vpwr vgnd scs8hd_fill_2
XANTENNA__104__D _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_8 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _214_/HI _176_/Y mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__129__A _095_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _201_/A mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_28_75 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_5_79 vpwr vgnd scs8hd_fill_2
XANTENNA__115__C _100_/X vgnd vpwr scs8hd_diode_2
XANTENNA__131__B _130_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_22 vgnd vpwr scs8hd_decap_6
XFILLER_14_44 vgnd vpwr scs8hd_fill_1
XFILLER_14_88 vpwr vgnd scs8hd_fill_2
XANTENNA__232__A _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_227 vgnd vpwr scs8hd_decap_4
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XANTENNA__126__B _143_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_271 vgnd vpwr scs8hd_decap_4
XANTENNA__142__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XANTENNA__227__A _227_/A vgnd vpwr scs8hd_diode_2
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _205_/Y mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_13.LATCH_0_.latch data_in _185_/A _133_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA__137__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_23_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_34 vpwr vgnd scs8hd_fill_2
X_175_ _175_/A _175_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__C _100_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_7 vpwr vgnd scs8hd_fill_2
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_148 vgnd vpwr scs8hd_decap_4
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_88 vgnd vpwr scs8hd_decap_4
XFILLER_22_22 vgnd vpwr scs8hd_decap_4
XFILLER_7_108 vpwr vgnd scs8hd_fill_2
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
X_227_ _227_/A chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_8_35 vpwr vgnd scs8hd_fill_2
XANTENNA__118__C _100_/X vgnd vpwr scs8hd_diode_2
XANTENNA__134__B _130_/B vgnd vpwr scs8hd_diode_2
X_158_ _170_/C _158_/B _158_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__150__A _135_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_77 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XFILLER_33_54 vgnd vpwr scs8hd_decap_6
XFILLER_33_10 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_12
XANTENNA__235__A _235_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_199 vpwr vgnd scs8hd_fill_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _175_/A mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _205_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_0_114 vgnd vpwr scs8hd_decap_4
XFILLER_28_87 vgnd vpwr scs8hd_decap_4
XANTENNA__115__D _169_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_14 vpwr vgnd scs8hd_fill_2
XFILLER_10_6 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_1_.latch data_in _206_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _196_/A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_11 vgnd vpwr scs8hd_decap_4
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XANTENNA__142__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA__126__C _100_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _179_/Y mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_154 vgnd vpwr scs8hd_decap_12
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XANTENNA__243__A _243_/A vgnd vpwr scs8hd_diode_2
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_264 vgnd vpwr scs8hd_decap_12
XFILLER_1_253 vgnd vpwr scs8hd_decap_4
XFILLER_17_132 vpwr vgnd scs8hd_fill_2
XFILLER_17_143 vpwr vgnd scs8hd_fill_2
XFILLER_17_154 vgnd vpwr scs8hd_decap_12
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__153__A _130_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_135 vgnd vpwr scs8hd_decap_12
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _184_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XANTENNA__238__A _238_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_0_.latch data_in _173_/A _107_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_102 vpwr vgnd scs8hd_fill_2
XFILLER_22_190 vgnd vpwr scs8hd_decap_12
X_243_ _243_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_157 vgnd vpwr scs8hd_decap_8
XFILLER_14_168 vgnd vpwr scs8hd_decap_12
X_174_ _174_/A _174_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__D _169_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__148__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_11_138 vpwr vgnd scs8hd_fill_2
XFILLER_22_67 vgnd vpwr scs8hd_decap_4
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
X_226_ _226_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_6_131 vgnd vpwr scs8hd_decap_3
XFILLER_8_58 vgnd vpwr scs8hd_decap_3
XANTENNA__134__C _130_/C vgnd vpwr scs8hd_diode_2
XANTENNA__118__D _110_/D vgnd vpwr scs8hd_diode_2
X_157_ _130_/A address[2] _139_/X _109_/A _158_/B vgnd vpwr scs8hd_or4_4
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_9_ mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__150__B _149_/X vgnd vpwr scs8hd_diode_2
XFILLER_25_208 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_167 vpwr vgnd scs8hd_fill_2
XFILLER_3_134 vgnd vpwr scs8hd_decap_4
XANTENNA__145__B _143_/X vgnd vpwr scs8hd_diode_2
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__161__A _170_/C vgnd vpwr scs8hd_diode_2
XFILLER_12_200 vgnd vpwr scs8hd_decap_12
XFILLER_8_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__156__A _169_/C vgnd vpwr scs8hd_diode_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XFILLER_14_35 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
Xmux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _218_/HI _200_/Y mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__126__D _110_/D vgnd vpwr scs8hd_diode_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_23 vpwr vgnd scs8hd_fill_2
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_27 vpwr vgnd scs8hd_fill_2
XFILLER_1_276 vgnd vpwr scs8hd_fill_1
XFILLER_17_111 vgnd vpwr scs8hd_decap_4
XFILLER_17_166 vgnd vpwr scs8hd_decap_12
XANTENNA__153__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_147 vgnd vpwr scs8hd_decap_12
XFILLER_11_69 vpwr vgnd scs8hd_fill_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_125 vpwr vgnd scs8hd_fill_2
XFILLER_14_136 vgnd vpwr scs8hd_decap_12
X_242_ _242_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
X_173_ _173_/A _173_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _199_/A mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__148__B _148_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vgnd vpwr scs8hd_decap_4
XANTENNA__164__A _170_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _223_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_8_26 vgnd vpwr scs8hd_fill_1
XANTENNA__134__D _110_/D vgnd vpwr scs8hd_diode_2
X_156_ _169_/C _156_/B _156_/Y vgnd vpwr scs8hd_nor2_4
X_225_ _225_/HI _225_/LO vgnd vpwr scs8hd_conb_1
XFILLER_40_7 vgnd vpwr scs8hd_decap_12
XFILLER_33_6 vpwr vgnd scs8hd_fill_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _169_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_3_102 vgnd vpwr scs8hd_decap_3
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__161__B _161_/B vgnd vpwr scs8hd_diode_2
X_139_ _163_/C _139_/X vgnd vpwr scs8hd_buf_1
Xmux_left_track_7.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_7_ mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_138 vpwr vgnd scs8hd_fill_2
XFILLER_12_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_38 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _156_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _174_/Y mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _242_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_14 vpwr vgnd scs8hd_fill_2
XFILLER_30_35 vgnd vpwr scs8hd_decap_12
XFILLER_39_11 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A _166_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_178 vgnd vpwr scs8hd_decap_12
XPHY_46 vgnd vpwr scs8hd_decap_3
Xmem_left_track_13.LATCH_1_.latch data_in _202_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_9_3 vpwr vgnd scs8hd_fill_2
XFILLER_17_178 vgnd vpwr scs8hd_decap_4
XANTENNA__153__C _139_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_159 vgnd vpwr scs8hd_decap_12
XFILLER_11_15 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_1_.latch data_in _180_/A _124_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_148 vgnd vpwr scs8hd_decap_4
X_172_ _172_/A _172_/Y vgnd vpwr scs8hd_inv_8
X_241_ _241_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__164__B _165_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_130 vpwr vgnd scs8hd_fill_2
XFILLER_13_170 vgnd vpwr scs8hd_decap_12
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _203_/Y mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XFILLER_22_47 vpwr vgnd scs8hd_fill_2
XFILLER_22_14 vpwr vgnd scs8hd_fill_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_0_.latch data_in _199_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_224_ _224_/HI _224_/LO vgnd vpwr scs8hd_conb_1
X_155_ address[0] _169_/C vgnd vpwr scs8hd_buf_1
XFILLER_26_6 vpwr vgnd scs8hd_fill_2
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _158_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_36 vpwr vgnd scs8hd_fill_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
XFILLER_30_202 vgnd vpwr scs8hd_decap_12
X_207_ _207_/A _207_/Y vgnd vpwr scs8hd_inv_8
X_138_ address[4] _166_/D _163_/C vgnd vpwr scs8hd_nand2_4
XFILLER_24_3 vgnd vpwr scs8hd_fill_1
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
XFILLER_0_83 vpwr vgnd scs8hd_fill_2
XFILLER_21_257 vgnd vpwr scs8hd_decap_12
XFILLER_9_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XFILLER_30_47 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _173_/A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_23 vgnd vpwr scs8hd_decap_12
XFILLER_29_110 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_5_ mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _181_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _185_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_25_36 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XFILLER_1_234 vgnd vpwr scs8hd_decap_8
XFILLER_1_212 vpwr vgnd scs8hd_fill_2
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _194_/A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__153__D _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_105 vgnd vpwr scs8hd_decap_12
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_171 vgnd vpwr scs8hd_decap_12
XFILLER_11_38 vgnd vpwr scs8hd_decap_4
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
X_240_ _240_/A chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
X_171_ _110_/D _169_/B _169_/C _171_/Y vgnd vpwr scs8hd_nor3_4
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _177_/Y mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_1_.latch data_in _188_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_164 vpwr vgnd scs8hd_fill_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_13_182 vgnd vpwr scs8hd_fill_1
XFILLER_9_197 vgnd vpwr scs8hd_decap_4
XFILLER_3_83 vpwr vgnd scs8hd_fill_2
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_26 vgnd vpwr scs8hd_fill_1
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
XFILLER_8_39 vpwr vgnd scs8hd_fill_2
XFILLER_10_141 vpwr vgnd scs8hd_fill_2
X_223_ _223_/HI _223_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_112 vpwr vgnd scs8hd_fill_2
XFILLER_6_145 vgnd vpwr scs8hd_decap_6
XFILLER_6_178 vgnd vpwr scs8hd_decap_6
XFILLER_10_163 vgnd vpwr scs8hd_decap_12
X_154_ _170_/C _156_/B _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _225_/HI _198_/Y mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _238_/A vgnd vpwr scs8hd_inv_1
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_15 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_14 vpwr vgnd scs8hd_fill_2
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_148 vpwr vgnd scs8hd_fill_2
X_206_ _206_/A _206_/Y vgnd vpwr scs8hd_inv_8
X_137_ address[5] _166_/D vgnd vpwr scs8hd_inv_8
XFILLER_17_3 vgnd vpwr scs8hd_decap_3
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XFILLER_9_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _187_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_25 vgnd vpwr scs8hd_decap_6
XFILLER_0_107 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _095_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_218 vgnd vpwr scs8hd_decap_8
XFILLER_8_229 vgnd vpwr scs8hd_decap_12
XFILLER_5_18 vgnd vpwr scs8hd_decap_4
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_59 vgnd vpwr scs8hd_decap_12
XFILLER_39_35 vgnd vpwr scs8hd_decap_12
XFILLER_4_232 vgnd vpwr scs8hd_fill_1
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _230_/A vgnd vpwr scs8hd_inv_1
XFILLER_6_72 vpwr vgnd scs8hd_fill_2
XFILLER_6_83 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _173_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_136 vpwr vgnd scs8hd_fill_2
XFILLER_17_147 vgnd vpwr scs8hd_decap_4
XFILLER_32_117 vgnd vpwr scs8hd_decap_12
XFILLER_15_92 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_3_ mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_117 vgnd vpwr scs8hd_decap_4
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
X_170_ _110_/D _169_/B _170_/C _170_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_14_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_62 vpwr vgnd scs8hd_fill_2
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.LATCH_1_.latch data_in _176_/A _116_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_222_ _222_/HI _222_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_102 vpwr vgnd scs8hd_fill_2
XFILLER_8_18 vpwr vgnd scs8hd_fill_2
XFILLER_8_29 vpwr vgnd scs8hd_fill_2
XFILLER_10_175 vpwr vgnd scs8hd_fill_2
XFILLER_10_186 vgnd vpwr scs8hd_decap_8
X_153_ _130_/A address[2] _139_/X _103_/A _156_/B vgnd vpwr scs8hd_or4_4
XFILLER_6_157 vpwr vgnd scs8hd_fill_2
XFILLER_10_197 vgnd vpwr scs8hd_decap_12
XFILLER_12_60 vgnd vpwr scs8hd_decap_8
XFILLER_12_71 vpwr vgnd scs8hd_fill_2
XFILLER_19_7 vgnd vpwr scs8hd_decap_4
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _197_/A mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_49 vpwr vgnd scs8hd_fill_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_138 vgnd vpwr scs8hd_fill_1
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
X_205_ _205_/A _205_/Y vgnd vpwr scs8hd_inv_8
Xmem_left_track_5.LATCH_0_.latch data_in _195_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_136_ _133_/A _135_/B _136_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_182 vpwr vgnd scs8hd_fill_2
XFILLER_0_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_15 vpwr vgnd scs8hd_fill_2
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
X_119_ _127_/A _118_/X _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_252 vgnd vpwr scs8hd_decap_3
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_28 vgnd vpwr scs8hd_fill_1
XFILLER_39_47 vgnd vpwr scs8hd_decap_12
XFILLER_29_123 vgnd vpwr scs8hd_decap_12
XFILLER_4_211 vgnd vpwr scs8hd_decap_3
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _208_/HI _172_/Y mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_32_129 vgnd vpwr scs8hd_decap_12
XFILLER_17_115 vgnd vpwr scs8hd_fill_1
XFILLER_15_71 vgnd vpwr scs8hd_decap_4
XFILLER_16_181 vgnd vpwr scs8hd_decap_12
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
XFILLER_26_70 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_1_ mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _224_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_232 vgnd vpwr scs8hd_decap_12
X_221_ _221_/HI _221_/LO vgnd vpwr scs8hd_conb_1
X_152_ _095_/Y _170_/C vgnd vpwr scs8hd_buf_1
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_13.LATCH_1_.latch data_in _184_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_202 vgnd vpwr scs8hd_decap_12
Xmux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _201_/Y mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_7.INVTX1_1_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
XFILLER_23_93 vgnd vpwr scs8hd_decap_12
XFILLER_23_60 vgnd vpwr scs8hd_fill_1
X_135_ _135_/A _135_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_31_7 vpwr vgnd scs8hd_fill_2
XFILLER_9_40 vpwr vgnd scs8hd_fill_2
XFILLER_12_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
X_118_ _118_/A _130_/B _100_/X _110_/D _118_/X vgnd vpwr scs8hd_or4_4
XFILLER_22_3 vpwr vgnd scs8hd_fill_2
XFILLER_14_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XFILLER_29_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_83 vpwr vgnd scs8hd_fill_2
XFILLER_28_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_105 vgnd vpwr scs8hd_decap_12
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_25_171 vgnd vpwr scs8hd_decap_12
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _205_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_193 vgnd vpwr scs8hd_decap_12
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_11_19 vpwr vgnd scs8hd_fill_2
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_14_119 vgnd vpwr scs8hd_decap_4
XFILLER_22_152 vgnd vpwr scs8hd_fill_1
XFILLER_26_93 vgnd vpwr scs8hd_decap_12
XFILLER_9_123 vpwr vgnd scs8hd_fill_2
XFILLER_9_134 vpwr vgnd scs8hd_fill_2
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _192_/A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_22_29 vpwr vgnd scs8hd_fill_2
XFILLER_22_18 vpwr vgnd scs8hd_fill_2
X_220_ _220_/HI _220_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
X_151_ _133_/A _149_/X _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _175_/Y mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
X_134_ _130_/A _130_/B _130_/C _110_/D _135_/B vgnd vpwr scs8hd_or4_4
Xmem_bottom_track_1.LATCH_1_.latch data_in _172_/A _105_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_10 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_0_76 vpwr vgnd scs8hd_fill_2
XFILLER_0_87 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _184_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _224_/HI _196_/Y mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_239 vgnd vpwr scs8hd_decap_12
XFILLER_18_50 vgnd vpwr scs8hd_decap_6
XFILLER_18_72 vpwr vgnd scs8hd_fill_2
XFILLER_18_83 vgnd vpwr scs8hd_decap_3
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _207_/A vgnd vpwr
+ scs8hd_diode_2
X_117_ _128_/A _115_/X _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_210 vgnd vpwr scs8hd_decap_4
XFILLER_7_221 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.INVTX1_1_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_232 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.LATCH_0_.latch data_in _191_/A _145_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_3 vgnd vpwr scs8hd_decap_4
XFILLER_29_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_224 vgnd vpwr scs8hd_decap_8
XFILLER_20_62 vpwr vgnd scs8hd_fill_2
XFILLER_26_117 vgnd vpwr scs8hd_decap_12
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_1_249 vpwr vgnd scs8hd_fill_2
XFILLER_1_216 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_39_220 vgnd vpwr scs8hd_decap_12
XFILLER_22_120 vgnd vpwr scs8hd_decap_12
XFILLER_26_83 vpwr vgnd scs8hd_fill_2
XFILLER_9_168 vpwr vgnd scs8hd_fill_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _186_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_12
X_150_ _135_/A _149_/X _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_127 vpwr vgnd scs8hd_fill_2
XFILLER_10_145 vgnd vpwr scs8hd_decap_6
XFILLER_12_96 vgnd vpwr scs8hd_decap_8
XFILLER_5_193 vpwr vgnd scs8hd_fill_2
XFILLER_17_19 vpwr vgnd scs8hd_fill_2
XFILLER_33_18 vgnd vpwr scs8hd_decap_12
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_62 vgnd vpwr scs8hd_decap_3
X_133_ _133_/A _130_/X _133_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__110__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_9_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _172_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _195_/A mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__105__A _127_/A vgnd vpwr scs8hd_diode_2
X_116_ _127_/A _115_/X _116_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_19 vgnd vpwr scs8hd_decap_12
XFILLER_29_159 vgnd vpwr scs8hd_decap_12
XFILLER_20_41 vgnd vpwr scs8hd_decap_8
XFILLER_6_21 vgnd vpwr scs8hd_fill_1
XFILLER_6_43 vgnd vpwr scs8hd_fill_1
XFILLER_6_76 vpwr vgnd scs8hd_fill_2
XFILLER_6_87 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_19 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.INVTX1_1_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_184 vgnd vpwr scs8hd_decap_12
XFILLER_15_30 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XANTENNA__102__B _101_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _199_/Y mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_110 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_232 vgnd vpwr scs8hd_decap_12
XFILLER_22_154 vgnd vpwr scs8hd_decap_12
XFILLER_22_132 vgnd vpwr scs8hd_decap_12
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_147 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_6_106 vgnd vpwr scs8hd_decap_4
XFILLER_10_124 vpwr vgnd scs8hd_fill_2
XFILLER_5_3 vpwr vgnd scs8hd_fill_2
XFILLER_18_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__108__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vpwr vgnd scs8hd_fill_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_74 vpwr vgnd scs8hd_fill_2
X_132_ address[0] _133_/A vgnd vpwr scs8hd_buf_1
XFILLER_2_186 vgnd vpwr scs8hd_decap_4
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B _143_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
XFILLER_28_19 vgnd vpwr scs8hd_decap_4
XFILLER_20_263 vgnd vpwr scs8hd_decap_12
XFILLER_18_41 vgnd vpwr scs8hd_decap_3
XANTENNA__105__B _104_/X vgnd vpwr scs8hd_diode_2
X_115_ _118_/A _130_/B _100_/X _169_/A _115_/X vgnd vpwr scs8hd_or4_4
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XANTENNA__121__A address[3] vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in _198_/A _158_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_237 vgnd vpwr scs8hd_decap_8
XFILLER_4_248 vgnd vpwr scs8hd_decap_8
XFILLER_29_62 vgnd vpwr scs8hd_decap_12
XFILLER_4_259 vgnd vpwr scs8hd_decap_12
XANTENNA__116__A _127_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_55 vgnd vpwr scs8hd_decap_8
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
XFILLER_19_182 vgnd vpwr scs8hd_fill_1
XFILLER_1_229 vgnd vpwr scs8hd_decap_3
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_196 vgnd vpwr scs8hd_decap_12
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XFILLER_31_41 vgnd vpwr scs8hd_decap_12
XFILLER_16_152 vgnd vpwr scs8hd_fill_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

