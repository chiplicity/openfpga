VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_top
  CLASS BLOCK ;
  FOREIGN grid_io_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 144.670 BY 120.000 ;
  PIN bottom_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.280 0.000 69.560 2.400 ;
    END
  END bottom_width_0_height_0__pin_0_
  PIN bottom_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.420 0.000 119.700 2.400 ;
    END
  END bottom_width_0_height_0__pin_1_lower
  PIN bottom_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.600 0.000 19.880 2.400 ;
    END
  END bottom_width_0_height_0__pin_1_upper
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 142.270 59.200 144.670 59.800 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 142.270 99.320 144.670 99.920 ;
    END
  END ccff_tail
  PIN gfpga_pad_GPIO_A
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.160 117.600 13.440 120.000 ;
    END
  END gfpga_pad_GPIO_A
  PIN gfpga_pad_GPIO_IE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.420 117.600 50.700 120.000 ;
    END
  END gfpga_pad_GPIO_IE
  PIN gfpga_pad_GPIO_OE
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.140 117.600 88.420 120.000 ;
    END
  END gfpga_pad_GPIO_OE
  PIN gfpga_pad_GPIO_Y
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 125.400 117.600 125.680 120.000 ;
    END
  END gfpga_pad_GPIO_Y
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 142.270 19.760 144.670 20.360 ;
    END
  END prog_clk
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.390 10.640 25.990 109.040 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.390 10.640 50.990 109.040 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.190 10.795 139.110 108.885 ;
      LAYER met1 ;
        RECT 0.190 10.640 139.110 109.780 ;
      LAYER met2 ;
        RECT 13.720 117.320 50.140 117.600 ;
        RECT 50.980 117.320 87.860 117.600 ;
        RECT 88.700 117.320 125.120 117.600 ;
        RECT 13.230 2.680 125.930 117.320 ;
        RECT 13.230 2.400 19.320 2.680 ;
        RECT 20.160 2.400 69.000 2.680 ;
        RECT 69.840 2.400 119.140 2.680 ;
        RECT 119.980 2.400 125.930 2.680 ;
      LAYER met3 ;
        RECT 14.975 100.320 142.270 108.965 ;
        RECT 14.975 98.920 141.870 100.320 ;
        RECT 14.975 60.200 142.270 98.920 ;
        RECT 14.975 58.800 141.870 60.200 ;
        RECT 14.975 20.760 142.270 58.800 ;
        RECT 14.975 19.360 141.870 20.760 ;
        RECT 14.975 10.715 142.270 19.360 ;
      LAYER met4 ;
        RECT 74.390 10.640 125.990 109.040 ;
  END
END grid_io_top
END LIBRARY

