VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 2.400 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.450 197.600 191.730 200.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 2.400 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.970 197.600 197.250 200.000 ;
    END
  END SC_OUT_TOP
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 2.400 ;
    END
  END Test_en
  PIN bottom_width_0_height_0__pin_50_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.400 ;
    END
  END bottom_width_0_height_0__pin_50_
  PIN bottom_width_0_height_0__pin_51_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.400 ;
    END
  END bottom_width_0_height_0__pin_51_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 51.040 200.000 51.640 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 2.400 ;
    END
  END clk
  PIN left_width_0_height_0__pin_52_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 2.400 167.240 ;
    END
  END left_width_0_height_0__pin_52_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END prog_clk
  PIN right_width_0_height_0__pin_16_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 57.160 200.000 57.760 ;
    END
  END right_width_0_height_0__pin_16_
  PIN right_width_0_height_0__pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 63.280 200.000 63.880 ;
    END
  END right_width_0_height_0__pin_17_
  PIN right_width_0_height_0__pin_18_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 69.400 200.000 70.000 ;
    END
  END right_width_0_height_0__pin_18_
  PIN right_width_0_height_0__pin_19_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 74.840 200.000 75.440 ;
    END
  END right_width_0_height_0__pin_19_
  PIN right_width_0_height_0__pin_20_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 80.960 200.000 81.560 ;
    END
  END right_width_0_height_0__pin_20_
  PIN right_width_0_height_0__pin_21_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 87.080 200.000 87.680 ;
    END
  END right_width_0_height_0__pin_21_
  PIN right_width_0_height_0__pin_22_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 93.200 200.000 93.800 ;
    END
  END right_width_0_height_0__pin_22_
  PIN right_width_0_height_0__pin_23_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 99.320 200.000 99.920 ;
    END
  END right_width_0_height_0__pin_23_
  PIN right_width_0_height_0__pin_24_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 105.440 200.000 106.040 ;
    END
  END right_width_0_height_0__pin_24_
  PIN right_width_0_height_0__pin_25_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 111.560 200.000 112.160 ;
    END
  END right_width_0_height_0__pin_25_
  PIN right_width_0_height_0__pin_26_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 117.680 200.000 118.280 ;
    END
  END right_width_0_height_0__pin_26_
  PIN right_width_0_height_0__pin_27_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 123.800 200.000 124.400 ;
    END
  END right_width_0_height_0__pin_27_
  PIN right_width_0_height_0__pin_28_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 129.920 200.000 130.520 ;
    END
  END right_width_0_height_0__pin_28_
  PIN right_width_0_height_0__pin_29_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 136.040 200.000 136.640 ;
    END
  END right_width_0_height_0__pin_29_
  PIN right_width_0_height_0__pin_30_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 141.480 200.000 142.080 ;
    END
  END right_width_0_height_0__pin_30_
  PIN right_width_0_height_0__pin_31_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 147.600 200.000 148.200 ;
    END
  END right_width_0_height_0__pin_31_
  PIN right_width_0_height_0__pin_42_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 2.760 200.000 3.360 ;
    END
  END right_width_0_height_0__pin_42_lower
  PIN right_width_0_height_0__pin_42_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 153.720 200.000 154.320 ;
    END
  END right_width_0_height_0__pin_42_upper
  PIN right_width_0_height_0__pin_43_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 8.200 200.000 8.800 ;
    END
  END right_width_0_height_0__pin_43_lower
  PIN right_width_0_height_0__pin_43_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 159.840 200.000 160.440 ;
    END
  END right_width_0_height_0__pin_43_upper
  PIN right_width_0_height_0__pin_44_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 14.320 200.000 14.920 ;
    END
  END right_width_0_height_0__pin_44_lower
  PIN right_width_0_height_0__pin_44_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 165.960 200.000 166.560 ;
    END
  END right_width_0_height_0__pin_44_upper
  PIN right_width_0_height_0__pin_45_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 20.440 200.000 21.040 ;
    END
  END right_width_0_height_0__pin_45_lower
  PIN right_width_0_height_0__pin_45_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 172.080 200.000 172.680 ;
    END
  END right_width_0_height_0__pin_45_upper
  PIN right_width_0_height_0__pin_46_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 26.560 200.000 27.160 ;
    END
  END right_width_0_height_0__pin_46_lower
  PIN right_width_0_height_0__pin_46_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 178.200 200.000 178.800 ;
    END
  END right_width_0_height_0__pin_46_upper
  PIN right_width_0_height_0__pin_47_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 32.680 200.000 33.280 ;
    END
  END right_width_0_height_0__pin_47_lower
  PIN right_width_0_height_0__pin_47_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 184.320 200.000 184.920 ;
    END
  END right_width_0_height_0__pin_47_upper
  PIN right_width_0_height_0__pin_48_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 38.800 200.000 39.400 ;
    END
  END right_width_0_height_0__pin_48_lower
  PIN right_width_0_height_0__pin_48_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 190.440 200.000 191.040 ;
    END
  END right_width_0_height_0__pin_48_upper
  PIN right_width_0_height_0__pin_49_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 44.920 200.000 45.520 ;
    END
  END right_width_0_height_0__pin_49_lower
  PIN right_width_0_height_0__pin_49_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 196.560 200.000 197.160 ;
    END
  END right_width_0_height_0__pin_49_upper
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 197.600 47.290 200.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.670 197.600 102.950 200.000 ;
    END
  END top_width_0_height_0__pin_10_
  PIN top_width_0_height_0__pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.190 197.600 108.470 200.000 ;
    END
  END top_width_0_height_0__pin_11_
  PIN top_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.710 197.600 113.990 200.000 ;
    END
  END top_width_0_height_0__pin_12_
  PIN top_width_0_height_0__pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.230 197.600 119.510 200.000 ;
    END
  END top_width_0_height_0__pin_13_
  PIN top_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.750 197.600 125.030 200.000 ;
    END
  END top_width_0_height_0__pin_14_
  PIN top_width_0_height_0__pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.270 197.600 130.550 200.000 ;
    END
  END top_width_0_height_0__pin_15_
  PIN top_width_0_height_0__pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 197.600 52.810 200.000 ;
    END
  END top_width_0_height_0__pin_1_
  PIN top_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 197.600 58.330 200.000 ;
    END
  END top_width_0_height_0__pin_2_
  PIN top_width_0_height_0__pin_32_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.250 197.600 136.530 200.000 ;
    END
  END top_width_0_height_0__pin_32_
  PIN top_width_0_height_0__pin_33_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.770 197.600 142.050 200.000 ;
    END
  END top_width_0_height_0__pin_33_
  PIN top_width_0_height_0__pin_34_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 147.290 197.600 147.570 200.000 ;
    END
  END top_width_0_height_0__pin_34_lower
  PIN top_width_0_height_0__pin_34_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 197.600 3.130 200.000 ;
    END
  END top_width_0_height_0__pin_34_upper
  PIN top_width_0_height_0__pin_35_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 152.810 197.600 153.090 200.000 ;
    END
  END top_width_0_height_0__pin_35_lower
  PIN top_width_0_height_0__pin_35_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 8.370 197.600 8.650 200.000 ;
    END
  END top_width_0_height_0__pin_35_upper
  PIN top_width_0_height_0__pin_36_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 158.330 197.600 158.610 200.000 ;
    END
  END top_width_0_height_0__pin_36_lower
  PIN top_width_0_height_0__pin_36_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 13.890 197.600 14.170 200.000 ;
    END
  END top_width_0_height_0__pin_36_upper
  PIN top_width_0_height_0__pin_37_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.850 197.600 164.130 200.000 ;
    END
  END top_width_0_height_0__pin_37_lower
  PIN top_width_0_height_0__pin_37_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.410 197.600 19.690 200.000 ;
    END
  END top_width_0_height_0__pin_37_upper
  PIN top_width_0_height_0__pin_38_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 169.370 197.600 169.650 200.000 ;
    END
  END top_width_0_height_0__pin_38_lower
  PIN top_width_0_height_0__pin_38_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 197.600 25.210 200.000 ;
    END
  END top_width_0_height_0__pin_38_upper
  PIN top_width_0_height_0__pin_39_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.890 197.600 175.170 200.000 ;
    END
  END top_width_0_height_0__pin_39_lower
  PIN top_width_0_height_0__pin_39_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.450 197.600 30.730 200.000 ;
    END
  END top_width_0_height_0__pin_39_upper
  PIN top_width_0_height_0__pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 197.600 63.850 200.000 ;
    END
  END top_width_0_height_0__pin_3_
  PIN top_width_0_height_0__pin_40_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.410 197.600 180.690 200.000 ;
    END
  END top_width_0_height_0__pin_40_lower
  PIN top_width_0_height_0__pin_40_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.970 197.600 36.250 200.000 ;
    END
  END top_width_0_height_0__pin_40_upper
  PIN top_width_0_height_0__pin_41_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.930 197.600 186.210 200.000 ;
    END
  END top_width_0_height_0__pin_41_lower
  PIN top_width_0_height_0__pin_41_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.490 197.600 41.770 200.000 ;
    END
  END top_width_0_height_0__pin_41_upper
  PIN top_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 197.600 69.830 200.000 ;
    END
  END top_width_0_height_0__pin_4_
  PIN top_width_0_height_0__pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.070 197.600 75.350 200.000 ;
    END
  END top_width_0_height_0__pin_5_
  PIN top_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.590 197.600 80.870 200.000 ;
    END
  END top_width_0_height_0__pin_6_
  PIN top_width_0_height_0__pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.110 197.600 86.390 200.000 ;
    END
  END top_width_0_height_0__pin_7_
  PIN top_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.630 197.600 91.910 200.000 ;
    END
  END top_width_0_height_0__pin_8_
  PIN top_width_0_height_0__pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.150 197.600 97.430 200.000 ;
    END
  END top_width_0_height_0__pin_9_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 2.830 10.640 194.120 187.920 ;
      LAYER met2 ;
        RECT 3.410 197.320 8.090 197.610 ;
        RECT 8.930 197.320 13.610 197.610 ;
        RECT 14.450 197.320 19.130 197.610 ;
        RECT 19.970 197.320 24.650 197.610 ;
        RECT 25.490 197.320 30.170 197.610 ;
        RECT 31.010 197.320 35.690 197.610 ;
        RECT 36.530 197.320 41.210 197.610 ;
        RECT 42.050 197.320 46.730 197.610 ;
        RECT 47.570 197.320 52.250 197.610 ;
        RECT 53.090 197.320 57.770 197.610 ;
        RECT 58.610 197.320 63.290 197.610 ;
        RECT 64.130 197.320 69.270 197.610 ;
        RECT 70.110 197.320 74.790 197.610 ;
        RECT 75.630 197.320 80.310 197.610 ;
        RECT 81.150 197.320 85.830 197.610 ;
        RECT 86.670 197.320 91.350 197.610 ;
        RECT 92.190 197.320 96.870 197.610 ;
        RECT 97.710 197.320 102.390 197.610 ;
        RECT 103.230 197.320 107.910 197.610 ;
        RECT 108.750 197.320 113.430 197.610 ;
        RECT 114.270 197.320 118.950 197.610 ;
        RECT 119.790 197.320 124.470 197.610 ;
        RECT 125.310 197.320 129.990 197.610 ;
        RECT 130.830 197.320 135.970 197.610 ;
        RECT 136.810 197.320 141.490 197.610 ;
        RECT 142.330 197.320 147.010 197.610 ;
        RECT 147.850 197.320 152.530 197.610 ;
        RECT 153.370 197.320 158.050 197.610 ;
        RECT 158.890 197.320 163.570 197.610 ;
        RECT 164.410 197.320 169.090 197.610 ;
        RECT 169.930 197.320 174.610 197.610 ;
        RECT 175.450 197.320 180.130 197.610 ;
        RECT 180.970 197.320 185.650 197.610 ;
        RECT 186.490 197.320 191.170 197.610 ;
        RECT 192.010 197.320 196.690 197.610 ;
        RECT 2.850 2.680 197.250 197.320 ;
        RECT 2.850 2.400 16.370 2.680 ;
        RECT 17.210 2.400 49.490 2.680 ;
        RECT 50.330 2.400 83.070 2.680 ;
        RECT 83.910 2.400 116.190 2.680 ;
        RECT 117.030 2.400 149.770 2.680 ;
        RECT 150.610 2.400 182.890 2.680 ;
        RECT 183.730 2.400 197.250 2.680 ;
      LAYER met3 ;
        RECT 2.400 196.160 197.200 197.025 ;
        RECT 2.400 191.440 197.600 196.160 ;
        RECT 2.400 190.040 197.200 191.440 ;
        RECT 2.400 185.320 197.600 190.040 ;
        RECT 2.400 183.920 197.200 185.320 ;
        RECT 2.400 179.200 197.600 183.920 ;
        RECT 2.400 177.800 197.200 179.200 ;
        RECT 2.400 173.080 197.600 177.800 ;
        RECT 2.400 171.680 197.200 173.080 ;
        RECT 2.400 167.640 197.600 171.680 ;
        RECT 2.800 166.960 197.600 167.640 ;
        RECT 2.800 166.240 197.200 166.960 ;
        RECT 2.400 165.560 197.200 166.240 ;
        RECT 2.400 160.840 197.600 165.560 ;
        RECT 2.400 159.440 197.200 160.840 ;
        RECT 2.400 154.720 197.600 159.440 ;
        RECT 2.400 153.320 197.200 154.720 ;
        RECT 2.400 148.600 197.600 153.320 ;
        RECT 2.400 147.200 197.200 148.600 ;
        RECT 2.400 142.480 197.600 147.200 ;
        RECT 2.400 141.080 197.200 142.480 ;
        RECT 2.400 137.040 197.600 141.080 ;
        RECT 2.400 135.640 197.200 137.040 ;
        RECT 2.400 130.920 197.600 135.640 ;
        RECT 2.400 129.520 197.200 130.920 ;
        RECT 2.400 124.800 197.600 129.520 ;
        RECT 2.400 123.400 197.200 124.800 ;
        RECT 2.400 118.680 197.600 123.400 ;
        RECT 2.400 117.280 197.200 118.680 ;
        RECT 2.400 112.560 197.600 117.280 ;
        RECT 2.400 111.160 197.200 112.560 ;
        RECT 2.400 106.440 197.600 111.160 ;
        RECT 2.400 105.040 197.200 106.440 ;
        RECT 2.400 101.000 197.600 105.040 ;
        RECT 2.800 100.320 197.600 101.000 ;
        RECT 2.800 99.600 197.200 100.320 ;
        RECT 2.400 98.920 197.200 99.600 ;
        RECT 2.400 94.200 197.600 98.920 ;
        RECT 2.400 92.800 197.200 94.200 ;
        RECT 2.400 88.080 197.600 92.800 ;
        RECT 2.400 86.680 197.200 88.080 ;
        RECT 2.400 81.960 197.600 86.680 ;
        RECT 2.400 80.560 197.200 81.960 ;
        RECT 2.400 75.840 197.600 80.560 ;
        RECT 2.400 74.440 197.200 75.840 ;
        RECT 2.400 70.400 197.600 74.440 ;
        RECT 2.400 69.000 197.200 70.400 ;
        RECT 2.400 64.280 197.600 69.000 ;
        RECT 2.400 62.880 197.200 64.280 ;
        RECT 2.400 58.160 197.600 62.880 ;
        RECT 2.400 56.760 197.200 58.160 ;
        RECT 2.400 52.040 197.600 56.760 ;
        RECT 2.400 50.640 197.200 52.040 ;
        RECT 2.400 45.920 197.600 50.640 ;
        RECT 2.400 44.520 197.200 45.920 ;
        RECT 2.400 39.800 197.600 44.520 ;
        RECT 2.400 38.400 197.200 39.800 ;
        RECT 2.400 34.360 197.600 38.400 ;
        RECT 2.800 33.680 197.600 34.360 ;
        RECT 2.800 32.960 197.200 33.680 ;
        RECT 2.400 32.280 197.200 32.960 ;
        RECT 2.400 27.560 197.600 32.280 ;
        RECT 2.400 26.160 197.200 27.560 ;
        RECT 2.400 21.440 197.600 26.160 ;
        RECT 2.400 20.040 197.200 21.440 ;
        RECT 2.400 15.320 197.600 20.040 ;
        RECT 2.400 13.920 197.200 15.320 ;
        RECT 2.400 9.200 197.600 13.920 ;
        RECT 2.400 7.800 197.200 9.200 ;
        RECT 2.400 3.760 197.600 7.800 ;
        RECT 2.400 2.895 197.200 3.760 ;
      LAYER met4 ;
        RECT 24.710 10.640 97.440 187.920 ;
        RECT 99.840 10.640 177.265 187.920 ;
      LAYER met5 ;
        RECT 24.500 174.300 125.460 179.300 ;
  END
END grid_clb
END LIBRARY

