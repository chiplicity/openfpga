VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 138.600 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.320 2.400 33.920 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.360 2.400 103.960 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 17.680 140.000 18.280 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 47.600 140.000 48.200 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 50.320 140.000 50.920 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 53.040 140.000 53.640 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 56.440 140.000 57.040 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 59.160 140.000 59.760 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 62.560 140.000 63.160 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 65.280 140.000 65.880 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 68.000 140.000 68.600 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 71.400 140.000 72.000 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 74.120 140.000 74.720 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 20.400 140.000 21.000 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 23.800 140.000 24.400 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 26.520 140.000 27.120 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 29.240 140.000 29.840 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 32.640 140.000 33.240 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 35.360 140.000 35.960 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 38.080 140.000 38.680 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 41.480 140.000 42.080 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.200 140.000 44.800 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 76.840 140.000 77.440 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 106.760 140.000 107.360 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 110.160 140.000 110.760 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 112.880 140.000 113.480 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 115.600 140.000 116.200 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 119.000 140.000 119.600 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 121.720 140.000 122.320 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 125.120 140.000 125.720 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 127.840 140.000 128.440 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 130.560 140.000 131.160 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 133.960 140.000 134.560 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 80.240 140.000 80.840 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 82.960 140.000 83.560 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 86.360 140.000 86.960 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 89.080 140.000 89.680 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 91.800 140.000 92.400 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 95.200 140.000 95.800 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 97.920 140.000 98.520 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 101.320 140.000 101.920 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 104.040 140.000 104.640 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 136.200 4.970 138.600 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 136.200 39.010 138.600 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 136.200 42.230 138.600 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 136.200 45.910 138.600 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 136.200 49.130 138.600 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 136.200 52.810 138.600 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 136.200 56.030 138.600 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 136.200 59.710 138.600 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 136.200 62.930 138.600 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 136.200 66.150 138.600 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 136.200 69.830 138.600 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 136.200 8.190 138.600 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 136.200 11.870 138.600 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 136.200 15.090 138.600 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 136.200 18.770 138.600 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 136.200 21.990 138.600 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.930 136.200 25.210 138.600 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 136.200 28.890 138.600 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 136.200 32.110 138.600 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 136.200 35.790 138.600 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 136.200 73.050 138.600 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 136.200 107.090 138.600 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 136.200 110.770 138.600 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.710 136.200 113.990 138.600 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.390 136.200 117.670 138.600 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 136.200 120.890 138.600 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.830 136.200 124.110 138.600 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.510 136.200 127.790 138.600 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 136.200 131.010 138.600 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.410 136.200 134.690 138.600 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 136.200 137.910 138.600 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.450 136.200 76.730 138.600 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.670 136.200 79.950 138.600 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 136.200 83.170 138.600 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.570 136.200 86.850 138.600 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 136.200 90.070 138.600 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.470 136.200 93.750 138.600 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 136.200 96.970 138.600 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.370 136.200 100.650 138.600 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 136.200 103.870 138.600 ;
    END
  END chany_top_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 136.680 140.000 137.280 ;
    END
  END prog_clk
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 14.280 140.000 14.880 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 0.000 140.000 0.600 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 2.720 140.000 3.320 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 5.440 140.000 6.040 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 8.840 140.000 9.440 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 11.560 140.000 12.160 ;
    END
  END right_bottom_grid_pin_9_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 136.200 1.750 138.600 ;
    END
  END top_left_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 28.055 9.240 29.655 126.680 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.385 9.240 52.985 126.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 9.395 134.320 126.525 ;
      LAYER met1 ;
        RECT 1.450 9.240 137.930 135.920 ;
      LAYER met2 ;
        RECT 2.030 135.920 4.410 137.165 ;
        RECT 5.250 135.920 7.630 137.165 ;
        RECT 8.470 135.920 11.310 137.165 ;
        RECT 12.150 135.920 14.530 137.165 ;
        RECT 15.370 135.920 18.210 137.165 ;
        RECT 19.050 135.920 21.430 137.165 ;
        RECT 22.270 135.920 24.650 137.165 ;
        RECT 25.490 135.920 28.330 137.165 ;
        RECT 29.170 135.920 31.550 137.165 ;
        RECT 32.390 135.920 35.230 137.165 ;
        RECT 36.070 135.920 38.450 137.165 ;
        RECT 39.290 135.920 41.670 137.165 ;
        RECT 42.510 135.920 45.350 137.165 ;
        RECT 46.190 135.920 48.570 137.165 ;
        RECT 49.410 135.920 52.250 137.165 ;
        RECT 53.090 135.920 55.470 137.165 ;
        RECT 56.310 135.920 59.150 137.165 ;
        RECT 59.990 135.920 62.370 137.165 ;
        RECT 63.210 135.920 65.590 137.165 ;
        RECT 66.430 135.920 69.270 137.165 ;
        RECT 70.110 135.920 72.490 137.165 ;
        RECT 73.330 135.920 76.170 137.165 ;
        RECT 77.010 135.920 79.390 137.165 ;
        RECT 80.230 135.920 82.610 137.165 ;
        RECT 83.450 135.920 86.290 137.165 ;
        RECT 87.130 135.920 89.510 137.165 ;
        RECT 90.350 135.920 93.190 137.165 ;
        RECT 94.030 135.920 96.410 137.165 ;
        RECT 97.250 135.920 100.090 137.165 ;
        RECT 100.930 135.920 103.310 137.165 ;
        RECT 104.150 135.920 106.530 137.165 ;
        RECT 107.370 135.920 110.210 137.165 ;
        RECT 111.050 135.920 113.430 137.165 ;
        RECT 114.270 135.920 117.110 137.165 ;
        RECT 117.950 135.920 120.330 137.165 ;
        RECT 121.170 135.920 123.550 137.165 ;
        RECT 124.390 135.920 127.230 137.165 ;
        RECT 128.070 135.920 130.450 137.165 ;
        RECT 131.290 135.920 134.130 137.165 ;
        RECT 134.970 135.920 137.350 137.165 ;
        RECT 1.480 0.115 137.900 135.920 ;
      LAYER met3 ;
        RECT 2.365 136.280 137.200 137.145 ;
        RECT 2.365 134.960 137.600 136.280 ;
        RECT 2.365 133.560 137.200 134.960 ;
        RECT 2.365 131.560 137.600 133.560 ;
        RECT 2.365 130.160 137.200 131.560 ;
        RECT 2.365 128.840 137.600 130.160 ;
        RECT 2.365 127.440 137.200 128.840 ;
        RECT 2.365 126.120 137.600 127.440 ;
        RECT 2.365 124.720 137.200 126.120 ;
        RECT 2.365 122.720 137.600 124.720 ;
        RECT 2.365 121.320 137.200 122.720 ;
        RECT 2.365 120.000 137.600 121.320 ;
        RECT 2.365 118.600 137.200 120.000 ;
        RECT 2.365 116.600 137.600 118.600 ;
        RECT 2.365 115.200 137.200 116.600 ;
        RECT 2.365 113.880 137.600 115.200 ;
        RECT 2.365 112.480 137.200 113.880 ;
        RECT 2.365 111.160 137.600 112.480 ;
        RECT 2.365 109.760 137.200 111.160 ;
        RECT 2.365 107.760 137.600 109.760 ;
        RECT 2.365 106.360 137.200 107.760 ;
        RECT 2.365 105.040 137.600 106.360 ;
        RECT 2.365 104.360 137.200 105.040 ;
        RECT 2.800 103.640 137.200 104.360 ;
        RECT 2.800 102.960 137.600 103.640 ;
        RECT 2.365 102.320 137.600 102.960 ;
        RECT 2.365 100.920 137.200 102.320 ;
        RECT 2.365 98.920 137.600 100.920 ;
        RECT 2.365 97.520 137.200 98.920 ;
        RECT 2.365 96.200 137.600 97.520 ;
        RECT 2.365 94.800 137.200 96.200 ;
        RECT 2.365 92.800 137.600 94.800 ;
        RECT 2.365 91.400 137.200 92.800 ;
        RECT 2.365 90.080 137.600 91.400 ;
        RECT 2.365 88.680 137.200 90.080 ;
        RECT 2.365 87.360 137.600 88.680 ;
        RECT 2.365 85.960 137.200 87.360 ;
        RECT 2.365 83.960 137.600 85.960 ;
        RECT 2.365 82.560 137.200 83.960 ;
        RECT 2.365 81.240 137.600 82.560 ;
        RECT 2.365 79.840 137.200 81.240 ;
        RECT 2.365 77.840 137.600 79.840 ;
        RECT 2.365 76.440 137.200 77.840 ;
        RECT 2.365 75.120 137.600 76.440 ;
        RECT 2.365 73.720 137.200 75.120 ;
        RECT 2.365 72.400 137.600 73.720 ;
        RECT 2.365 71.000 137.200 72.400 ;
        RECT 2.365 69.000 137.600 71.000 ;
        RECT 2.365 67.600 137.200 69.000 ;
        RECT 2.365 66.280 137.600 67.600 ;
        RECT 2.365 64.880 137.200 66.280 ;
        RECT 2.365 63.560 137.600 64.880 ;
        RECT 2.365 62.160 137.200 63.560 ;
        RECT 2.365 60.160 137.600 62.160 ;
        RECT 2.365 58.760 137.200 60.160 ;
        RECT 2.365 57.440 137.600 58.760 ;
        RECT 2.365 56.040 137.200 57.440 ;
        RECT 2.365 54.040 137.600 56.040 ;
        RECT 2.365 52.640 137.200 54.040 ;
        RECT 2.365 51.320 137.600 52.640 ;
        RECT 2.365 49.920 137.200 51.320 ;
        RECT 2.365 48.600 137.600 49.920 ;
        RECT 2.365 47.200 137.200 48.600 ;
        RECT 2.365 45.200 137.600 47.200 ;
        RECT 2.365 43.800 137.200 45.200 ;
        RECT 2.365 42.480 137.600 43.800 ;
        RECT 2.365 41.080 137.200 42.480 ;
        RECT 2.365 39.080 137.600 41.080 ;
        RECT 2.365 37.680 137.200 39.080 ;
        RECT 2.365 36.360 137.600 37.680 ;
        RECT 2.365 34.960 137.200 36.360 ;
        RECT 2.365 34.320 137.600 34.960 ;
        RECT 2.800 33.640 137.600 34.320 ;
        RECT 2.800 32.920 137.200 33.640 ;
        RECT 2.365 32.240 137.200 32.920 ;
        RECT 2.365 30.240 137.600 32.240 ;
        RECT 2.365 28.840 137.200 30.240 ;
        RECT 2.365 27.520 137.600 28.840 ;
        RECT 2.365 26.120 137.200 27.520 ;
        RECT 2.365 24.800 137.600 26.120 ;
        RECT 2.365 23.400 137.200 24.800 ;
        RECT 2.365 21.400 137.600 23.400 ;
        RECT 2.365 20.000 137.200 21.400 ;
        RECT 2.365 18.680 137.600 20.000 ;
        RECT 2.365 17.280 137.200 18.680 ;
        RECT 2.365 15.280 137.600 17.280 ;
        RECT 2.365 13.880 137.200 15.280 ;
        RECT 2.365 12.560 137.600 13.880 ;
        RECT 2.365 11.160 137.200 12.560 ;
        RECT 2.365 9.840 137.600 11.160 ;
        RECT 2.365 8.440 137.200 9.840 ;
        RECT 2.365 6.440 137.600 8.440 ;
        RECT 2.365 5.040 137.200 6.440 ;
        RECT 2.365 3.720 137.600 5.040 ;
        RECT 2.365 2.320 137.200 3.720 ;
        RECT 2.365 1.000 137.600 2.320 ;
        RECT 2.365 0.135 137.200 1.000 ;
      LAYER met4 ;
        RECT 30.055 9.240 50.985 126.680 ;
        RECT 53.385 9.240 122.985 126.680 ;
  END
END sb_0__0_
END LIBRARY

