magic
tech EFS8A
magscale 1 2
timestamp 1602095416
<< locali >>
rect 2547 18785 2582 18819
rect 6371 16745 6377 16779
rect 11891 16745 11897 16779
rect 6371 16677 6405 16745
rect 11891 16677 11925 16745
rect 15243 16609 15370 16643
rect 6469 15895 6503 15997
rect 4439 14569 4445 14603
rect 4439 14501 4473 14569
rect 7843 13719 7877 13787
rect 7843 13685 7849 13719
rect 17635 12257 17670 12291
rect 12483 11645 12610 11679
rect 15209 11611 15243 11713
rect 15939 11305 15945 11339
rect 15939 11237 15973 11305
rect 4905 10523 4939 10761
rect 3427 10455 3461 10523
rect 3427 10421 3433 10455
rect 1547 10217 1685 10251
rect 6837 9979 6871 10149
rect 10051 9129 10057 9163
rect 10051 9061 10085 9129
rect 4387 7973 4432 8007
rect 14611 7497 14749 7531
rect 1972 6885 2040 6919
rect 5273 6103 5307 6409
rect 5687 6273 5825 6307
rect 12081 6103 12115 6205
rect 8251 5729 8286 5763
rect 9781 5151 9815 5321
rect 8217 4063 8251 4233
rect 5779 3145 5917 3179
rect 9597 2839 9631 3145
rect 6561 2499 6595 2601
<< viali >>
rect 10000 20961 10034 20995
rect 10103 20757 10137 20791
rect 4537 20553 4571 20587
rect 6101 20553 6135 20587
rect 7389 20553 7423 20587
rect 8953 20553 8987 20587
rect 9965 20553 9999 20587
rect 10977 20553 11011 20587
rect 14013 20553 14047 20587
rect 14749 20553 14783 20587
rect 16957 20553 16991 20587
rect 18613 20553 18647 20587
rect 21465 20553 21499 20587
rect 1444 20349 1478 20383
rect 1869 20349 1903 20383
rect 4144 20349 4178 20383
rect 5708 20349 5742 20383
rect 6904 20349 6938 20383
rect 8769 20349 8803 20383
rect 10492 20349 10526 20383
rect 13528 20349 13562 20383
rect 14565 20349 14599 20383
rect 15117 20349 15151 20383
rect 16472 20349 16506 20383
rect 18128 20349 18162 20383
rect 20980 20349 21014 20383
rect 1547 20213 1581 20247
rect 4215 20213 4249 20247
rect 5779 20213 5813 20247
rect 6975 20213 7009 20247
rect 9413 20213 9447 20247
rect 10563 20213 10597 20247
rect 13599 20213 13633 20247
rect 16543 20213 16577 20247
rect 18199 20213 18233 20247
rect 21051 20213 21085 20247
rect 1593 20009 1627 20043
rect 9827 20009 9861 20043
rect 10977 19941 11011 19975
rect 11069 19941 11103 19975
rect 12633 19941 12667 19975
rect 1409 19873 1443 19907
rect 2580 19873 2614 19907
rect 6101 19873 6135 19907
rect 9756 19873 9790 19907
rect 18036 19873 18070 19907
rect 12541 19805 12575 19839
rect 12817 19805 12851 19839
rect 11529 19737 11563 19771
rect 2651 19669 2685 19703
rect 6469 19669 6503 19703
rect 10149 19669 10183 19703
rect 18107 19669 18141 19703
rect 2973 19465 3007 19499
rect 6561 19465 6595 19499
rect 10241 19465 10275 19499
rect 12265 19465 12299 19499
rect 12909 19465 12943 19499
rect 19073 19465 19107 19499
rect 1593 19397 1627 19431
rect 5273 19329 5307 19363
rect 11529 19329 11563 19363
rect 13277 19329 13311 19363
rect 1409 19261 1443 19295
rect 4772 19261 4806 19295
rect 8953 19261 8987 19295
rect 9505 19261 9539 19295
rect 10701 19261 10735 19295
rect 11345 19261 11379 19295
rect 12516 19261 12550 19295
rect 18220 19261 18254 19295
rect 2421 19193 2455 19227
rect 4859 19193 4893 19227
rect 5733 19193 5767 19227
rect 6285 19193 6319 19227
rect 6929 19193 6963 19227
rect 7021 19193 7055 19227
rect 7573 19193 7607 19227
rect 9781 19193 9815 19227
rect 18705 19193 18739 19227
rect 1961 19125 1995 19159
rect 2513 19125 2547 19159
rect 5641 19125 5675 19159
rect 12587 19125 12621 19159
rect 18291 19125 18325 19159
rect 1593 18921 1627 18955
rect 2053 18921 2087 18955
rect 12449 18921 12483 18955
rect 6745 18853 6779 18887
rect 9873 18853 9907 18887
rect 12909 18853 12943 18887
rect 1409 18785 1443 18819
rect 2513 18785 2547 18819
rect 4353 18785 4387 18819
rect 20980 18785 21014 18819
rect 4077 18717 4111 18751
rect 6653 18717 6687 18751
rect 6929 18717 6963 18751
rect 8585 18717 8619 18751
rect 9781 18717 9815 18751
rect 10057 18717 10091 18751
rect 12817 18717 12851 18751
rect 13277 18717 13311 18751
rect 2421 18649 2455 18683
rect 2651 18581 2685 18615
rect 9413 18581 9447 18615
rect 10885 18581 10919 18615
rect 21051 18581 21085 18615
rect 4353 18377 4387 18411
rect 5043 18377 5077 18411
rect 6653 18377 6687 18411
rect 9137 18377 9171 18411
rect 10333 18377 10367 18411
rect 11897 18377 11931 18411
rect 21005 18377 21039 18411
rect 1777 18241 1811 18275
rect 3433 18241 3467 18275
rect 5917 18241 5951 18275
rect 6929 18241 6963 18275
rect 7573 18241 7607 18275
rect 9413 18241 9447 18275
rect 10057 18241 10091 18275
rect 12541 18241 12575 18275
rect 13185 18241 13219 18275
rect 4940 18173 4974 18207
rect 5365 18173 5399 18207
rect 1869 18105 1903 18139
rect 2421 18105 2455 18139
rect 3525 18105 3559 18139
rect 4077 18105 4111 18139
rect 6285 18105 6319 18139
rect 7021 18105 7055 18139
rect 9505 18105 9539 18139
rect 12633 18105 12667 18139
rect 2697 18037 2731 18071
rect 3249 18037 3283 18071
rect 12265 18037 12299 18071
rect 13461 18037 13495 18071
rect 3433 17833 3467 17867
rect 7297 17833 7331 17867
rect 8769 17833 8803 17867
rect 2329 17765 2363 17799
rect 4261 17765 4295 17799
rect 6469 17765 6503 17799
rect 7021 17765 7055 17799
rect 9873 17765 9907 17799
rect 12265 17765 12299 17799
rect 12909 17697 12943 17731
rect 2237 17629 2271 17663
rect 2513 17629 2547 17663
rect 4169 17629 4203 17663
rect 4445 17629 4479 17663
rect 6377 17629 6411 17663
rect 9781 17629 9815 17663
rect 10057 17629 10091 17663
rect 13829 17629 13863 17663
rect 1685 17493 1719 17527
rect 9321 17493 9355 17527
rect 3341 17289 3375 17323
rect 4721 17289 4755 17323
rect 12725 17289 12759 17323
rect 9413 17221 9447 17255
rect 1685 17153 1719 17187
rect 3801 17153 3835 17187
rect 6377 17153 6411 17187
rect 6837 17153 6871 17187
rect 8861 17153 8895 17187
rect 10241 17153 10275 17187
rect 12265 17153 12299 17187
rect 13001 17153 13035 17187
rect 1777 17085 1811 17119
rect 2697 17085 2731 17119
rect 6929 17085 6963 17119
rect 10793 17085 10827 17119
rect 11253 17085 11287 17119
rect 14381 17085 14415 17119
rect 14565 17085 14599 17119
rect 4122 17017 4156 17051
rect 8953 17017 8987 17051
rect 11529 17017 11563 17051
rect 13093 17017 13127 17051
rect 13645 17017 13679 17051
rect 14473 17017 14507 17051
rect 3617 16949 3651 16983
rect 4997 16949 5031 16983
rect 5917 16949 5951 16983
rect 8677 16949 8711 16983
rect 9781 16949 9815 16983
rect 10609 16949 10643 16983
rect 1777 16745 1811 16779
rect 2789 16745 2823 16779
rect 4169 16745 4203 16779
rect 6377 16745 6411 16779
rect 6929 16745 6963 16779
rect 7205 16745 7239 16779
rect 11897 16745 11931 16779
rect 12449 16745 12483 16779
rect 13001 16745 13035 16779
rect 2190 16677 2224 16711
rect 3157 16677 3191 16711
rect 9689 16677 9723 16711
rect 13461 16677 13495 16711
rect 4169 16609 4203 16643
rect 4629 16609 4663 16643
rect 8309 16609 8343 16643
rect 8493 16609 8527 16643
rect 9781 16609 9815 16643
rect 15209 16609 15243 16643
rect 1869 16541 1903 16575
rect 6009 16541 6043 16575
rect 8585 16541 8619 16575
rect 11529 16541 11563 16575
rect 13369 16541 13403 16575
rect 13645 16541 13679 16575
rect 3893 16405 3927 16439
rect 5825 16405 5859 16439
rect 10793 16405 10827 16439
rect 15439 16405 15473 16439
rect 1593 16201 1627 16235
rect 2421 16201 2455 16235
rect 8125 16201 8159 16235
rect 11253 16201 11287 16235
rect 13645 16201 13679 16235
rect 14013 16201 14047 16235
rect 15393 16201 15427 16235
rect 13369 16133 13403 16167
rect 5825 16065 5859 16099
rect 8401 16065 8435 16099
rect 8585 16065 8619 16099
rect 1409 15997 1443 16031
rect 2881 15997 2915 16031
rect 3617 15997 3651 16031
rect 5089 15997 5123 16031
rect 5457 15997 5491 16031
rect 5733 15997 5767 16031
rect 6469 15997 6503 16031
rect 6837 15997 6871 16031
rect 7297 15997 7331 16031
rect 9781 15997 9815 16031
rect 10333 15997 10367 16031
rect 12449 15997 12483 16031
rect 14248 15997 14282 16031
rect 14657 15997 14691 16031
rect 2973 15929 3007 15963
rect 8906 15929 8940 15963
rect 10149 15929 10183 15963
rect 10654 15929 10688 15963
rect 11529 15929 11563 15963
rect 12173 15929 12207 15963
rect 12770 15929 12804 15963
rect 14335 15929 14369 15963
rect 2053 15861 2087 15895
rect 4077 15861 4111 15895
rect 4537 15861 4571 15895
rect 6285 15861 6319 15895
rect 6469 15861 6503 15895
rect 6561 15861 6595 15895
rect 6929 15861 6963 15895
rect 9505 15861 9539 15895
rect 1961 15657 1995 15691
rect 4169 15657 4203 15691
rect 5273 15657 5307 15691
rect 6837 15657 6871 15691
rect 9045 15657 9079 15691
rect 9873 15657 9907 15691
rect 11897 15657 11931 15691
rect 14657 15657 14691 15691
rect 2421 15589 2455 15623
rect 6279 15589 6313 15623
rect 8769 15589 8803 15623
rect 10333 15589 10367 15623
rect 11621 15589 11655 15623
rect 12817 15589 12851 15623
rect 13829 15589 13863 15623
rect 4353 15521 4387 15555
rect 4537 15521 4571 15555
rect 5917 15521 5951 15555
rect 8033 15521 8067 15555
rect 8585 15521 8619 15555
rect 10885 15521 10919 15555
rect 11345 15521 11379 15555
rect 2329 15453 2363 15487
rect 2973 15453 3007 15487
rect 13737 15453 13771 15487
rect 7113 15385 7147 15419
rect 14289 15385 14323 15419
rect 1685 15317 1719 15351
rect 10701 15317 10735 15351
rect 12449 15317 12483 15351
rect 2881 15113 2915 15147
rect 3893 15113 3927 15147
rect 5457 15113 5491 15147
rect 10241 15113 10275 15147
rect 11345 15113 11379 15147
rect 12173 15113 12207 15147
rect 13369 15113 13403 15147
rect 13737 15113 13771 15147
rect 3525 15045 3559 15079
rect 4629 15045 4663 15079
rect 1869 14977 1903 15011
rect 2329 14977 2363 15011
rect 4077 14977 4111 15011
rect 5687 14977 5721 15011
rect 14289 14977 14323 15011
rect 14565 14977 14599 15011
rect 5600 14909 5634 14943
rect 6009 14909 6043 14943
rect 9965 14909 9999 14943
rect 10425 14909 10459 14943
rect 12449 14909 12483 14943
rect 18832 14909 18866 14943
rect 19257 14909 19291 14943
rect 1685 14841 1719 14875
rect 1961 14841 1995 14875
rect 4169 14841 4203 14875
rect 10746 14841 10780 14875
rect 11621 14841 11655 14875
rect 12770 14841 12804 14875
rect 14381 14841 14415 14875
rect 4997 14773 5031 14807
rect 6377 14773 6411 14807
rect 8033 14773 8067 14807
rect 8493 14773 8527 14807
rect 14105 14773 14139 14807
rect 18935 14773 18969 14807
rect 2697 14569 2731 14603
rect 3157 14569 3191 14603
rect 4445 14569 4479 14603
rect 4997 14569 5031 14603
rect 10333 14569 10367 14603
rect 14473 14569 14507 14603
rect 19901 14569 19935 14603
rect 1869 14501 1903 14535
rect 3893 14501 3927 14535
rect 6279 14501 6313 14535
rect 12357 14501 12391 14535
rect 14105 14501 14139 14535
rect 16773 14501 16807 14535
rect 10149 14433 10183 14467
rect 10517 14433 10551 14467
rect 11897 14433 11931 14467
rect 12173 14433 12207 14467
rect 13737 14433 13771 14467
rect 18797 14433 18831 14467
rect 19717 14433 19751 14467
rect 1777 14365 1811 14399
rect 4077 14365 4111 14399
rect 5917 14365 5951 14399
rect 8401 14365 8435 14399
rect 9965 14365 9999 14399
rect 16681 14365 16715 14399
rect 17325 14365 17359 14399
rect 2329 14297 2363 14331
rect 6837 14297 6871 14331
rect 11437 14297 11471 14331
rect 11069 14229 11103 14263
rect 12817 14229 12851 14263
rect 15485 14229 15519 14263
rect 18429 14229 18463 14263
rect 1869 14025 1903 14059
rect 2605 14025 2639 14059
rect 3709 14025 3743 14059
rect 6561 14025 6595 14059
rect 11069 14025 11103 14059
rect 12173 14025 12207 14059
rect 13737 14025 13771 14059
rect 16773 14025 16807 14059
rect 19073 14025 19107 14059
rect 20085 14025 20119 14059
rect 5503 13957 5537 13991
rect 10333 13957 10367 13991
rect 17049 13957 17083 13991
rect 9321 13889 9355 13923
rect 10701 13889 10735 13923
rect 11161 13889 11195 13923
rect 11897 13889 11931 13923
rect 15485 13889 15519 13923
rect 2237 13821 2271 13855
rect 3801 13821 3835 13855
rect 4353 13821 4387 13855
rect 5432 13821 5466 13855
rect 5825 13821 5859 13855
rect 7481 13821 7515 13855
rect 10793 13821 10827 13855
rect 10940 13821 10974 13855
rect 12817 13821 12851 13855
rect 9413 13753 9447 13787
rect 9965 13753 9999 13787
rect 15806 13753 15840 13787
rect 17509 13753 17543 13787
rect 18153 13753 18187 13787
rect 18245 13753 18279 13787
rect 18797 13753 18831 13787
rect 19625 13753 19659 13787
rect 3341 13685 3375 13719
rect 4077 13685 4111 13719
rect 4905 13685 4939 13719
rect 6285 13685 6319 13719
rect 7389 13685 7423 13719
rect 7849 13685 7883 13719
rect 8401 13685 8435 13719
rect 9045 13685 9079 13719
rect 11437 13685 11471 13719
rect 13185 13685 13219 13719
rect 15393 13685 15427 13719
rect 16405 13685 16439 13719
rect 17877 13685 17911 13719
rect 1777 13481 1811 13515
rect 3249 13481 3283 13515
rect 4169 13481 4203 13515
rect 6101 13481 6135 13515
rect 7481 13481 7515 13515
rect 9321 13481 9355 13515
rect 11529 13481 11563 13515
rect 13001 13481 13035 13515
rect 13369 13481 13403 13515
rect 16405 13481 16439 13515
rect 2237 13413 2271 13447
rect 2329 13413 2363 13447
rect 12402 13413 12436 13447
rect 15847 13413 15881 13447
rect 17969 13413 18003 13447
rect 18521 13413 18555 13447
rect 4353 13345 4387 13379
rect 4629 13345 4663 13379
rect 6101 13345 6135 13379
rect 6561 13345 6595 13379
rect 8125 13345 8159 13379
rect 10517 13345 10551 13379
rect 11069 13345 11103 13379
rect 2513 13277 2547 13311
rect 11253 13277 11287 13311
rect 12081 13277 12115 13311
rect 13829 13277 13863 13311
rect 15485 13277 15519 13311
rect 17877 13277 17911 13311
rect 3893 13141 3927 13175
rect 7113 13141 7147 13175
rect 8493 13141 8527 13175
rect 10241 13141 10275 13175
rect 3341 12937 3375 12971
rect 4629 12937 4663 12971
rect 8125 12937 8159 12971
rect 8493 12937 8527 12971
rect 10314 12937 10348 12971
rect 10793 12937 10827 12971
rect 11529 12937 11563 12971
rect 12081 12937 12115 12971
rect 12633 12937 12667 12971
rect 13001 12937 13035 12971
rect 16313 12937 16347 12971
rect 17417 12937 17451 12971
rect 4077 12869 4111 12903
rect 4445 12869 4479 12903
rect 10425 12869 10459 12903
rect 18705 12869 18739 12903
rect 19441 12869 19475 12903
rect 3709 12801 3743 12835
rect 4537 12801 4571 12835
rect 7481 12801 7515 12835
rect 8677 12801 8711 12835
rect 10517 12801 10551 12835
rect 13277 12801 13311 12835
rect 13737 12801 13771 12835
rect 15393 12801 15427 12835
rect 18153 12801 18187 12835
rect 19073 12801 19107 12835
rect 1869 12733 1903 12767
rect 4316 12733 4350 12767
rect 5641 12733 5675 12767
rect 6837 12733 6871 12767
rect 7297 12733 7331 12767
rect 9321 12733 9355 12767
rect 14657 12733 14691 12767
rect 14749 12733 14783 12767
rect 15209 12733 15243 12767
rect 16773 12733 16807 12767
rect 1777 12665 1811 12699
rect 2190 12665 2224 12699
rect 4169 12665 4203 12699
rect 8769 12665 8803 12699
rect 10149 12665 10183 12699
rect 13369 12665 13403 12699
rect 17141 12665 17175 12699
rect 17785 12665 17819 12699
rect 18245 12665 18279 12699
rect 2789 12597 2823 12631
rect 5273 12597 5307 12631
rect 5733 12597 5767 12631
rect 6193 12597 6227 12631
rect 6561 12597 6595 12631
rect 9597 12597 9631 12631
rect 10057 12597 10091 12631
rect 11161 12597 11195 12631
rect 15853 12597 15887 12631
rect 3157 12393 3191 12427
rect 3893 12393 3927 12427
rect 7941 12393 7975 12427
rect 8677 12393 8711 12427
rect 10701 12393 10735 12427
rect 11069 12393 11103 12427
rect 12633 12393 12667 12427
rect 14749 12393 14783 12427
rect 15577 12393 15611 12427
rect 16313 12393 16347 12427
rect 17739 12393 17773 12427
rect 21097 12393 21131 12427
rect 1869 12325 1903 12359
rect 4077 12325 4111 12359
rect 8033 12325 8067 12359
rect 13093 12325 13127 12359
rect 13645 12325 13679 12359
rect 18797 12325 18831 12359
rect 2789 12257 2823 12291
rect 4629 12257 4663 12291
rect 6377 12257 6411 12291
rect 10057 12257 10091 12291
rect 11688 12257 11722 12291
rect 12081 12257 12115 12291
rect 15301 12257 15335 12291
rect 15761 12257 15795 12291
rect 17601 12257 17635 12291
rect 20913 12257 20947 12291
rect 1777 12189 1811 12223
rect 6745 12189 6779 12223
rect 8180 12189 8214 12223
rect 8401 12189 8435 12223
rect 10425 12189 10459 12223
rect 13001 12189 13035 12223
rect 18705 12189 18739 12223
rect 18981 12189 19015 12223
rect 2329 12121 2363 12155
rect 5917 12121 5951 12155
rect 6837 12121 6871 12155
rect 11759 12121 11793 12155
rect 5273 12053 5307 12087
rect 6193 12053 6227 12087
rect 6515 12053 6549 12087
rect 6653 12053 6687 12087
rect 7389 12053 7423 12087
rect 8309 12053 8343 12087
rect 9137 12053 9171 12087
rect 9873 12053 9907 12087
rect 10195 12053 10229 12087
rect 10333 12053 10367 12087
rect 14013 12053 14047 12087
rect 18337 12053 18371 12087
rect 2053 11849 2087 11883
rect 4629 11849 4663 11883
rect 10425 11849 10459 11883
rect 10609 11849 10643 11883
rect 11161 11849 11195 11883
rect 11529 11849 11563 11883
rect 13369 11849 13403 11883
rect 15301 11849 15335 11883
rect 16681 11849 16715 11883
rect 1593 11781 1627 11815
rect 3617 11781 3651 11815
rect 6377 11781 6411 11815
rect 8493 11781 8527 11815
rect 10287 11781 10321 11815
rect 13093 11781 13127 11815
rect 16405 11781 16439 11815
rect 20959 11781 20993 11815
rect 21649 11781 21683 11815
rect 3985 11713 4019 11747
rect 7205 11713 7239 11747
rect 9321 11713 9355 11747
rect 10517 11713 10551 11747
rect 12679 11713 12713 11747
rect 14933 11713 14967 11747
rect 15209 11713 15243 11747
rect 18981 11713 19015 11747
rect 21281 11713 21315 11747
rect 1409 11645 1443 11679
rect 5457 11645 5491 11679
rect 5641 11645 5675 11679
rect 8677 11645 8711 11679
rect 9597 11645 9631 11679
rect 12449 11645 12483 11679
rect 13921 11645 13955 11679
rect 14381 11645 14415 11679
rect 14657 11645 14691 11679
rect 15485 11645 15519 11679
rect 17049 11645 17083 11679
rect 20856 11645 20890 11679
rect 2697 11577 2731 11611
rect 2789 11577 2823 11611
rect 3341 11577 3375 11611
rect 5917 11577 5951 11611
rect 6929 11577 6963 11611
rect 7021 11577 7055 11611
rect 10149 11577 10183 11611
rect 11897 11577 11931 11611
rect 15209 11577 15243 11611
rect 15806 11577 15840 11611
rect 18337 11577 18371 11611
rect 18429 11577 18463 11611
rect 19809 11577 19843 11611
rect 2513 11509 2547 11543
rect 4169 11509 4203 11543
rect 5089 11509 5123 11543
rect 8125 11509 8159 11543
rect 9965 11509 9999 11543
rect 13737 11509 13771 11543
rect 17693 11509 17727 11543
rect 19349 11509 19383 11543
rect 1547 11305 1581 11339
rect 4997 11305 5031 11339
rect 6837 11305 6871 11339
rect 8217 11305 8251 11339
rect 10425 11305 10459 11339
rect 15945 11305 15979 11339
rect 18705 11305 18739 11339
rect 19441 11305 19475 11339
rect 1961 11237 1995 11271
rect 2605 11237 2639 11271
rect 6238 11237 6272 11271
rect 8493 11237 8527 11271
rect 10793 11237 10827 11271
rect 11707 11237 11741 11271
rect 13277 11237 13311 11271
rect 17785 11237 17819 11271
rect 18337 11237 18371 11271
rect 18981 11237 19015 11271
rect 1476 11169 1510 11203
rect 4353 11169 4387 11203
rect 5733 11169 5767 11203
rect 7700 11169 7734 11203
rect 9781 11169 9815 11203
rect 19257 11169 19291 11203
rect 20913 11169 20947 11203
rect 2513 11101 2547 11135
rect 2973 11101 3007 11135
rect 4721 11101 4755 11135
rect 5917 11101 5951 11135
rect 9928 11101 9962 11135
rect 10149 11101 10183 11135
rect 11345 11101 11379 11135
rect 13185 11101 13219 11135
rect 13461 11101 13495 11135
rect 15577 11101 15611 11135
rect 17693 11101 17727 11135
rect 7481 11033 7515 11067
rect 2237 10965 2271 10999
rect 4518 10965 4552 10999
rect 4629 10965 4663 10999
rect 5457 10965 5491 10999
rect 7113 10965 7147 10999
rect 7803 10965 7837 10999
rect 8861 10965 8895 10999
rect 9505 10965 9539 10999
rect 10057 10965 10091 10999
rect 12265 10965 12299 10999
rect 12725 10965 12759 10999
rect 16497 10965 16531 10999
rect 21097 10965 21131 10999
rect 1961 10761 1995 10795
rect 2973 10761 3007 10795
rect 4353 10761 4387 10795
rect 4905 10761 4939 10795
rect 6009 10761 6043 10795
rect 7941 10761 7975 10795
rect 9413 10761 9447 10795
rect 10149 10761 10183 10795
rect 11529 10761 11563 10795
rect 13645 10761 13679 10795
rect 15761 10761 15795 10795
rect 17417 10761 17451 10795
rect 19165 10761 19199 10795
rect 20913 10761 20947 10795
rect 1593 10693 1627 10727
rect 2513 10693 2547 10727
rect 3985 10693 4019 10727
rect 4813 10625 4847 10659
rect 1409 10557 1443 10591
rect 3065 10557 3099 10591
rect 5135 10693 5169 10727
rect 5273 10693 5307 10727
rect 8566 10693 8600 10727
rect 8677 10693 8711 10727
rect 17141 10693 17175 10727
rect 5365 10625 5399 10659
rect 8309 10625 8343 10659
rect 8769 10625 8803 10659
rect 11161 10625 11195 10659
rect 11805 10625 11839 10659
rect 12725 10625 12759 10659
rect 13369 10625 13403 10659
rect 14565 10625 14599 10659
rect 15393 10625 15427 10659
rect 16037 10625 16071 10659
rect 18429 10625 18463 10659
rect 6837 10557 6871 10591
rect 7021 10557 7055 10591
rect 10517 10557 10551 10591
rect 10885 10557 10919 10591
rect 14933 10557 14967 10591
rect 15117 10557 15151 10591
rect 4905 10489 4939 10523
rect 4997 10489 5031 10523
rect 8401 10489 8435 10523
rect 12265 10489 12299 10523
rect 12817 10489 12851 10523
rect 18153 10489 18187 10523
rect 18245 10489 18279 10523
rect 3433 10421 3467 10455
rect 5641 10421 5675 10455
rect 6377 10421 6411 10455
rect 9045 10421 9079 10455
rect 9781 10421 9815 10455
rect 17785 10421 17819 10455
rect 1685 10217 1719 10251
rect 2237 10217 2271 10251
rect 3433 10217 3467 10251
rect 4537 10217 4571 10251
rect 5549 10217 5583 10251
rect 7021 10217 7055 10251
rect 7389 10217 7423 10251
rect 9045 10217 9079 10251
rect 9413 10217 9447 10251
rect 9965 10217 9999 10251
rect 11069 10217 11103 10251
rect 12541 10217 12575 10251
rect 13277 10217 13311 10251
rect 14657 10217 14691 10251
rect 2605 10149 2639 10183
rect 3157 10149 3191 10183
rect 4261 10149 4295 10183
rect 6745 10149 6779 10183
rect 6837 10149 6871 10183
rect 7941 10149 7975 10183
rect 17785 10149 17819 10183
rect 1476 10081 1510 10115
rect 4721 10081 4755 10115
rect 4905 10081 4939 10115
rect 6009 10081 6043 10115
rect 2513 10013 2547 10047
rect 6377 10013 6411 10047
rect 8309 10081 8343 10115
rect 8493 10081 8527 10115
rect 9781 10081 9815 10115
rect 12357 10081 12391 10115
rect 13864 10081 13898 10115
rect 17417 10081 17451 10115
rect 8769 10013 8803 10047
rect 1961 9945 1995 9979
rect 6174 9945 6208 9979
rect 6837 9945 6871 9979
rect 3893 9877 3927 9911
rect 5825 9877 5859 9911
rect 6285 9877 6319 9911
rect 10793 9877 10827 9911
rect 13967 9877 14001 9911
rect 18061 9877 18095 9911
rect 2145 9673 2179 9707
rect 4445 9673 4479 9707
rect 4813 9673 4847 9707
rect 6193 9673 6227 9707
rect 6469 9673 6503 9707
rect 8493 9673 8527 9707
rect 12909 9673 12943 9707
rect 13829 9673 13863 9707
rect 17003 9673 17037 9707
rect 1593 9605 1627 9639
rect 8125 9605 8159 9639
rect 17693 9605 17727 9639
rect 2513 9537 2547 9571
rect 2697 9537 2731 9571
rect 9413 9537 9447 9571
rect 12449 9537 12483 9571
rect 1409 9469 1443 9503
rect 2881 9469 2915 9503
rect 5733 9469 5767 9503
rect 7205 9469 7239 9503
rect 16932 9469 16966 9503
rect 7113 9401 7147 9435
rect 7567 9401 7601 9435
rect 8769 9401 8803 9435
rect 10149 9401 10183 9435
rect 10241 9401 10275 9435
rect 10793 9401 10827 9435
rect 5365 9333 5399 9367
rect 9689 9333 9723 9367
rect 11069 9333 11103 9367
rect 17417 9333 17451 9367
rect 2789 9129 2823 9163
rect 3065 9129 3099 9163
rect 4215 9129 4249 9163
rect 4997 9129 5031 9163
rect 6469 9129 6503 9163
rect 7205 9129 7239 9163
rect 7481 9129 7515 9163
rect 10057 9129 10091 9163
rect 10609 9129 10643 9163
rect 5273 9061 5307 9095
rect 5825 9061 5859 9095
rect 1961 8993 1995 9027
rect 4144 8993 4178 9027
rect 4537 8993 4571 9027
rect 7665 8993 7699 9027
rect 7849 8993 7883 9027
rect 9689 8993 9723 9027
rect 13737 8993 13771 9027
rect 5181 8925 5215 8959
rect 13645 8925 13679 8959
rect 1777 8789 1811 8823
rect 6101 8789 6135 8823
rect 10885 8789 10919 8823
rect 5089 8585 5123 8619
rect 6653 8585 6687 8619
rect 9229 8585 9263 8619
rect 9965 8585 9999 8619
rect 2237 8449 2271 8483
rect 5273 8449 5307 8483
rect 5917 8449 5951 8483
rect 9413 8449 9447 8483
rect 10517 8449 10551 8483
rect 3433 8381 3467 8415
rect 3801 8381 3835 8415
rect 3985 8381 4019 8415
rect 6285 8381 6319 8415
rect 7113 8381 7147 8415
rect 1593 8313 1627 8347
rect 1685 8313 1719 8347
rect 5365 8313 5399 8347
rect 10609 8313 10643 8347
rect 11161 8313 11195 8347
rect 2605 8245 2639 8279
rect 2881 8245 2915 8279
rect 3801 8245 3835 8279
rect 4721 8245 4755 8279
rect 7297 8245 7331 8279
rect 8125 8245 8159 8279
rect 10333 8245 10367 8279
rect 13737 8245 13771 8279
rect 1685 8041 1719 8075
rect 2789 8041 2823 8075
rect 3617 8041 3651 8075
rect 4997 8041 5031 8075
rect 5641 8041 5675 8075
rect 10333 8041 10367 8075
rect 1961 7973 1995 8007
rect 2513 7973 2547 8007
rect 4353 7973 4387 8007
rect 7297 7973 7331 8007
rect 4077 7905 4111 7939
rect 10241 7905 10275 7939
rect 11897 7905 11931 7939
rect 12081 7905 12115 7939
rect 19292 7905 19326 7939
rect 1869 7837 1903 7871
rect 3157 7837 3191 7871
rect 6101 7837 6135 7871
rect 7205 7837 7239 7871
rect 7849 7837 7883 7871
rect 12357 7837 12391 7871
rect 5273 7701 5307 7735
rect 6837 7701 6871 7735
rect 8677 7701 8711 7735
rect 12909 7701 12943 7735
rect 19395 7701 19429 7735
rect 2881 7497 2915 7531
rect 4077 7497 4111 7531
rect 5871 7497 5905 7531
rect 6285 7497 6319 7531
rect 7757 7497 7791 7531
rect 10057 7497 10091 7531
rect 11713 7497 11747 7531
rect 12081 7497 12115 7531
rect 14749 7497 14783 7531
rect 19257 7497 19291 7531
rect 21465 7497 21499 7531
rect 2145 7429 2179 7463
rect 4307 7429 4341 7463
rect 4445 7429 4479 7463
rect 4537 7361 4571 7395
rect 8677 7361 8711 7395
rect 13461 7361 13495 7395
rect 3100 7293 3134 7327
rect 5800 7293 5834 7327
rect 6837 7293 6871 7327
rect 9689 7293 9723 7327
rect 10241 7293 10275 7327
rect 14540 7293 14574 7327
rect 14933 7293 14967 7327
rect 20980 7293 21014 7327
rect 1593 7225 1627 7259
rect 1685 7225 1719 7259
rect 4169 7225 4203 7259
rect 6561 7225 6595 7259
rect 7158 7225 7192 7259
rect 8769 7225 8803 7259
rect 9321 7225 9355 7259
rect 10149 7225 10183 7259
rect 13001 7225 13035 7259
rect 13093 7225 13127 7259
rect 2513 7157 2547 7191
rect 3203 7157 3237 7191
rect 3709 7157 3743 7191
rect 4813 7157 4847 7191
rect 5181 7157 5215 7191
rect 5641 7157 5675 7191
rect 8493 7157 8527 7191
rect 12817 7157 12851 7191
rect 21051 7157 21085 7191
rect 2881 6953 2915 6987
rect 3525 6953 3559 6987
rect 4169 6953 4203 6987
rect 6837 6953 6871 6987
rect 7297 6953 7331 6987
rect 11713 6953 11747 6987
rect 12449 6953 12483 6987
rect 1938 6885 1972 6919
rect 5825 6885 5859 6919
rect 7941 6885 7975 6919
rect 8033 6885 8067 6919
rect 9873 6885 9907 6919
rect 12909 6885 12943 6919
rect 13461 6885 13495 6919
rect 1685 6817 1719 6851
rect 4353 6817 4387 6851
rect 4537 6817 4571 6851
rect 6193 6817 6227 6851
rect 6745 6817 6779 6851
rect 6929 6817 6963 6851
rect 8217 6749 8251 6783
rect 9781 6749 9815 6783
rect 12817 6749 12851 6783
rect 10333 6681 10367 6715
rect 2605 6613 2639 6647
rect 3893 6613 3927 6647
rect 7665 6613 7699 6647
rect 3433 6409 3467 6443
rect 3801 6409 3835 6443
rect 5273 6409 5307 6443
rect 5457 6409 5491 6443
rect 6377 6409 6411 6443
rect 9137 6409 9171 6443
rect 10517 6409 10551 6443
rect 2145 6341 2179 6375
rect 4077 6341 4111 6375
rect 4261 6205 4295 6239
rect 4537 6205 4571 6239
rect 1593 6137 1627 6171
rect 1685 6137 1719 6171
rect 5089 6137 5123 6171
rect 5825 6273 5859 6307
rect 11253 6273 11287 6307
rect 12449 6273 12483 6307
rect 13645 6273 13679 6307
rect 5616 6205 5650 6239
rect 6009 6205 6043 6239
rect 7757 6205 7791 6239
rect 8125 6205 8159 6239
rect 8493 6205 8527 6239
rect 8769 6205 8803 6239
rect 9597 6205 9631 6239
rect 10793 6205 10827 6239
rect 12081 6205 12115 6239
rect 14197 6205 14231 6239
rect 14381 6205 14415 6239
rect 14841 6205 14875 6239
rect 9505 6137 9539 6171
rect 9959 6137 9993 6171
rect 11897 6137 11931 6171
rect 12770 6137 12804 6171
rect 15117 6137 15151 6171
rect 2513 6069 2547 6103
rect 2881 6069 2915 6103
rect 5273 6069 5307 6103
rect 7021 6069 7055 6103
rect 7481 6069 7515 6103
rect 12081 6069 12115 6103
rect 12173 6069 12207 6103
rect 13369 6069 13403 6103
rect 2421 5865 2455 5899
rect 2973 5865 3007 5899
rect 3893 5865 3927 5899
rect 8033 5865 8067 5899
rect 8769 5865 8803 5899
rect 12817 5865 12851 5899
rect 14473 5865 14507 5899
rect 15577 5865 15611 5899
rect 2145 5797 2179 5831
rect 5089 5797 5123 5831
rect 1961 5729 1995 5763
rect 4353 5729 4387 5763
rect 6009 5729 6043 5763
rect 8217 5729 8251 5763
rect 10057 5729 10091 5763
rect 10204 5729 10238 5763
rect 12633 5729 12667 5763
rect 4721 5661 4755 5695
rect 7757 5661 7791 5695
rect 10425 5661 10459 5695
rect 10793 5661 10827 5695
rect 2789 5593 2823 5627
rect 4629 5593 4663 5627
rect 8355 5593 8389 5627
rect 10333 5593 10367 5627
rect 4491 5525 4525 5559
rect 5365 5525 5399 5559
rect 5733 5525 5767 5559
rect 6193 5525 6227 5559
rect 9873 5525 9907 5559
rect 2973 5321 3007 5355
rect 4537 5321 4571 5355
rect 6009 5321 6043 5355
rect 6469 5321 6503 5355
rect 9781 5321 9815 5355
rect 9965 5321 9999 5355
rect 10333 5321 10367 5355
rect 10701 5321 10735 5355
rect 12265 5321 12299 5355
rect 5273 5253 5307 5287
rect 2605 5185 2639 5219
rect 4169 5185 4203 5219
rect 5365 5185 5399 5219
rect 9505 5185 9539 5219
rect 10195 5253 10229 5287
rect 11069 5253 11103 5287
rect 11437 5253 11471 5287
rect 10425 5185 10459 5219
rect 15577 5185 15611 5219
rect 2237 5117 2271 5151
rect 3341 5117 3375 5151
rect 3525 5117 3559 5151
rect 4997 5117 5031 5151
rect 5144 5117 5178 5151
rect 6872 5117 6906 5151
rect 7297 5117 7331 5151
rect 7757 5117 7791 5151
rect 8585 5117 8619 5151
rect 9781 5117 9815 5151
rect 12484 5117 12518 5151
rect 12909 5117 12943 5151
rect 13553 5117 13587 5151
rect 13645 5117 13679 5151
rect 14197 5117 14231 5151
rect 1961 5049 1995 5083
rect 2053 5049 2087 5083
rect 6975 5049 7009 5083
rect 8953 5049 8987 5083
rect 10057 5049 10091 5083
rect 11805 5049 11839 5083
rect 12587 5049 12621 5083
rect 14381 5049 14415 5083
rect 15898 5049 15932 5083
rect 4813 4981 4847 5015
rect 5641 4981 5675 5015
rect 8125 4981 8159 5015
rect 15393 4981 15427 5015
rect 16497 4981 16531 5015
rect 1961 4777 1995 4811
rect 4353 4777 4387 4811
rect 5549 4777 5583 4811
rect 6009 4777 6043 4811
rect 7113 4777 7147 4811
rect 13231 4777 13265 4811
rect 13737 4777 13771 4811
rect 14289 4777 14323 4811
rect 2329 4709 2363 4743
rect 6285 4709 6319 4743
rect 9505 4709 9539 4743
rect 10793 4709 10827 4743
rect 11707 4709 11741 4743
rect 17325 4709 17359 4743
rect 1476 4641 1510 4675
rect 2697 4641 2731 4675
rect 2973 4641 3007 4675
rect 4537 4641 4571 4675
rect 5089 4641 5123 4675
rect 7665 4641 7699 4675
rect 8217 4641 8251 4675
rect 8493 4641 8527 4675
rect 10057 4641 10091 4675
rect 10333 4641 10367 4675
rect 12541 4641 12575 4675
rect 13160 4641 13194 4675
rect 15945 4641 15979 4675
rect 3157 4573 3191 4607
rect 5273 4573 5307 4607
rect 6193 4573 6227 4607
rect 10517 4573 10551 4607
rect 11345 4573 11379 4607
rect 17233 4573 17267 4607
rect 17877 4573 17911 4607
rect 1547 4505 1581 4539
rect 6745 4505 6779 4539
rect 7481 4437 7515 4471
rect 8769 4437 8803 4471
rect 12265 4437 12299 4471
rect 15577 4437 15611 4471
rect 18153 4437 18187 4471
rect 1593 4233 1627 4267
rect 3249 4233 3283 4267
rect 4905 4233 4939 4267
rect 5365 4233 5399 4267
rect 8217 4233 8251 4267
rect 10701 4233 10735 4267
rect 11161 4233 11195 4267
rect 11805 4233 11839 4267
rect 17233 4233 17267 4267
rect 3709 4097 3743 4131
rect 6653 4097 6687 4131
rect 7757 4097 7791 4131
rect 14013 4165 14047 4199
rect 15117 4165 15151 4199
rect 15485 4165 15519 4199
rect 15853 4165 15887 4199
rect 9137 4097 9171 4131
rect 10425 4097 10459 4131
rect 12541 4097 12575 4131
rect 12817 4097 12851 4131
rect 14197 4097 14231 4131
rect 16313 4097 16347 4131
rect 18429 4097 18463 4131
rect 2513 4029 2547 4063
rect 2881 4029 2915 4063
rect 5492 4029 5526 4063
rect 5917 4029 5951 4063
rect 7021 4029 7055 4063
rect 7849 4029 7883 4063
rect 8217 4029 8251 4063
rect 11380 4029 11414 4063
rect 2329 3961 2363 3995
rect 4030 3961 4064 3995
rect 8401 3961 8435 3995
rect 9458 3961 9492 3995
rect 12265 3961 12299 3995
rect 12633 3961 12667 3995
rect 14518 3961 14552 3995
rect 16037 3961 16071 3995
rect 16129 3961 16163 3995
rect 18153 3961 18187 3995
rect 18245 3961 18279 3995
rect 2145 3893 2179 3927
rect 3525 3893 3559 3927
rect 4629 3893 4663 3927
rect 5595 3893 5629 3927
rect 7297 3893 7331 3927
rect 8953 3893 8987 3927
rect 10057 3893 10091 3927
rect 11483 3893 11517 3927
rect 13461 3893 13495 3927
rect 17785 3893 17819 3927
rect 3709 3689 3743 3723
rect 4629 3689 4663 3723
rect 6193 3689 6227 3723
rect 7481 3689 7515 3723
rect 8493 3689 8527 3723
rect 9137 3689 9171 3723
rect 17877 3689 17911 3723
rect 5594 3621 5628 3655
rect 7894 3621 7928 3655
rect 10149 3621 10183 3655
rect 12081 3621 12115 3655
rect 12633 3621 12667 3655
rect 13461 3621 13495 3655
rect 15485 3621 15519 3655
rect 16037 3621 16071 3655
rect 17601 3621 17635 3655
rect 2237 3553 2271 3587
rect 2789 3553 2823 3587
rect 3065 3553 3099 3587
rect 4144 3553 4178 3587
rect 5273 3553 5307 3587
rect 7573 3553 7607 3587
rect 8769 3553 8803 3587
rect 13553 3553 13587 3587
rect 17325 3553 17359 3587
rect 7021 3485 7055 3519
rect 10057 3485 10091 3519
rect 11989 3485 12023 3519
rect 15393 3485 15427 3519
rect 16405 3485 16439 3519
rect 10609 3417 10643 3451
rect 1961 3349 1995 3383
rect 4215 3349 4249 3383
rect 6469 3349 6503 3383
rect 11345 3349 11379 3383
rect 1547 3145 1581 3179
rect 5365 3145 5399 3179
rect 5917 3145 5951 3179
rect 7205 3145 7239 3179
rect 8125 3145 8159 3179
rect 9597 3145 9631 3179
rect 9689 3145 9723 3179
rect 11897 3145 11931 3179
rect 13553 3145 13587 3179
rect 15761 3145 15795 3179
rect 16129 3145 16163 3179
rect 16957 3145 16991 3179
rect 18199 3145 18233 3179
rect 7435 3077 7469 3111
rect 8401 3009 8435 3043
rect 9045 3009 9079 3043
rect 1444 2941 1478 2975
rect 1869 2941 1903 2975
rect 2513 2941 2547 2975
rect 3433 2941 3467 2975
rect 5708 2941 5742 2975
rect 7364 2941 7398 2975
rect 9321 2941 9355 2975
rect 3157 2873 3191 2907
rect 4077 2873 4111 2907
rect 4169 2873 4203 2907
rect 4721 2873 4755 2907
rect 8493 2873 8527 2907
rect 10885 3077 10919 3111
rect 15209 3077 15243 3111
rect 10241 3009 10275 3043
rect 11253 3009 11287 3043
rect 16313 3009 16347 3043
rect 12265 2941 12299 2975
rect 12541 2941 12575 2975
rect 14197 2941 14231 2975
rect 15336 2941 15370 2975
rect 18128 2941 18162 2975
rect 9965 2873 9999 2907
rect 10057 2873 10091 2907
rect 12449 2873 12483 2907
rect 14841 2873 14875 2907
rect 15439 2873 15473 2907
rect 2237 2805 2271 2839
rect 3893 2805 3927 2839
rect 6193 2805 6227 2839
rect 7849 2805 7883 2839
rect 9597 2805 9631 2839
rect 14381 2805 14415 2839
rect 18613 2805 18647 2839
rect 3525 2601 3559 2635
rect 5365 2601 5399 2635
rect 5825 2601 5859 2635
rect 6561 2601 6595 2635
rect 8401 2601 8435 2635
rect 11989 2601 12023 2635
rect 3801 2533 3835 2567
rect 4445 2533 4479 2567
rect 4997 2533 5031 2567
rect 6285 2533 6319 2567
rect 7021 2533 7055 2567
rect 7113 2533 7147 2567
rect 10333 2533 10367 2567
rect 10609 2533 10643 2567
rect 11161 2533 11195 2567
rect 16037 2533 16071 2567
rect 2329 2465 2363 2499
rect 2881 2465 2915 2499
rect 6561 2465 6595 2499
rect 6653 2465 6687 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 13737 2465 13771 2499
rect 14289 2465 14323 2499
rect 15485 2465 15519 2499
rect 17268 2465 17302 2499
rect 17371 2465 17405 2499
rect 18613 2465 18647 2499
rect 19165 2465 19199 2499
rect 19993 2465 20027 2499
rect 20545 2465 20579 2499
rect 2697 2397 2731 2431
rect 4353 2397 4387 2431
rect 5641 2397 5675 2431
rect 7665 2397 7699 2431
rect 8677 2397 8711 2431
rect 9505 2397 9539 2431
rect 10517 2397 10551 2431
rect 17693 2397 17727 2431
rect 13921 2329 13955 2363
rect 1777 2261 1811 2295
rect 2145 2261 2179 2295
rect 12817 2261 12851 2295
rect 15669 2261 15703 2295
rect 18797 2261 18831 2295
rect 20177 2261 20211 2295
<< metal1 >>
rect 14 23536 20 23588
rect 72 23576 78 23588
rect 842 23576 848 23588
rect 72 23548 848 23576
rect 72 23536 78 23548
rect 842 23536 848 23548
rect 900 23536 906 23588
rect 1104 21786 22816 21808
rect 1104 21734 4982 21786
rect 5034 21734 5046 21786
rect 5098 21734 5110 21786
rect 5162 21734 5174 21786
rect 5226 21734 12982 21786
rect 13034 21734 13046 21786
rect 13098 21734 13110 21786
rect 13162 21734 13174 21786
rect 13226 21734 20982 21786
rect 21034 21734 21046 21786
rect 21098 21734 21110 21786
rect 21162 21734 21174 21786
rect 21226 21734 22816 21786
rect 1104 21712 22816 21734
rect 1104 21242 22816 21264
rect 1104 21190 8982 21242
rect 9034 21190 9046 21242
rect 9098 21190 9110 21242
rect 9162 21190 9174 21242
rect 9226 21190 16982 21242
rect 17034 21190 17046 21242
rect 17098 21190 17110 21242
rect 17162 21190 17174 21242
rect 17226 21190 22816 21242
rect 1104 21168 22816 21190
rect 106 20952 112 21004
rect 164 20992 170 21004
rect 9950 20992 9956 21004
rect 10008 21001 10014 21004
rect 10008 20995 10046 21001
rect 164 20964 9956 20992
rect 164 20952 170 20964
rect 9950 20952 9956 20964
rect 10034 20961 10046 20995
rect 10008 20955 10046 20961
rect 10008 20952 10014 20955
rect 10091 20791 10149 20797
rect 10091 20757 10103 20791
rect 10137 20788 10149 20791
rect 10226 20788 10232 20800
rect 10137 20760 10232 20788
rect 10137 20757 10149 20760
rect 10091 20751 10149 20757
rect 10226 20748 10232 20760
rect 10284 20748 10290 20800
rect 1104 20698 22816 20720
rect 1104 20646 4982 20698
rect 5034 20646 5046 20698
rect 5098 20646 5110 20698
rect 5162 20646 5174 20698
rect 5226 20646 12982 20698
rect 13034 20646 13046 20698
rect 13098 20646 13110 20698
rect 13162 20646 13174 20698
rect 13226 20646 20982 20698
rect 21034 20646 21046 20698
rect 21098 20646 21110 20698
rect 21162 20646 21174 20698
rect 21226 20646 22816 20698
rect 1104 20624 22816 20646
rect 4522 20584 4528 20596
rect 4483 20556 4528 20584
rect 4522 20544 4528 20556
rect 4580 20544 4586 20596
rect 6086 20584 6092 20596
rect 6047 20556 6092 20584
rect 6086 20544 6092 20556
rect 6144 20544 6150 20596
rect 7374 20584 7380 20596
rect 7335 20556 7380 20584
rect 7374 20544 7380 20556
rect 7432 20544 7438 20596
rect 8941 20587 8999 20593
rect 8941 20553 8953 20587
rect 8987 20584 8999 20587
rect 9306 20584 9312 20596
rect 8987 20556 9312 20584
rect 8987 20553 8999 20556
rect 8941 20547 8999 20553
rect 9306 20544 9312 20556
rect 9364 20544 9370 20596
rect 9950 20584 9956 20596
rect 9911 20556 9956 20584
rect 9950 20544 9956 20556
rect 10008 20544 10014 20596
rect 10962 20584 10968 20596
rect 10923 20556 10968 20584
rect 10962 20544 10968 20556
rect 11020 20544 11026 20596
rect 14001 20587 14059 20593
rect 14001 20584 14013 20587
rect 13786 20556 14013 20584
rect 1210 20340 1216 20392
rect 1268 20380 1274 20392
rect 1432 20383 1490 20389
rect 1432 20380 1444 20383
rect 1268 20352 1444 20380
rect 1268 20340 1274 20352
rect 1432 20349 1444 20352
rect 1478 20380 1490 20383
rect 1857 20383 1915 20389
rect 1857 20380 1869 20383
rect 1478 20352 1869 20380
rect 1478 20349 1490 20352
rect 1432 20343 1490 20349
rect 1857 20349 1869 20352
rect 1903 20349 1915 20383
rect 1857 20343 1915 20349
rect 4132 20383 4190 20389
rect 4132 20349 4144 20383
rect 4178 20380 4190 20383
rect 4522 20380 4528 20392
rect 4178 20352 4528 20380
rect 4178 20349 4190 20352
rect 4132 20343 4190 20349
rect 4522 20340 4528 20352
rect 4580 20340 4586 20392
rect 5696 20383 5754 20389
rect 5696 20349 5708 20383
rect 5742 20380 5754 20383
rect 6086 20380 6092 20392
rect 5742 20352 6092 20380
rect 5742 20349 5754 20352
rect 5696 20343 5754 20349
rect 6086 20340 6092 20352
rect 6144 20340 6150 20392
rect 6892 20383 6950 20389
rect 6892 20349 6904 20383
rect 6938 20380 6950 20383
rect 7374 20380 7380 20392
rect 6938 20352 7380 20380
rect 6938 20349 6950 20352
rect 6892 20343 6950 20349
rect 7374 20340 7380 20352
rect 7432 20340 7438 20392
rect 8757 20383 8815 20389
rect 8757 20349 8769 20383
rect 8803 20380 8815 20383
rect 10480 20383 10538 20389
rect 8803 20352 9444 20380
rect 8803 20349 8815 20352
rect 8757 20343 8815 20349
rect 9416 20256 9444 20352
rect 10480 20349 10492 20383
rect 10526 20380 10538 20383
rect 10962 20380 10968 20392
rect 10526 20352 10968 20380
rect 10526 20349 10538 20352
rect 10480 20343 10538 20349
rect 10962 20340 10968 20352
rect 11020 20340 11026 20392
rect 13516 20383 13574 20389
rect 13516 20349 13528 20383
rect 13562 20380 13574 20383
rect 13786 20380 13814 20556
rect 14001 20553 14013 20556
rect 14047 20584 14059 20587
rect 14274 20584 14280 20596
rect 14047 20556 14280 20584
rect 14047 20553 14059 20556
rect 14001 20547 14059 20553
rect 14274 20544 14280 20556
rect 14332 20544 14338 20596
rect 14737 20587 14795 20593
rect 14737 20553 14749 20587
rect 14783 20584 14795 20587
rect 15838 20584 15844 20596
rect 14783 20556 15844 20584
rect 14783 20553 14795 20556
rect 14737 20547 14795 20553
rect 15838 20544 15844 20556
rect 15896 20544 15902 20596
rect 16945 20587 17003 20593
rect 16945 20553 16957 20587
rect 16991 20584 17003 20587
rect 17678 20584 17684 20596
rect 16991 20556 17684 20584
rect 16991 20553 17003 20556
rect 16945 20547 17003 20553
rect 14550 20380 14556 20392
rect 13562 20352 13814 20380
rect 14511 20352 14556 20380
rect 13562 20349 13574 20352
rect 13516 20343 13574 20349
rect 14550 20340 14556 20352
rect 14608 20380 14614 20392
rect 15105 20383 15163 20389
rect 15105 20380 15117 20383
rect 14608 20352 15117 20380
rect 14608 20340 14614 20352
rect 15105 20349 15117 20352
rect 15151 20349 15163 20383
rect 15105 20343 15163 20349
rect 16460 20383 16518 20389
rect 16460 20349 16472 20383
rect 16506 20380 16518 20383
rect 16960 20380 16988 20547
rect 17678 20544 17684 20556
rect 17736 20544 17742 20596
rect 18601 20587 18659 20593
rect 18601 20553 18613 20587
rect 18647 20584 18659 20587
rect 21266 20584 21272 20596
rect 18647 20556 21272 20584
rect 18647 20553 18659 20556
rect 18601 20547 18659 20553
rect 16506 20352 16988 20380
rect 18116 20383 18174 20389
rect 16506 20349 16518 20352
rect 16460 20343 16518 20349
rect 18116 20349 18128 20383
rect 18162 20380 18174 20383
rect 18616 20380 18644 20547
rect 21266 20544 21272 20556
rect 21324 20544 21330 20596
rect 21450 20584 21456 20596
rect 21411 20556 21456 20584
rect 21450 20544 21456 20556
rect 21508 20544 21514 20596
rect 18162 20352 18644 20380
rect 20968 20383 21026 20389
rect 18162 20349 18174 20352
rect 18116 20343 18174 20349
rect 20968 20349 20980 20383
rect 21014 20380 21026 20383
rect 21450 20380 21456 20392
rect 21014 20352 21456 20380
rect 21014 20349 21026 20352
rect 20968 20343 21026 20349
rect 21450 20340 21456 20352
rect 21508 20340 21514 20392
rect 1535 20247 1593 20253
rect 1535 20213 1547 20247
rect 1581 20244 1593 20247
rect 1946 20244 1952 20256
rect 1581 20216 1952 20244
rect 1581 20213 1593 20216
rect 1535 20207 1593 20213
rect 1946 20204 1952 20216
rect 2004 20204 2010 20256
rect 3786 20204 3792 20256
rect 3844 20244 3850 20256
rect 4203 20247 4261 20253
rect 4203 20244 4215 20247
rect 3844 20216 4215 20244
rect 3844 20204 3850 20216
rect 4203 20213 4215 20216
rect 4249 20213 4261 20247
rect 4203 20207 4261 20213
rect 5767 20247 5825 20253
rect 5767 20213 5779 20247
rect 5813 20244 5825 20247
rect 6270 20244 6276 20256
rect 5813 20216 6276 20244
rect 5813 20213 5825 20216
rect 5767 20207 5825 20213
rect 6270 20204 6276 20216
rect 6328 20204 6334 20256
rect 6638 20204 6644 20256
rect 6696 20244 6702 20256
rect 6963 20247 7021 20253
rect 6963 20244 6975 20247
rect 6696 20216 6975 20244
rect 6696 20204 6702 20216
rect 6963 20213 6975 20216
rect 7009 20213 7021 20247
rect 9398 20244 9404 20256
rect 9359 20216 9404 20244
rect 6963 20207 7021 20213
rect 9398 20204 9404 20216
rect 9456 20204 9462 20256
rect 10551 20247 10609 20253
rect 10551 20213 10563 20247
rect 10597 20244 10609 20247
rect 12526 20244 12532 20256
rect 10597 20216 12532 20244
rect 10597 20213 10609 20216
rect 10551 20207 10609 20213
rect 12526 20204 12532 20216
rect 12584 20204 12590 20256
rect 13354 20204 13360 20256
rect 13412 20244 13418 20256
rect 13587 20247 13645 20253
rect 13587 20244 13599 20247
rect 13412 20216 13599 20244
rect 13412 20204 13418 20216
rect 13587 20213 13599 20216
rect 13633 20213 13645 20247
rect 13587 20207 13645 20213
rect 14918 20204 14924 20256
rect 14976 20244 14982 20256
rect 16531 20247 16589 20253
rect 16531 20244 16543 20247
rect 14976 20216 16543 20244
rect 14976 20204 14982 20216
rect 16531 20213 16543 20216
rect 16577 20213 16589 20247
rect 16531 20207 16589 20213
rect 17494 20204 17500 20256
rect 17552 20244 17558 20256
rect 18187 20247 18245 20253
rect 18187 20244 18199 20247
rect 17552 20216 18199 20244
rect 17552 20204 17558 20216
rect 18187 20213 18199 20216
rect 18233 20213 18245 20247
rect 18187 20207 18245 20213
rect 20622 20204 20628 20256
rect 20680 20244 20686 20256
rect 21039 20247 21097 20253
rect 21039 20244 21051 20247
rect 20680 20216 21051 20244
rect 20680 20204 20686 20216
rect 21039 20213 21051 20216
rect 21085 20213 21097 20247
rect 21039 20207 21097 20213
rect 1104 20154 22816 20176
rect 1104 20102 8982 20154
rect 9034 20102 9046 20154
rect 9098 20102 9110 20154
rect 9162 20102 9174 20154
rect 9226 20102 16982 20154
rect 17034 20102 17046 20154
rect 17098 20102 17110 20154
rect 17162 20102 17174 20154
rect 17226 20102 22816 20154
rect 1104 20080 22816 20102
rect 1578 20040 1584 20052
rect 1539 20012 1584 20040
rect 1578 20000 1584 20012
rect 1636 20000 1642 20052
rect 9398 20000 9404 20052
rect 9456 20040 9462 20052
rect 9815 20043 9873 20049
rect 9815 20040 9827 20043
rect 9456 20012 9827 20040
rect 9456 20000 9462 20012
rect 9815 20009 9827 20012
rect 9861 20009 9873 20043
rect 9815 20003 9873 20009
rect 10226 19932 10232 19984
rect 10284 19972 10290 19984
rect 10965 19975 11023 19981
rect 10965 19972 10977 19975
rect 10284 19944 10977 19972
rect 10284 19932 10290 19944
rect 10965 19941 10977 19944
rect 11011 19941 11023 19975
rect 10965 19935 11023 19941
rect 11057 19975 11115 19981
rect 11057 19941 11069 19975
rect 11103 19972 11115 19975
rect 11330 19972 11336 19984
rect 11103 19944 11336 19972
rect 11103 19941 11115 19944
rect 11057 19935 11115 19941
rect 11330 19932 11336 19944
rect 11388 19932 11394 19984
rect 12618 19972 12624 19984
rect 12579 19944 12624 19972
rect 12618 19932 12624 19944
rect 12676 19932 12682 19984
rect 1302 19864 1308 19916
rect 1360 19904 1366 19916
rect 1397 19907 1455 19913
rect 1397 19904 1409 19907
rect 1360 19876 1409 19904
rect 1360 19864 1366 19876
rect 1397 19873 1409 19876
rect 1443 19873 1455 19907
rect 1397 19867 1455 19873
rect 2568 19907 2626 19913
rect 2568 19873 2580 19907
rect 2614 19904 2626 19907
rect 2774 19904 2780 19916
rect 2614 19876 2780 19904
rect 2614 19873 2626 19876
rect 2568 19867 2626 19873
rect 2774 19864 2780 19876
rect 2832 19864 2838 19916
rect 5626 19864 5632 19916
rect 5684 19904 5690 19916
rect 6089 19907 6147 19913
rect 6089 19904 6101 19907
rect 5684 19876 6101 19904
rect 5684 19864 5690 19876
rect 6089 19873 6101 19876
rect 6135 19873 6147 19907
rect 6089 19867 6147 19873
rect 9744 19907 9802 19913
rect 9744 19873 9756 19907
rect 9790 19904 9802 19907
rect 10042 19904 10048 19916
rect 9790 19876 10048 19904
rect 9790 19873 9802 19876
rect 9744 19867 9802 19873
rect 10042 19864 10048 19876
rect 10100 19864 10106 19916
rect 18024 19907 18082 19913
rect 18024 19873 18036 19907
rect 18070 19904 18082 19907
rect 18690 19904 18696 19916
rect 18070 19876 18696 19904
rect 18070 19873 18082 19876
rect 18024 19867 18082 19873
rect 18690 19864 18696 19876
rect 18748 19864 18754 19916
rect 12526 19836 12532 19848
rect 12487 19808 12532 19836
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 12710 19796 12716 19848
rect 12768 19836 12774 19848
rect 12805 19839 12863 19845
rect 12805 19836 12817 19839
rect 12768 19808 12817 19836
rect 12768 19796 12774 19808
rect 12805 19805 12817 19808
rect 12851 19805 12863 19839
rect 12805 19799 12863 19805
rect 11517 19771 11575 19777
rect 11517 19737 11529 19771
rect 11563 19768 11575 19771
rect 12728 19768 12756 19796
rect 11563 19740 12756 19768
rect 11563 19737 11575 19740
rect 11517 19731 11575 19737
rect 2639 19703 2697 19709
rect 2639 19669 2651 19703
rect 2685 19700 2697 19703
rect 3418 19700 3424 19712
rect 2685 19672 3424 19700
rect 2685 19669 2697 19672
rect 2639 19663 2697 19669
rect 3418 19660 3424 19672
rect 3476 19660 3482 19712
rect 6454 19700 6460 19712
rect 6415 19672 6460 19700
rect 6454 19660 6460 19672
rect 6512 19660 6518 19712
rect 10042 19660 10048 19712
rect 10100 19700 10106 19712
rect 10137 19703 10195 19709
rect 10137 19700 10149 19703
rect 10100 19672 10149 19700
rect 10100 19660 10106 19672
rect 10137 19669 10149 19672
rect 10183 19669 10195 19703
rect 10137 19663 10195 19669
rect 17862 19660 17868 19712
rect 17920 19700 17926 19712
rect 18095 19703 18153 19709
rect 18095 19700 18107 19703
rect 17920 19672 18107 19700
rect 17920 19660 17926 19672
rect 18095 19669 18107 19672
rect 18141 19669 18153 19703
rect 18095 19663 18153 19669
rect 1104 19610 22816 19632
rect 1104 19558 4982 19610
rect 5034 19558 5046 19610
rect 5098 19558 5110 19610
rect 5162 19558 5174 19610
rect 5226 19558 12982 19610
rect 13034 19558 13046 19610
rect 13098 19558 13110 19610
rect 13162 19558 13174 19610
rect 13226 19558 20982 19610
rect 21034 19558 21046 19610
rect 21098 19558 21110 19610
rect 21162 19558 21174 19610
rect 21226 19558 22816 19610
rect 1104 19536 22816 19558
rect 2774 19456 2780 19508
rect 2832 19496 2838 19508
rect 2961 19499 3019 19505
rect 2961 19496 2973 19499
rect 2832 19468 2973 19496
rect 2832 19456 2838 19468
rect 2961 19465 2973 19468
rect 3007 19465 3019 19499
rect 2961 19459 3019 19465
rect 6454 19456 6460 19508
rect 6512 19496 6518 19508
rect 6549 19499 6607 19505
rect 6549 19496 6561 19499
rect 6512 19468 6561 19496
rect 6512 19456 6518 19468
rect 6549 19465 6561 19468
rect 6595 19465 6607 19499
rect 10226 19496 10232 19508
rect 10187 19468 10232 19496
rect 6549 19459 6607 19465
rect 10226 19456 10232 19468
rect 10284 19456 10290 19508
rect 12253 19499 12311 19505
rect 12253 19465 12265 19499
rect 12299 19496 12311 19499
rect 12526 19496 12532 19508
rect 12299 19468 12532 19496
rect 12299 19465 12311 19468
rect 12253 19459 12311 19465
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 12802 19456 12808 19508
rect 12860 19496 12866 19508
rect 12897 19499 12955 19505
rect 12897 19496 12909 19499
rect 12860 19468 12909 19496
rect 12860 19456 12866 19468
rect 12897 19465 12909 19468
rect 12943 19465 12955 19499
rect 12897 19459 12955 19465
rect 19061 19499 19119 19505
rect 19061 19465 19073 19499
rect 19107 19496 19119 19499
rect 19426 19496 19432 19508
rect 19107 19468 19432 19496
rect 19107 19465 19119 19468
rect 19061 19459 19119 19465
rect 1578 19428 1584 19440
rect 1539 19400 1584 19428
rect 1578 19388 1584 19400
rect 1636 19388 1642 19440
rect 5261 19363 5319 19369
rect 5261 19360 5273 19363
rect 4775 19332 5273 19360
rect 4775 19301 4803 19332
rect 5261 19329 5273 19332
rect 5307 19360 5319 19363
rect 11517 19363 11575 19369
rect 5307 19332 7604 19360
rect 5307 19329 5319 19332
rect 5261 19323 5319 19329
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19261 1455 19295
rect 1397 19255 1455 19261
rect 4760 19295 4818 19301
rect 4760 19261 4772 19295
rect 4806 19261 4818 19295
rect 4760 19255 4818 19261
rect 1412 19224 1440 19255
rect 7576 19236 7604 19332
rect 11517 19329 11529 19363
rect 11563 19360 11575 19363
rect 12618 19360 12624 19372
rect 11563 19332 12624 19360
rect 11563 19329 11575 19332
rect 11517 19323 11575 19329
rect 12618 19320 12624 19332
rect 12676 19360 12682 19372
rect 13265 19363 13323 19369
rect 13265 19360 13277 19363
rect 12676 19332 13277 19360
rect 12676 19320 12682 19332
rect 13265 19329 13277 19332
rect 13311 19329 13323 19363
rect 13265 19323 13323 19329
rect 8941 19295 8999 19301
rect 8941 19261 8953 19295
rect 8987 19292 8999 19295
rect 9490 19292 9496 19304
rect 8987 19264 9496 19292
rect 8987 19261 8999 19264
rect 8941 19255 8999 19261
rect 9490 19252 9496 19264
rect 9548 19252 9554 19304
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19292 10747 19295
rect 11330 19292 11336 19304
rect 10735 19264 11336 19292
rect 10735 19261 10747 19264
rect 10689 19255 10747 19261
rect 11330 19252 11336 19264
rect 11388 19252 11394 19304
rect 12504 19295 12562 19301
rect 12504 19261 12516 19295
rect 12550 19292 12562 19295
rect 12802 19292 12808 19304
rect 12550 19264 12808 19292
rect 12550 19261 12562 19264
rect 12504 19255 12562 19261
rect 12802 19252 12808 19264
rect 12860 19252 12866 19304
rect 18208 19295 18266 19301
rect 18208 19261 18220 19295
rect 18254 19292 18266 19295
rect 19076 19292 19104 19459
rect 19426 19456 19432 19468
rect 19484 19456 19490 19508
rect 18254 19264 19104 19292
rect 18254 19261 18266 19264
rect 18208 19255 18266 19261
rect 2409 19227 2467 19233
rect 2409 19224 2421 19227
rect 1412 19196 2421 19224
rect 2409 19193 2421 19196
rect 2455 19224 2467 19227
rect 4847 19227 4905 19233
rect 4847 19224 4859 19227
rect 2455 19196 4859 19224
rect 2455 19193 2467 19196
rect 2409 19187 2467 19193
rect 4847 19193 4859 19196
rect 4893 19193 4905 19227
rect 4847 19187 4905 19193
rect 5721 19227 5779 19233
rect 5721 19193 5733 19227
rect 5767 19224 5779 19227
rect 6273 19227 6331 19233
rect 6273 19224 6285 19227
rect 5767 19196 6285 19224
rect 5767 19193 5779 19196
rect 5721 19187 5779 19193
rect 6273 19193 6285 19196
rect 6319 19224 6331 19227
rect 6917 19227 6975 19233
rect 6917 19224 6929 19227
rect 6319 19196 6929 19224
rect 6319 19193 6331 19196
rect 6273 19187 6331 19193
rect 6917 19193 6929 19196
rect 6963 19193 6975 19227
rect 6917 19187 6975 19193
rect 7009 19227 7067 19233
rect 7009 19193 7021 19227
rect 7055 19193 7067 19227
rect 7558 19224 7564 19236
rect 7519 19196 7564 19224
rect 7009 19187 7067 19193
rect 1302 19116 1308 19168
rect 1360 19156 1366 19168
rect 1949 19159 2007 19165
rect 1949 19156 1961 19159
rect 1360 19128 1961 19156
rect 1360 19116 1366 19128
rect 1949 19125 1961 19128
rect 1995 19125 2007 19159
rect 1949 19119 2007 19125
rect 2038 19116 2044 19168
rect 2096 19156 2102 19168
rect 2501 19159 2559 19165
rect 2501 19156 2513 19159
rect 2096 19128 2513 19156
rect 2096 19116 2102 19128
rect 2501 19125 2513 19128
rect 2547 19125 2559 19159
rect 5626 19156 5632 19168
rect 5587 19128 5632 19156
rect 2501 19119 2559 19125
rect 5626 19116 5632 19128
rect 5684 19116 5690 19168
rect 6454 19116 6460 19168
rect 6512 19156 6518 19168
rect 7024 19156 7052 19187
rect 7558 19184 7564 19196
rect 7616 19184 7622 19236
rect 9766 19224 9772 19236
rect 9727 19196 9772 19224
rect 9766 19184 9772 19196
rect 9824 19184 9830 19236
rect 18690 19224 18696 19236
rect 18603 19196 18696 19224
rect 18690 19184 18696 19196
rect 18748 19224 18754 19236
rect 22830 19224 22836 19236
rect 18748 19196 22836 19224
rect 18748 19184 18754 19196
rect 22830 19184 22836 19196
rect 22888 19184 22894 19236
rect 6512 19128 7052 19156
rect 6512 19116 6518 19128
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 12575 19159 12633 19165
rect 12575 19156 12587 19159
rect 12492 19128 12587 19156
rect 12492 19116 12498 19128
rect 12575 19125 12587 19128
rect 12621 19125 12633 19159
rect 12575 19119 12633 19125
rect 12802 19116 12808 19168
rect 12860 19156 12866 19168
rect 18279 19159 18337 19165
rect 18279 19156 18291 19159
rect 12860 19128 18291 19156
rect 12860 19116 12866 19128
rect 18279 19125 18291 19128
rect 18325 19125 18337 19159
rect 18279 19119 18337 19125
rect 1104 19066 22816 19088
rect 1104 19014 8982 19066
rect 9034 19014 9046 19066
rect 9098 19014 9110 19066
rect 9162 19014 9174 19066
rect 9226 19014 16982 19066
rect 17034 19014 17046 19066
rect 17098 19014 17110 19066
rect 17162 19014 17174 19066
rect 17226 19014 22816 19066
rect 1104 18992 22816 19014
rect 106 18912 112 18964
rect 164 18952 170 18964
rect 1581 18955 1639 18961
rect 1581 18952 1593 18955
rect 164 18924 1593 18952
rect 164 18912 170 18924
rect 1581 18921 1593 18924
rect 1627 18921 1639 18955
rect 2038 18952 2044 18964
rect 1999 18924 2044 18952
rect 1581 18915 1639 18921
rect 2038 18912 2044 18924
rect 2096 18912 2102 18964
rect 12434 18952 12440 18964
rect 12395 18924 12440 18952
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 6730 18884 6736 18896
rect 6691 18856 6736 18884
rect 6730 18844 6736 18856
rect 6788 18844 6794 18896
rect 9766 18844 9772 18896
rect 9824 18884 9830 18896
rect 9861 18887 9919 18893
rect 9861 18884 9873 18887
rect 9824 18856 9873 18884
rect 9824 18844 9830 18856
rect 9861 18853 9873 18856
rect 9907 18853 9919 18887
rect 12894 18884 12900 18896
rect 12855 18856 12900 18884
rect 9861 18847 9919 18853
rect 12894 18844 12900 18856
rect 12952 18844 12958 18896
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 2501 18819 2559 18825
rect 1443 18788 2452 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 2424 18689 2452 18788
rect 2501 18785 2513 18819
rect 2547 18816 2559 18819
rect 2590 18816 2596 18828
rect 2547 18788 2596 18816
rect 2547 18785 2559 18788
rect 2501 18779 2559 18785
rect 2590 18776 2596 18788
rect 2648 18776 2654 18828
rect 4338 18816 4344 18828
rect 4299 18788 4344 18816
rect 4338 18776 4344 18788
rect 4396 18776 4402 18828
rect 20968 18819 21026 18825
rect 20968 18785 20980 18819
rect 21014 18816 21026 18819
rect 21266 18816 21272 18828
rect 21014 18788 21272 18816
rect 21014 18785 21026 18788
rect 20968 18779 21026 18785
rect 21266 18776 21272 18788
rect 21324 18776 21330 18828
rect 3510 18708 3516 18760
rect 3568 18748 3574 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 3568 18720 4077 18748
rect 3568 18708 3574 18720
rect 4065 18717 4077 18720
rect 4111 18717 4123 18751
rect 6638 18748 6644 18760
rect 6599 18720 6644 18748
rect 4065 18711 4123 18717
rect 6638 18708 6644 18720
rect 6696 18708 6702 18760
rect 6914 18748 6920 18760
rect 6875 18720 6920 18748
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 8573 18751 8631 18757
rect 8573 18717 8585 18751
rect 8619 18748 8631 18751
rect 9122 18748 9128 18760
rect 8619 18720 9128 18748
rect 8619 18717 8631 18720
rect 8573 18711 8631 18717
rect 9122 18708 9128 18720
rect 9180 18748 9186 18760
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 9180 18720 9781 18748
rect 9180 18708 9186 18720
rect 9769 18717 9781 18720
rect 9815 18717 9827 18751
rect 10042 18748 10048 18760
rect 10003 18720 10048 18748
rect 9769 18711 9827 18717
rect 10042 18708 10048 18720
rect 10100 18708 10106 18760
rect 11882 18708 11888 18760
rect 11940 18748 11946 18760
rect 12802 18748 12808 18760
rect 11940 18720 12808 18748
rect 11940 18708 11946 18720
rect 12802 18708 12808 18720
rect 12860 18708 12866 18760
rect 13262 18748 13268 18760
rect 13223 18720 13268 18748
rect 13262 18708 13268 18720
rect 13320 18708 13326 18760
rect 2409 18683 2467 18689
rect 2409 18649 2421 18683
rect 2455 18680 2467 18683
rect 4798 18680 4804 18692
rect 2455 18652 4804 18680
rect 2455 18649 2467 18652
rect 2409 18643 2467 18649
rect 4798 18640 4804 18652
rect 4856 18640 4862 18692
rect 2639 18615 2697 18621
rect 2639 18581 2651 18615
rect 2685 18612 2697 18615
rect 8754 18612 8760 18624
rect 2685 18584 8760 18612
rect 2685 18581 2697 18584
rect 2639 18575 2697 18581
rect 8754 18572 8760 18584
rect 8812 18572 8818 18624
rect 9398 18612 9404 18624
rect 9359 18584 9404 18612
rect 9398 18572 9404 18584
rect 9456 18572 9462 18624
rect 10873 18615 10931 18621
rect 10873 18581 10885 18615
rect 10919 18612 10931 18615
rect 11330 18612 11336 18624
rect 10919 18584 11336 18612
rect 10919 18581 10931 18584
rect 10873 18575 10931 18581
rect 11330 18572 11336 18584
rect 11388 18572 11394 18624
rect 16390 18572 16396 18624
rect 16448 18612 16454 18624
rect 21039 18615 21097 18621
rect 21039 18612 21051 18615
rect 16448 18584 21051 18612
rect 16448 18572 16454 18584
rect 21039 18581 21051 18584
rect 21085 18581 21097 18615
rect 21039 18575 21097 18581
rect 1104 18522 22816 18544
rect 1104 18470 4982 18522
rect 5034 18470 5046 18522
rect 5098 18470 5110 18522
rect 5162 18470 5174 18522
rect 5226 18470 12982 18522
rect 13034 18470 13046 18522
rect 13098 18470 13110 18522
rect 13162 18470 13174 18522
rect 13226 18470 20982 18522
rect 21034 18470 21046 18522
rect 21098 18470 21110 18522
rect 21162 18470 21174 18522
rect 21226 18470 22816 18522
rect 1104 18448 22816 18470
rect 4338 18408 4344 18420
rect 4299 18380 4344 18408
rect 4338 18368 4344 18380
rect 4396 18368 4402 18420
rect 4798 18368 4804 18420
rect 4856 18408 4862 18420
rect 5031 18411 5089 18417
rect 5031 18408 5043 18411
rect 4856 18380 5043 18408
rect 4856 18368 4862 18380
rect 5031 18377 5043 18380
rect 5077 18377 5089 18411
rect 5031 18371 5089 18377
rect 6641 18411 6699 18417
rect 6641 18377 6653 18411
rect 6687 18408 6699 18411
rect 6730 18408 6736 18420
rect 6687 18380 6736 18408
rect 6687 18377 6699 18380
rect 6641 18371 6699 18377
rect 6730 18368 6736 18380
rect 6788 18368 6794 18420
rect 9122 18408 9128 18420
rect 9083 18380 9128 18408
rect 9122 18368 9128 18380
rect 9180 18368 9186 18420
rect 9766 18368 9772 18420
rect 9824 18408 9830 18420
rect 10321 18411 10379 18417
rect 10321 18408 10333 18411
rect 9824 18380 10333 18408
rect 9824 18368 9830 18380
rect 10321 18377 10333 18380
rect 10367 18377 10379 18411
rect 11882 18408 11888 18420
rect 11843 18380 11888 18408
rect 10321 18371 10379 18377
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 20993 18411 21051 18417
rect 20993 18377 21005 18411
rect 21039 18408 21051 18411
rect 21266 18408 21272 18420
rect 21039 18380 21272 18408
rect 21039 18377 21051 18380
rect 20993 18371 21051 18377
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 2498 18300 2504 18352
rect 2556 18340 2562 18352
rect 2556 18312 4154 18340
rect 2556 18300 2562 18312
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 2038 18272 2044 18284
rect 1811 18244 2044 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 3418 18272 3424 18284
rect 3379 18244 3424 18272
rect 3418 18232 3424 18244
rect 3476 18232 3482 18284
rect 4126 18204 4154 18312
rect 12434 18300 12440 18352
rect 12492 18340 12498 18352
rect 12492 18312 12572 18340
rect 12492 18300 12498 18312
rect 5905 18275 5963 18281
rect 5905 18241 5917 18275
rect 5951 18272 5963 18275
rect 6638 18272 6644 18284
rect 5951 18244 6644 18272
rect 5951 18241 5963 18244
rect 5905 18235 5963 18241
rect 6638 18232 6644 18244
rect 6696 18232 6702 18284
rect 6914 18272 6920 18284
rect 6875 18244 6920 18272
rect 6914 18232 6920 18244
rect 6972 18232 6978 18284
rect 7558 18272 7564 18284
rect 7519 18244 7564 18272
rect 7558 18232 7564 18244
rect 7616 18232 7622 18284
rect 9398 18272 9404 18284
rect 9359 18244 9404 18272
rect 9398 18232 9404 18244
rect 9456 18232 9462 18284
rect 10042 18272 10048 18284
rect 10003 18244 10048 18272
rect 10042 18232 10048 18244
rect 10100 18232 10106 18284
rect 12544 18281 12572 18312
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12529 18235 12587 18241
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18272 13231 18275
rect 13262 18272 13268 18284
rect 13219 18244 13268 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 13262 18232 13268 18244
rect 13320 18232 13326 18284
rect 4928 18207 4986 18213
rect 4928 18204 4940 18207
rect 4126 18176 4940 18204
rect 4928 18173 4940 18176
rect 4974 18204 4986 18207
rect 5353 18207 5411 18213
rect 5353 18204 5365 18207
rect 4974 18176 5365 18204
rect 4974 18173 4986 18176
rect 4928 18167 4986 18173
rect 5353 18173 5365 18176
rect 5399 18173 5411 18207
rect 5353 18167 5411 18173
rect 1857 18139 1915 18145
rect 1857 18105 1869 18139
rect 1903 18105 1915 18139
rect 1857 18099 1915 18105
rect 2409 18139 2467 18145
rect 2409 18105 2421 18139
rect 2455 18136 2467 18139
rect 2498 18136 2504 18148
rect 2455 18108 2504 18136
rect 2455 18105 2467 18108
rect 2409 18099 2467 18105
rect 1670 18028 1676 18080
rect 1728 18068 1734 18080
rect 1872 18068 1900 18099
rect 2498 18096 2504 18108
rect 2556 18096 2562 18148
rect 3510 18096 3516 18148
rect 3568 18136 3574 18148
rect 4062 18136 4068 18148
rect 3568 18108 3613 18136
rect 4023 18108 4068 18136
rect 3568 18096 3574 18108
rect 4062 18096 4068 18108
rect 4120 18096 4126 18148
rect 5626 18096 5632 18148
rect 5684 18136 5690 18148
rect 6273 18139 6331 18145
rect 6273 18136 6285 18139
rect 5684 18108 6285 18136
rect 5684 18096 5690 18108
rect 6273 18105 6285 18108
rect 6319 18136 6331 18139
rect 7006 18136 7012 18148
rect 6319 18108 7012 18136
rect 6319 18105 6331 18108
rect 6273 18099 6331 18105
rect 7006 18096 7012 18108
rect 7064 18096 7070 18148
rect 9490 18136 9496 18148
rect 9451 18108 9496 18136
rect 9490 18096 9496 18108
rect 9548 18096 9554 18148
rect 12621 18139 12679 18145
rect 12621 18105 12633 18139
rect 12667 18105 12679 18139
rect 12621 18099 12679 18105
rect 1728 18040 1900 18068
rect 1728 18028 1734 18040
rect 2130 18028 2136 18080
rect 2188 18068 2194 18080
rect 2590 18068 2596 18080
rect 2188 18040 2596 18068
rect 2188 18028 2194 18040
rect 2590 18028 2596 18040
rect 2648 18068 2654 18080
rect 2685 18071 2743 18077
rect 2685 18068 2697 18071
rect 2648 18040 2697 18068
rect 2648 18028 2654 18040
rect 2685 18037 2697 18040
rect 2731 18037 2743 18071
rect 2685 18031 2743 18037
rect 3237 18071 3295 18077
rect 3237 18037 3249 18071
rect 3283 18068 3295 18071
rect 3528 18068 3556 18096
rect 12250 18068 12256 18080
rect 3283 18040 3556 18068
rect 12211 18040 12256 18068
rect 3283 18037 3295 18040
rect 3237 18031 3295 18037
rect 12250 18028 12256 18040
rect 12308 18068 12314 18080
rect 12636 18068 12664 18099
rect 12308 18040 12664 18068
rect 12308 18028 12314 18040
rect 12894 18028 12900 18080
rect 12952 18068 12958 18080
rect 13449 18071 13507 18077
rect 13449 18068 13461 18071
rect 12952 18040 13461 18068
rect 12952 18028 12958 18040
rect 13449 18037 13461 18040
rect 13495 18037 13507 18071
rect 13449 18031 13507 18037
rect 1104 17978 22816 18000
rect 1104 17926 8982 17978
rect 9034 17926 9046 17978
rect 9098 17926 9110 17978
rect 9162 17926 9174 17978
rect 9226 17926 16982 17978
rect 17034 17926 17046 17978
rect 17098 17926 17110 17978
rect 17162 17926 17174 17978
rect 17226 17926 22816 17978
rect 1104 17904 22816 17926
rect 3418 17864 3424 17876
rect 3379 17836 3424 17864
rect 3418 17824 3424 17836
rect 3476 17824 3482 17876
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7285 17867 7343 17873
rect 7285 17864 7297 17867
rect 6972 17836 7297 17864
rect 6972 17824 6978 17836
rect 2314 17796 2320 17808
rect 2275 17768 2320 17796
rect 2314 17756 2320 17768
rect 2372 17756 2378 17808
rect 4249 17799 4307 17805
rect 4249 17765 4261 17799
rect 4295 17796 4307 17799
rect 4338 17796 4344 17808
rect 4295 17768 4344 17796
rect 4295 17765 4307 17768
rect 4249 17759 4307 17765
rect 4338 17756 4344 17768
rect 4396 17756 4402 17808
rect 6454 17796 6460 17808
rect 6415 17768 6460 17796
rect 6454 17756 6460 17768
rect 6512 17756 6518 17808
rect 7024 17805 7052 17836
rect 7285 17833 7297 17836
rect 7331 17833 7343 17867
rect 8754 17864 8760 17876
rect 8715 17836 8760 17864
rect 7285 17827 7343 17833
rect 8754 17824 8760 17836
rect 8812 17824 8818 17876
rect 7009 17799 7067 17805
rect 7009 17796 7021 17799
rect 6987 17768 7021 17796
rect 7009 17765 7021 17768
rect 7055 17765 7067 17799
rect 7009 17759 7067 17765
rect 9766 17756 9772 17808
rect 9824 17796 9830 17808
rect 9861 17799 9919 17805
rect 9861 17796 9873 17799
rect 9824 17768 9873 17796
rect 9824 17756 9830 17768
rect 9861 17765 9873 17768
rect 9907 17765 9919 17799
rect 12250 17796 12256 17808
rect 12211 17768 12256 17796
rect 9861 17759 9919 17765
rect 12250 17756 12256 17768
rect 12308 17756 12314 17808
rect 12894 17728 12900 17740
rect 12855 17700 12900 17728
rect 12894 17688 12900 17700
rect 12952 17688 12958 17740
rect 2225 17663 2283 17669
rect 2225 17629 2237 17663
rect 2271 17629 2283 17663
rect 2498 17660 2504 17672
rect 2459 17632 2504 17660
rect 2225 17623 2283 17629
rect 2240 17592 2268 17623
rect 2498 17620 2504 17632
rect 2556 17620 2562 17672
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17660 4215 17663
rect 4246 17660 4252 17672
rect 4203 17632 4252 17660
rect 4203 17629 4215 17632
rect 4157 17623 4215 17629
rect 4246 17620 4252 17632
rect 4304 17620 4310 17672
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17629 4491 17663
rect 4433 17623 4491 17629
rect 4062 17592 4068 17604
rect 2240 17564 4068 17592
rect 4062 17552 4068 17564
rect 4120 17592 4126 17604
rect 4448 17592 4476 17623
rect 5902 17620 5908 17672
rect 5960 17660 5966 17672
rect 6365 17663 6423 17669
rect 6365 17660 6377 17663
rect 5960 17632 6377 17660
rect 5960 17620 5966 17632
rect 6365 17629 6377 17632
rect 6411 17629 6423 17663
rect 6365 17623 6423 17629
rect 9769 17663 9827 17669
rect 9769 17629 9781 17663
rect 9815 17660 9827 17663
rect 9858 17660 9864 17672
rect 9815 17632 9864 17660
rect 9815 17629 9827 17632
rect 9769 17623 9827 17629
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17629 10103 17663
rect 10045 17623 10103 17629
rect 4120 17564 4476 17592
rect 4120 17552 4126 17564
rect 9398 17552 9404 17604
rect 9456 17592 9462 17604
rect 10060 17592 10088 17623
rect 13722 17620 13728 17672
rect 13780 17660 13786 17672
rect 13817 17663 13875 17669
rect 13817 17660 13829 17663
rect 13780 17632 13829 17660
rect 13780 17620 13786 17632
rect 13817 17629 13829 17632
rect 13863 17629 13875 17663
rect 13817 17623 13875 17629
rect 9456 17564 10088 17592
rect 9456 17552 9462 17564
rect 1670 17524 1676 17536
rect 1631 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 9309 17527 9367 17533
rect 9309 17493 9321 17527
rect 9355 17524 9367 17527
rect 9490 17524 9496 17536
rect 9355 17496 9496 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 9490 17484 9496 17496
rect 9548 17524 9554 17536
rect 11238 17524 11244 17536
rect 9548 17496 11244 17524
rect 9548 17484 9554 17496
rect 11238 17484 11244 17496
rect 11296 17484 11302 17536
rect 1104 17434 22816 17456
rect 1104 17382 4982 17434
rect 5034 17382 5046 17434
rect 5098 17382 5110 17434
rect 5162 17382 5174 17434
rect 5226 17382 12982 17434
rect 13034 17382 13046 17434
rect 13098 17382 13110 17434
rect 13162 17382 13174 17434
rect 13226 17382 20982 17434
rect 21034 17382 21046 17434
rect 21098 17382 21110 17434
rect 21162 17382 21174 17434
rect 21226 17382 22816 17434
rect 1104 17360 22816 17382
rect 3329 17323 3387 17329
rect 3329 17289 3341 17323
rect 3375 17320 3387 17323
rect 4338 17320 4344 17332
rect 3375 17292 4344 17320
rect 3375 17289 3387 17292
rect 3329 17283 3387 17289
rect 4338 17280 4344 17292
rect 4396 17320 4402 17332
rect 4709 17323 4767 17329
rect 4709 17320 4721 17323
rect 4396 17292 4721 17320
rect 4396 17280 4402 17292
rect 4709 17289 4721 17292
rect 4755 17289 4767 17323
rect 4709 17283 4767 17289
rect 12713 17323 12771 17329
rect 12713 17289 12725 17323
rect 12759 17320 12771 17323
rect 12802 17320 12808 17332
rect 12759 17292 12808 17320
rect 12759 17289 12771 17292
rect 12713 17283 12771 17289
rect 12802 17280 12808 17292
rect 12860 17280 12866 17332
rect 8754 17212 8760 17264
rect 8812 17252 8818 17264
rect 9398 17252 9404 17264
rect 8812 17224 8892 17252
rect 9359 17224 9404 17252
rect 8812 17212 8818 17224
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 3789 17187 3847 17193
rect 3789 17153 3801 17187
rect 3835 17184 3847 17187
rect 4154 17184 4160 17196
rect 3835 17156 4160 17184
rect 3835 17153 3847 17156
rect 3789 17147 3847 17153
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17184 6423 17187
rect 6454 17184 6460 17196
rect 6411 17156 6460 17184
rect 6411 17153 6423 17156
rect 6365 17147 6423 17153
rect 6454 17144 6460 17156
rect 6512 17184 6518 17196
rect 8864 17193 8892 17224
rect 9398 17212 9404 17224
rect 9456 17212 9462 17264
rect 6825 17187 6883 17193
rect 6825 17184 6837 17187
rect 6512 17156 6837 17184
rect 6512 17144 6518 17156
rect 6825 17153 6837 17156
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 8849 17187 8907 17193
rect 8849 17153 8861 17187
rect 8895 17153 8907 17187
rect 8849 17147 8907 17153
rect 9858 17144 9864 17196
rect 9916 17184 9922 17196
rect 10226 17184 10232 17196
rect 9916 17156 10232 17184
rect 9916 17144 9922 17156
rect 10226 17144 10232 17156
rect 10284 17144 10290 17196
rect 12253 17187 12311 17193
rect 12253 17153 12265 17187
rect 12299 17184 12311 17187
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 12299 17156 13001 17184
rect 12299 17153 12311 17156
rect 12253 17147 12311 17153
rect 12989 17153 13001 17156
rect 13035 17184 13047 17187
rect 13262 17184 13268 17196
rect 13035 17156 13268 17184
rect 13035 17153 13047 17156
rect 12989 17147 13047 17153
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17116 1826 17128
rect 2314 17116 2320 17128
rect 1820 17088 2320 17116
rect 1820 17076 1826 17088
rect 2314 17076 2320 17088
rect 2372 17116 2378 17128
rect 2685 17119 2743 17125
rect 2685 17116 2697 17119
rect 2372 17088 2697 17116
rect 2372 17076 2378 17088
rect 2685 17085 2697 17088
rect 2731 17085 2743 17119
rect 2685 17079 2743 17085
rect 6730 17076 6736 17128
rect 6788 17116 6794 17128
rect 6917 17119 6975 17125
rect 6917 17116 6929 17119
rect 6788 17088 6929 17116
rect 6788 17076 6794 17088
rect 6917 17085 6929 17088
rect 6963 17085 6975 17119
rect 10781 17119 10839 17125
rect 10781 17116 10793 17119
rect 6917 17079 6975 17085
rect 10612 17088 10793 17116
rect 4110 17051 4168 17057
rect 4110 17017 4122 17051
rect 4156 17017 4168 17051
rect 4110 17011 4168 17017
rect 8941 17051 8999 17057
rect 8941 17017 8953 17051
rect 8987 17048 8999 17051
rect 9306 17048 9312 17060
rect 8987 17020 9312 17048
rect 8987 17017 8999 17020
rect 8941 17011 8999 17017
rect 2038 16940 2044 16992
rect 2096 16980 2102 16992
rect 3605 16983 3663 16989
rect 3605 16980 3617 16983
rect 2096 16952 3617 16980
rect 2096 16940 2102 16952
rect 3605 16949 3617 16952
rect 3651 16980 3663 16983
rect 4125 16980 4153 17011
rect 3651 16952 4153 16980
rect 3651 16949 3663 16952
rect 3605 16943 3663 16949
rect 4246 16940 4252 16992
rect 4304 16980 4310 16992
rect 4985 16983 5043 16989
rect 4985 16980 4997 16983
rect 4304 16952 4997 16980
rect 4304 16940 4310 16952
rect 4985 16949 4997 16952
rect 5031 16949 5043 16983
rect 5902 16980 5908 16992
rect 5863 16952 5908 16980
rect 4985 16943 5043 16949
rect 5902 16940 5908 16952
rect 5960 16940 5966 16992
rect 8665 16983 8723 16989
rect 8665 16949 8677 16983
rect 8711 16980 8723 16983
rect 8956 16980 8984 17011
rect 9306 17008 9312 17020
rect 9364 17008 9370 17060
rect 9766 16980 9772 16992
rect 8711 16952 8984 16980
rect 9727 16952 9772 16980
rect 8711 16949 8723 16952
rect 8665 16943 8723 16949
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10612 16989 10640 17088
rect 10781 17085 10793 17088
rect 10827 17085 10839 17119
rect 10781 17079 10839 17085
rect 11241 17119 11299 17125
rect 11241 17085 11253 17119
rect 11287 17085 11299 17119
rect 14369 17119 14427 17125
rect 14369 17116 14381 17119
rect 11241 17079 11299 17085
rect 13786 17088 14381 17116
rect 10686 17008 10692 17060
rect 10744 17048 10750 17060
rect 11256 17048 11284 17079
rect 11514 17048 11520 17060
rect 10744 17020 11284 17048
rect 11475 17020 11520 17048
rect 10744 17008 10750 17020
rect 11514 17008 11520 17020
rect 11572 17008 11578 17060
rect 13081 17051 13139 17057
rect 13081 17017 13093 17051
rect 13127 17017 13139 17051
rect 13630 17048 13636 17060
rect 13591 17020 13636 17048
rect 13081 17011 13139 17017
rect 10597 16983 10655 16989
rect 10597 16980 10609 16983
rect 10192 16952 10609 16980
rect 10192 16940 10198 16952
rect 10597 16949 10609 16952
rect 10643 16949 10655 16983
rect 10597 16943 10655 16949
rect 12986 16940 12992 16992
rect 13044 16980 13050 16992
rect 13096 16980 13124 17011
rect 13630 17008 13636 17020
rect 13688 17008 13694 17060
rect 13262 16980 13268 16992
rect 13044 16952 13268 16980
rect 13044 16940 13050 16952
rect 13262 16940 13268 16952
rect 13320 16980 13326 16992
rect 13786 16980 13814 17088
rect 14369 17085 14381 17088
rect 14415 17116 14427 17119
rect 14553 17119 14611 17125
rect 14553 17116 14565 17119
rect 14415 17088 14565 17116
rect 14415 17085 14427 17088
rect 14369 17079 14427 17085
rect 14553 17085 14565 17088
rect 14599 17085 14611 17119
rect 14553 17079 14611 17085
rect 14458 17048 14464 17060
rect 14419 17020 14464 17048
rect 14458 17008 14464 17020
rect 14516 17008 14522 17060
rect 13320 16952 13814 16980
rect 13320 16940 13326 16952
rect 1104 16890 22816 16912
rect 1104 16838 8982 16890
rect 9034 16838 9046 16890
rect 9098 16838 9110 16890
rect 9162 16838 9174 16890
rect 9226 16838 16982 16890
rect 17034 16838 17046 16890
rect 17098 16838 17110 16890
rect 17162 16838 17174 16890
rect 17226 16838 22816 16890
rect 1104 16816 22816 16838
rect 1762 16776 1768 16788
rect 1723 16748 1768 16776
rect 1762 16736 1768 16748
rect 1820 16776 1826 16788
rect 2777 16779 2835 16785
rect 2777 16776 2789 16779
rect 1820 16748 2789 16776
rect 1820 16736 1826 16748
rect 2777 16745 2789 16748
rect 2823 16745 2835 16779
rect 2777 16739 2835 16745
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 4157 16779 4215 16785
rect 4157 16776 4169 16779
rect 2924 16748 4169 16776
rect 2924 16736 2930 16748
rect 4157 16745 4169 16748
rect 4203 16745 4215 16779
rect 6362 16776 6368 16788
rect 6323 16748 6368 16776
rect 4157 16739 4215 16745
rect 6362 16736 6368 16748
rect 6420 16736 6426 16788
rect 6730 16736 6736 16788
rect 6788 16776 6794 16788
rect 6917 16779 6975 16785
rect 6917 16776 6929 16779
rect 6788 16748 6929 16776
rect 6788 16736 6794 16748
rect 6917 16745 6929 16748
rect 6963 16776 6975 16779
rect 7193 16779 7251 16785
rect 7193 16776 7205 16779
rect 6963 16748 7205 16776
rect 6963 16745 6975 16748
rect 6917 16739 6975 16745
rect 7193 16745 7205 16748
rect 7239 16745 7251 16779
rect 10134 16776 10140 16788
rect 7193 16739 7251 16745
rect 8312 16748 10140 16776
rect 2038 16668 2044 16720
rect 2096 16708 2102 16720
rect 2178 16711 2236 16717
rect 2178 16708 2190 16711
rect 2096 16680 2190 16708
rect 2096 16668 2102 16680
rect 2178 16677 2190 16680
rect 2224 16677 2236 16711
rect 2178 16671 2236 16677
rect 3145 16711 3203 16717
rect 3145 16677 3157 16711
rect 3191 16708 3203 16711
rect 4062 16708 4068 16720
rect 3191 16680 4068 16708
rect 3191 16677 3203 16680
rect 3145 16671 3203 16677
rect 4062 16668 4068 16680
rect 4120 16668 4126 16720
rect 3878 16600 3884 16652
rect 3936 16640 3942 16652
rect 4157 16643 4215 16649
rect 4157 16640 4169 16643
rect 3936 16612 4169 16640
rect 3936 16600 3942 16612
rect 4157 16609 4169 16612
rect 4203 16609 4215 16643
rect 4157 16603 4215 16609
rect 4617 16643 4675 16649
rect 4617 16609 4629 16643
rect 4663 16640 4675 16643
rect 4706 16640 4712 16652
rect 4663 16612 4712 16640
rect 4663 16609 4675 16612
rect 4617 16603 4675 16609
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 5442 16600 5448 16652
rect 5500 16640 5506 16652
rect 8110 16640 8116 16652
rect 5500 16612 8116 16640
rect 5500 16600 5506 16612
rect 8110 16600 8116 16612
rect 8168 16640 8174 16652
rect 8312 16649 8340 16748
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 11882 16776 11888 16788
rect 11843 16748 11888 16776
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12437 16779 12495 16785
rect 12437 16745 12449 16779
rect 12483 16776 12495 16779
rect 12802 16776 12808 16788
rect 12483 16748 12808 16776
rect 12483 16745 12495 16748
rect 12437 16739 12495 16745
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 12986 16776 12992 16788
rect 12947 16748 12992 16776
rect 12986 16736 12992 16748
rect 13044 16736 13050 16788
rect 9306 16668 9312 16720
rect 9364 16708 9370 16720
rect 9677 16711 9735 16717
rect 9677 16708 9689 16711
rect 9364 16680 9689 16708
rect 9364 16668 9370 16680
rect 9677 16677 9689 16680
rect 9723 16677 9735 16711
rect 13446 16708 13452 16720
rect 13407 16680 13452 16708
rect 9677 16671 9735 16677
rect 13446 16668 13452 16680
rect 13504 16708 13510 16720
rect 14458 16708 14464 16720
rect 13504 16680 14464 16708
rect 13504 16668 13510 16680
rect 14458 16668 14464 16680
rect 14516 16668 14522 16720
rect 8297 16643 8355 16649
rect 8297 16640 8309 16643
rect 8168 16612 8309 16640
rect 8168 16600 8174 16612
rect 8297 16609 8309 16612
rect 8343 16609 8355 16643
rect 8297 16603 8355 16609
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16640 8539 16643
rect 8662 16640 8668 16652
rect 8527 16612 8668 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 9490 16600 9496 16652
rect 9548 16640 9554 16652
rect 9766 16640 9772 16652
rect 9548 16612 9772 16640
rect 9548 16600 9554 16612
rect 9766 16600 9772 16612
rect 9824 16600 9830 16652
rect 15197 16643 15255 16649
rect 15197 16609 15209 16643
rect 15243 16640 15255 16643
rect 15378 16640 15384 16652
rect 15243 16612 15384 16640
rect 15243 16609 15255 16612
rect 15197 16603 15255 16609
rect 15378 16600 15384 16612
rect 15436 16600 15442 16652
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16572 1915 16575
rect 2866 16572 2872 16584
rect 1903 16544 2872 16572
rect 1903 16541 1915 16544
rect 1857 16535 1915 16541
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 5997 16575 6055 16581
rect 5997 16572 6009 16575
rect 5828 16544 6009 16572
rect 5828 16448 5856 16544
rect 5997 16541 6009 16544
rect 6043 16541 6055 16575
rect 8570 16572 8576 16584
rect 8531 16544 8576 16572
rect 5997 16535 6055 16541
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 11514 16572 11520 16584
rect 11475 16544 11520 16572
rect 11514 16532 11520 16544
rect 11572 16532 11578 16584
rect 13357 16575 13415 16581
rect 13357 16541 13369 16575
rect 13403 16541 13415 16575
rect 13630 16572 13636 16584
rect 13591 16544 13636 16572
rect 13357 16535 13415 16541
rect 13372 16504 13400 16535
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 13722 16504 13728 16516
rect 13372 16476 13728 16504
rect 13722 16464 13728 16476
rect 13780 16464 13786 16516
rect 3881 16439 3939 16445
rect 3881 16405 3893 16439
rect 3927 16436 3939 16439
rect 4154 16436 4160 16448
rect 3927 16408 4160 16436
rect 3927 16405 3939 16408
rect 3881 16399 3939 16405
rect 4154 16396 4160 16408
rect 4212 16396 4218 16448
rect 5810 16436 5816 16448
rect 5771 16408 5816 16436
rect 5810 16396 5816 16408
rect 5868 16396 5874 16448
rect 10686 16396 10692 16448
rect 10744 16436 10750 16448
rect 10781 16439 10839 16445
rect 10781 16436 10793 16439
rect 10744 16408 10793 16436
rect 10744 16396 10750 16408
rect 10781 16405 10793 16408
rect 10827 16405 10839 16439
rect 10781 16399 10839 16405
rect 14458 16396 14464 16448
rect 14516 16436 14522 16448
rect 15427 16439 15485 16445
rect 15427 16436 15439 16439
rect 14516 16408 15439 16436
rect 14516 16396 14522 16408
rect 15427 16405 15439 16408
rect 15473 16405 15485 16439
rect 15427 16399 15485 16405
rect 1104 16346 22816 16368
rect 1104 16294 4982 16346
rect 5034 16294 5046 16346
rect 5098 16294 5110 16346
rect 5162 16294 5174 16346
rect 5226 16294 12982 16346
rect 13034 16294 13046 16346
rect 13098 16294 13110 16346
rect 13162 16294 13174 16346
rect 13226 16294 20982 16346
rect 21034 16294 21046 16346
rect 21098 16294 21110 16346
rect 21162 16294 21174 16346
rect 21226 16294 22816 16346
rect 1104 16272 22816 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 2409 16235 2467 16241
rect 2409 16201 2421 16235
rect 2455 16232 2467 16235
rect 2866 16232 2872 16244
rect 2455 16204 2872 16232
rect 2455 16201 2467 16204
rect 2409 16195 2467 16201
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 8110 16232 8116 16244
rect 8071 16204 8116 16232
rect 8110 16192 8116 16204
rect 8168 16192 8174 16244
rect 11238 16232 11244 16244
rect 11199 16204 11244 16232
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 13446 16192 13452 16244
rect 13504 16232 13510 16244
rect 13633 16235 13691 16241
rect 13633 16232 13645 16235
rect 13504 16204 13645 16232
rect 13504 16192 13510 16204
rect 13633 16201 13645 16204
rect 13679 16201 13691 16235
rect 13633 16195 13691 16201
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 14001 16235 14059 16241
rect 14001 16232 14013 16235
rect 13780 16204 14013 16232
rect 13780 16192 13786 16204
rect 14001 16201 14013 16204
rect 14047 16201 14059 16235
rect 15378 16232 15384 16244
rect 15339 16204 15384 16232
rect 14001 16195 14059 16201
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 13262 16124 13268 16176
rect 13320 16164 13326 16176
rect 13357 16167 13415 16173
rect 13357 16164 13369 16167
rect 13320 16136 13369 16164
rect 13320 16124 13326 16136
rect 13357 16133 13369 16136
rect 13403 16133 13415 16167
rect 13357 16127 13415 16133
rect 5810 16096 5816 16108
rect 5771 16068 5816 16096
rect 5810 16056 5816 16068
rect 5868 16056 5874 16108
rect 6638 16056 6644 16108
rect 6696 16096 6702 16108
rect 8389 16099 8447 16105
rect 8389 16096 8401 16099
rect 6696 16068 8401 16096
rect 6696 16056 6702 16068
rect 8389 16065 8401 16068
rect 8435 16065 8447 16099
rect 8570 16096 8576 16108
rect 8531 16068 8576 16096
rect 8389 16059 8447 16065
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 15988 1458 16040
rect 2869 16031 2927 16037
rect 2869 15997 2881 16031
rect 2915 16028 2927 16031
rect 3602 16028 3608 16040
rect 2915 16000 3608 16028
rect 2915 15997 2927 16000
rect 2869 15991 2927 15997
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 4338 15988 4344 16040
rect 4396 16028 4402 16040
rect 5077 16031 5135 16037
rect 5077 16028 5089 16031
rect 4396 16000 5089 16028
rect 4396 15988 4402 16000
rect 5077 15997 5089 16000
rect 5123 16028 5135 16031
rect 5442 16028 5448 16040
rect 5123 16000 5448 16028
rect 5123 15997 5135 16000
rect 5077 15991 5135 15997
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 5721 16031 5779 16037
rect 5721 15997 5733 16031
rect 5767 15997 5779 16031
rect 5721 15991 5779 15997
rect 6457 16031 6515 16037
rect 6457 15997 6469 16031
rect 6503 16028 6515 16031
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6503 16000 6837 16028
rect 6503 15997 6515 16000
rect 6457 15991 6515 15997
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 7282 16028 7288 16040
rect 7243 16000 7288 16028
rect 6825 15991 6883 15997
rect 2958 15960 2964 15972
rect 2919 15932 2964 15960
rect 2958 15920 2964 15932
rect 3016 15920 3022 15972
rect 5258 15920 5264 15972
rect 5316 15960 5322 15972
rect 5736 15960 5764 15991
rect 7282 15988 7288 16000
rect 7340 15988 7346 16040
rect 7300 15960 7328 15988
rect 5316 15932 7328 15960
rect 8404 15960 8432 16059
rect 8570 16056 8576 16068
rect 8628 16056 8634 16108
rect 8662 15988 8668 16040
rect 8720 16028 8726 16040
rect 9769 16031 9827 16037
rect 9769 16028 9781 16031
rect 8720 16000 9781 16028
rect 8720 15988 8726 16000
rect 9769 15997 9781 16000
rect 9815 15997 9827 16031
rect 10318 16028 10324 16040
rect 10279 16000 10324 16028
rect 9769 15991 9827 15997
rect 10318 15988 10324 16000
rect 10376 15988 10382 16040
rect 12434 16028 12440 16040
rect 12395 16000 12440 16028
rect 12434 15988 12440 16000
rect 12492 15988 12498 16040
rect 13630 15988 13636 16040
rect 13688 16028 13694 16040
rect 14236 16031 14294 16037
rect 14236 16028 14248 16031
rect 13688 16000 14248 16028
rect 13688 15988 13694 16000
rect 14236 15997 14248 16000
rect 14282 16028 14294 16031
rect 14645 16031 14703 16037
rect 14645 16028 14657 16031
rect 14282 16000 14657 16028
rect 14282 15997 14294 16000
rect 14236 15991 14294 15997
rect 14645 15997 14657 16000
rect 14691 15997 14703 16031
rect 14645 15991 14703 15997
rect 8894 15963 8952 15969
rect 8894 15960 8906 15963
rect 8404 15932 8906 15960
rect 5316 15920 5322 15932
rect 8894 15929 8906 15932
rect 8940 15960 8952 15963
rect 10137 15963 10195 15969
rect 10137 15960 10149 15963
rect 8940 15932 10149 15960
rect 8940 15929 8952 15932
rect 8894 15923 8952 15929
rect 10137 15929 10149 15932
rect 10183 15960 10195 15963
rect 10226 15960 10232 15972
rect 10183 15932 10232 15960
rect 10183 15929 10195 15932
rect 10137 15923 10195 15929
rect 10226 15920 10232 15932
rect 10284 15960 10290 15972
rect 10642 15963 10700 15969
rect 10642 15960 10654 15963
rect 10284 15932 10654 15960
rect 10284 15920 10290 15932
rect 10642 15929 10654 15932
rect 10688 15960 10700 15963
rect 11517 15963 11575 15969
rect 11517 15960 11529 15963
rect 10688 15932 11529 15960
rect 10688 15929 10700 15932
rect 10642 15923 10700 15929
rect 11517 15929 11529 15932
rect 11563 15960 11575 15963
rect 11882 15960 11888 15972
rect 11563 15932 11888 15960
rect 11563 15929 11575 15932
rect 11517 15923 11575 15929
rect 11882 15920 11888 15932
rect 11940 15960 11946 15972
rect 12066 15960 12072 15972
rect 11940 15932 12072 15960
rect 11940 15920 11946 15932
rect 12066 15920 12072 15932
rect 12124 15960 12130 15972
rect 12161 15963 12219 15969
rect 12161 15960 12173 15963
rect 12124 15932 12173 15960
rect 12124 15920 12130 15932
rect 12161 15929 12173 15932
rect 12207 15960 12219 15963
rect 12758 15963 12816 15969
rect 12758 15960 12770 15963
rect 12207 15932 12770 15960
rect 12207 15929 12219 15932
rect 12161 15923 12219 15929
rect 12758 15929 12770 15932
rect 12804 15929 12816 15963
rect 14323 15963 14381 15969
rect 14323 15960 14335 15963
rect 12758 15923 12816 15929
rect 13786 15932 14335 15960
rect 2038 15892 2044 15904
rect 1999 15864 2044 15892
rect 2038 15852 2044 15864
rect 2096 15852 2102 15904
rect 3878 15852 3884 15904
rect 3936 15892 3942 15904
rect 4065 15895 4123 15901
rect 4065 15892 4077 15895
rect 3936 15864 4077 15892
rect 3936 15852 3942 15864
rect 4065 15861 4077 15864
rect 4111 15861 4123 15895
rect 4065 15855 4123 15861
rect 4525 15895 4583 15901
rect 4525 15861 4537 15895
rect 4571 15892 4583 15895
rect 4706 15892 4712 15904
rect 4571 15864 4712 15892
rect 4571 15861 4583 15864
rect 4525 15855 4583 15861
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 6273 15895 6331 15901
rect 6273 15861 6285 15895
rect 6319 15892 6331 15895
rect 6362 15892 6368 15904
rect 6319 15864 6368 15892
rect 6319 15861 6331 15864
rect 6273 15855 6331 15861
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 6454 15852 6460 15904
rect 6512 15892 6518 15904
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 6512 15864 6561 15892
rect 6512 15852 6518 15864
rect 6549 15861 6561 15864
rect 6595 15861 6607 15895
rect 6914 15892 6920 15904
rect 6875 15864 6920 15892
rect 6549 15855 6607 15861
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 9490 15892 9496 15904
rect 9451 15864 9496 15892
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 13630 15852 13636 15904
rect 13688 15892 13694 15904
rect 13786 15892 13814 15932
rect 14323 15929 14335 15932
rect 14369 15929 14381 15963
rect 14323 15923 14381 15929
rect 13688 15864 13814 15892
rect 13688 15852 13694 15864
rect 1104 15802 22816 15824
rect 1104 15750 8982 15802
rect 9034 15750 9046 15802
rect 9098 15750 9110 15802
rect 9162 15750 9174 15802
rect 9226 15750 16982 15802
rect 17034 15750 17046 15802
rect 17098 15750 17110 15802
rect 17162 15750 17174 15802
rect 17226 15750 22816 15802
rect 1104 15728 22816 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 5258 15688 5264 15700
rect 4212 15660 4257 15688
rect 5219 15660 5264 15688
rect 4212 15648 4218 15660
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 6825 15691 6883 15697
rect 6825 15657 6837 15691
rect 6871 15688 6883 15691
rect 7006 15688 7012 15700
rect 6871 15660 7012 15688
rect 6871 15657 6883 15660
rect 6825 15651 6883 15657
rect 7006 15648 7012 15660
rect 7064 15648 7070 15700
rect 8570 15648 8576 15700
rect 8628 15688 8634 15700
rect 9033 15691 9091 15697
rect 9033 15688 9045 15691
rect 8628 15660 9045 15688
rect 8628 15648 8634 15660
rect 9033 15657 9045 15660
rect 9079 15657 9091 15691
rect 9033 15651 9091 15657
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9548 15660 9873 15688
rect 9548 15648 9554 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 9861 15651 9919 15657
rect 11514 15648 11520 15700
rect 11572 15688 11578 15700
rect 11885 15691 11943 15697
rect 11885 15688 11897 15691
rect 11572 15660 11897 15688
rect 11572 15648 11578 15660
rect 11885 15657 11897 15660
rect 11931 15657 11943 15691
rect 11885 15651 11943 15657
rect 13354 15648 13360 15700
rect 13412 15688 13418 15700
rect 14274 15688 14280 15700
rect 13412 15660 14280 15688
rect 13412 15648 13418 15660
rect 14274 15648 14280 15660
rect 14332 15688 14338 15700
rect 14645 15691 14703 15697
rect 14645 15688 14657 15691
rect 14332 15660 14657 15688
rect 14332 15648 14338 15660
rect 14645 15657 14657 15660
rect 14691 15657 14703 15691
rect 14645 15651 14703 15657
rect 2409 15623 2467 15629
rect 2409 15589 2421 15623
rect 2455 15620 2467 15623
rect 2958 15620 2964 15632
rect 2455 15592 2964 15620
rect 2455 15589 2467 15592
rect 2409 15583 2467 15589
rect 2958 15580 2964 15592
rect 3016 15580 3022 15632
rect 6267 15623 6325 15629
rect 6267 15589 6279 15623
rect 6313 15620 6325 15623
rect 6362 15620 6368 15632
rect 6313 15592 6368 15620
rect 6313 15589 6325 15592
rect 6267 15583 6325 15589
rect 6362 15580 6368 15592
rect 6420 15580 6426 15632
rect 8757 15623 8815 15629
rect 8757 15589 8769 15623
rect 8803 15620 8815 15623
rect 10318 15620 10324 15632
rect 8803 15592 10324 15620
rect 8803 15589 8815 15592
rect 8757 15583 8815 15589
rect 10318 15580 10324 15592
rect 10376 15580 10382 15632
rect 11609 15623 11667 15629
rect 11609 15589 11621 15623
rect 11655 15620 11667 15623
rect 12434 15620 12440 15632
rect 11655 15592 12440 15620
rect 11655 15589 11667 15592
rect 11609 15583 11667 15589
rect 12434 15580 12440 15592
rect 12492 15620 12498 15632
rect 12805 15623 12863 15629
rect 12805 15620 12817 15623
rect 12492 15592 12817 15620
rect 12492 15580 12498 15592
rect 12805 15589 12817 15592
rect 12851 15589 12863 15623
rect 12805 15583 12863 15589
rect 13722 15580 13728 15632
rect 13780 15620 13786 15632
rect 13817 15623 13875 15629
rect 13817 15620 13829 15623
rect 13780 15592 13829 15620
rect 13780 15580 13786 15592
rect 13817 15589 13829 15592
rect 13863 15589 13875 15623
rect 13817 15583 13875 15589
rect 4338 15552 4344 15564
rect 4299 15524 4344 15552
rect 4338 15512 4344 15524
rect 4396 15512 4402 15564
rect 4525 15555 4583 15561
rect 4525 15521 4537 15555
rect 4571 15552 4583 15555
rect 4706 15552 4712 15564
rect 4571 15524 4712 15552
rect 4571 15521 4583 15524
rect 4525 15515 4583 15521
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 5442 15512 5448 15564
rect 5500 15552 5506 15564
rect 5905 15555 5963 15561
rect 5905 15552 5917 15555
rect 5500 15524 5917 15552
rect 5500 15512 5506 15524
rect 5905 15521 5917 15524
rect 5951 15552 5963 15555
rect 6914 15552 6920 15564
rect 5951 15524 6920 15552
rect 5951 15521 5963 15524
rect 5905 15515 5963 15521
rect 6914 15512 6920 15524
rect 6972 15512 6978 15564
rect 8018 15552 8024 15564
rect 7979 15524 8024 15552
rect 8018 15512 8024 15524
rect 8076 15512 8082 15564
rect 8573 15555 8631 15561
rect 8573 15521 8585 15555
rect 8619 15552 8631 15555
rect 8662 15552 8668 15564
rect 8619 15524 8668 15552
rect 8619 15521 8631 15524
rect 8573 15515 8631 15521
rect 8662 15512 8668 15524
rect 8720 15512 8726 15564
rect 10870 15552 10876 15564
rect 10831 15524 10876 15552
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 11333 15555 11391 15561
rect 11333 15521 11345 15555
rect 11379 15521 11391 15555
rect 11333 15515 11391 15521
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15484 2375 15487
rect 2682 15484 2688 15496
rect 2363 15456 2688 15484
rect 2363 15453 2375 15456
rect 2317 15447 2375 15453
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 3234 15484 3240 15496
rect 3007 15456 3240 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 3234 15444 3240 15456
rect 3292 15484 3298 15496
rect 4614 15484 4620 15496
rect 3292 15456 4620 15484
rect 3292 15444 3298 15456
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 11348 15484 11376 15515
rect 10704 15456 11376 15484
rect 13725 15487 13783 15493
rect 6730 15376 6736 15428
rect 6788 15416 6794 15428
rect 7101 15419 7159 15425
rect 7101 15416 7113 15419
rect 6788 15388 7113 15416
rect 6788 15376 6794 15388
rect 7101 15385 7113 15388
rect 7147 15416 7159 15419
rect 7282 15416 7288 15428
rect 7147 15388 7288 15416
rect 7147 15385 7159 15388
rect 7101 15379 7159 15385
rect 7282 15376 7288 15388
rect 7340 15376 7346 15428
rect 10704 15360 10732 15456
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 14458 15484 14464 15496
rect 13771 15456 14464 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 13446 15376 13452 15428
rect 13504 15416 13510 15428
rect 14277 15419 14335 15425
rect 14277 15416 14289 15419
rect 13504 15388 14289 15416
rect 13504 15376 13510 15388
rect 14277 15385 14289 15388
rect 14323 15385 14335 15419
rect 14277 15379 14335 15385
rect 1394 15308 1400 15360
rect 1452 15348 1458 15360
rect 1673 15351 1731 15357
rect 1673 15348 1685 15351
rect 1452 15320 1685 15348
rect 1452 15308 1458 15320
rect 1673 15317 1685 15320
rect 1719 15348 1731 15351
rect 3510 15348 3516 15360
rect 1719 15320 3516 15348
rect 1719 15317 1731 15320
rect 1673 15311 1731 15317
rect 3510 15308 3516 15320
rect 3568 15308 3574 15360
rect 10686 15348 10692 15360
rect 10647 15320 10692 15348
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 12342 15308 12348 15360
rect 12400 15348 12406 15360
rect 12437 15351 12495 15357
rect 12437 15348 12449 15351
rect 12400 15320 12449 15348
rect 12400 15308 12406 15320
rect 12437 15317 12449 15320
rect 12483 15317 12495 15351
rect 12437 15311 12495 15317
rect 1104 15258 22816 15280
rect 1104 15206 4982 15258
rect 5034 15206 5046 15258
rect 5098 15206 5110 15258
rect 5162 15206 5174 15258
rect 5226 15206 12982 15258
rect 13034 15206 13046 15258
rect 13098 15206 13110 15258
rect 13162 15206 13174 15258
rect 13226 15206 20982 15258
rect 21034 15206 21046 15258
rect 21098 15206 21110 15258
rect 21162 15206 21174 15258
rect 21226 15206 22816 15258
rect 1104 15184 22816 15206
rect 2869 15147 2927 15153
rect 2869 15113 2881 15147
rect 2915 15144 2927 15147
rect 2958 15144 2964 15156
rect 2915 15116 2964 15144
rect 2915 15113 2927 15116
rect 2869 15107 2927 15113
rect 2958 15104 2964 15116
rect 3016 15104 3022 15156
rect 3694 15104 3700 15156
rect 3752 15144 3758 15156
rect 3881 15147 3939 15153
rect 3881 15144 3893 15147
rect 3752 15116 3893 15144
rect 3752 15104 3758 15116
rect 3881 15113 3893 15116
rect 3927 15144 3939 15147
rect 4338 15144 4344 15156
rect 3927 15116 4344 15144
rect 3927 15113 3939 15116
rect 3881 15107 3939 15113
rect 4338 15104 4344 15116
rect 4396 15104 4402 15156
rect 4706 15144 4712 15156
rect 4448 15116 4712 15144
rect 3513 15079 3571 15085
rect 3513 15045 3525 15079
rect 3559 15076 3571 15079
rect 4448 15076 4476 15116
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 5442 15144 5448 15156
rect 5403 15116 5448 15144
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 10226 15144 10232 15156
rect 10187 15116 10232 15144
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 11330 15144 11336 15156
rect 11291 15116 11336 15144
rect 11330 15104 11336 15116
rect 11388 15104 11394 15156
rect 12066 15104 12072 15156
rect 12124 15144 12130 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 12124 15116 12173 15144
rect 12124 15104 12130 15116
rect 12161 15113 12173 15116
rect 12207 15113 12219 15147
rect 12161 15107 12219 15113
rect 13357 15147 13415 15153
rect 13357 15113 13369 15147
rect 13403 15144 13415 15147
rect 13722 15144 13728 15156
rect 13403 15116 13728 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 4614 15076 4620 15088
rect 3559 15048 4476 15076
rect 4575 15048 4620 15076
rect 3559 15045 3571 15048
rect 3513 15039 3571 15045
rect 4614 15036 4620 15048
rect 4672 15036 4678 15088
rect 13446 15036 13452 15088
rect 13504 15076 13510 15088
rect 13504 15048 14596 15076
rect 13504 15036 13510 15048
rect 1857 15011 1915 15017
rect 1857 14977 1869 15011
rect 1903 15008 1915 15011
rect 1946 15008 1952 15020
rect 1903 14980 1952 15008
rect 1903 14977 1915 14980
rect 1857 14971 1915 14977
rect 1946 14968 1952 14980
rect 2004 14968 2010 15020
rect 2314 15008 2320 15020
rect 2275 14980 2320 15008
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 4062 15008 4068 15020
rect 4023 14980 4068 15008
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 4246 14968 4252 15020
rect 4304 15008 4310 15020
rect 5675 15011 5733 15017
rect 5675 15008 5687 15011
rect 4304 14980 5687 15008
rect 4304 14968 4310 14980
rect 5675 14977 5687 14980
rect 5721 14977 5733 15011
rect 14274 15008 14280 15020
rect 14235 14980 14280 15008
rect 5675 14971 5733 14977
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 14568 15017 14596 15048
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 5588 14943 5646 14949
rect 5588 14909 5600 14943
rect 5634 14940 5646 14943
rect 5994 14940 6000 14952
rect 5634 14912 6000 14940
rect 5634 14909 5646 14912
rect 5588 14903 5646 14909
rect 5994 14900 6000 14912
rect 6052 14900 6058 14952
rect 9953 14943 10011 14949
rect 9953 14909 9965 14943
rect 9999 14940 10011 14943
rect 10318 14940 10324 14952
rect 9999 14912 10324 14940
rect 9999 14909 10011 14912
rect 9953 14903 10011 14909
rect 10318 14900 10324 14912
rect 10376 14940 10382 14952
rect 10413 14943 10471 14949
rect 10413 14940 10425 14943
rect 10376 14912 10425 14940
rect 10376 14900 10382 14912
rect 10413 14909 10425 14912
rect 10459 14909 10471 14943
rect 10413 14903 10471 14909
rect 12342 14900 12348 14952
rect 12400 14940 12406 14952
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 12400 14912 12449 14940
rect 12400 14900 12406 14912
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 18506 14900 18512 14952
rect 18564 14940 18570 14952
rect 18820 14943 18878 14949
rect 18820 14940 18832 14943
rect 18564 14912 18832 14940
rect 18564 14900 18570 14912
rect 18820 14909 18832 14912
rect 18866 14940 18878 14943
rect 19245 14943 19303 14949
rect 19245 14940 19257 14943
rect 18866 14912 19257 14940
rect 18866 14909 18878 14912
rect 18820 14903 18878 14909
rect 19245 14909 19257 14912
rect 19291 14909 19303 14943
rect 19245 14903 19303 14909
rect 1673 14875 1731 14881
rect 1673 14841 1685 14875
rect 1719 14872 1731 14875
rect 1949 14875 2007 14881
rect 1949 14872 1961 14875
rect 1719 14844 1961 14872
rect 1719 14841 1731 14844
rect 1673 14835 1731 14841
rect 1949 14841 1961 14844
rect 1995 14872 2007 14875
rect 2590 14872 2596 14884
rect 1995 14844 2596 14872
rect 1995 14841 2007 14844
rect 1949 14835 2007 14841
rect 2590 14832 2596 14844
rect 2648 14832 2654 14884
rect 3602 14832 3608 14884
rect 3660 14872 3666 14884
rect 4157 14875 4215 14881
rect 4157 14872 4169 14875
rect 3660 14844 4169 14872
rect 3660 14832 3666 14844
rect 4157 14841 4169 14844
rect 4203 14841 4215 14875
rect 4157 14835 4215 14841
rect 4172 14804 4200 14835
rect 10226 14832 10232 14884
rect 10284 14872 10290 14884
rect 10734 14875 10792 14881
rect 10734 14872 10746 14875
rect 10284 14844 10746 14872
rect 10284 14832 10290 14844
rect 10734 14841 10746 14844
rect 10780 14841 10792 14875
rect 10734 14835 10792 14841
rect 10870 14832 10876 14884
rect 10928 14872 10934 14884
rect 11609 14875 11667 14881
rect 11609 14872 11621 14875
rect 10928 14844 11621 14872
rect 10928 14832 10934 14844
rect 11609 14841 11621 14844
rect 11655 14841 11667 14875
rect 11609 14835 11667 14841
rect 12066 14832 12072 14884
rect 12124 14872 12130 14884
rect 12758 14875 12816 14881
rect 12758 14872 12770 14875
rect 12124 14844 12770 14872
rect 12124 14832 12130 14844
rect 12758 14841 12770 14844
rect 12804 14841 12816 14875
rect 12758 14835 12816 14841
rect 14369 14875 14427 14881
rect 14369 14841 14381 14875
rect 14415 14841 14427 14875
rect 14369 14835 14427 14841
rect 4982 14804 4988 14816
rect 4172 14776 4988 14804
rect 4982 14764 4988 14776
rect 5040 14764 5046 14816
rect 6362 14804 6368 14816
rect 6323 14776 6368 14804
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 6454 14764 6460 14816
rect 6512 14804 6518 14816
rect 8018 14804 8024 14816
rect 6512 14776 8024 14804
rect 6512 14764 6518 14776
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 8481 14807 8539 14813
rect 8481 14773 8493 14807
rect 8527 14804 8539 14807
rect 8662 14804 8668 14816
rect 8527 14776 8668 14804
rect 8527 14773 8539 14776
rect 8481 14767 8539 14773
rect 8662 14764 8668 14776
rect 8720 14764 8726 14816
rect 14090 14804 14096 14816
rect 14051 14776 14096 14804
rect 14090 14764 14096 14776
rect 14148 14804 14154 14816
rect 14384 14804 14412 14835
rect 14148 14776 14412 14804
rect 18923 14807 18981 14813
rect 14148 14764 14154 14776
rect 18923 14773 18935 14807
rect 18969 14804 18981 14807
rect 19702 14804 19708 14816
rect 18969 14776 19708 14804
rect 18969 14773 18981 14776
rect 18923 14767 18981 14773
rect 19702 14764 19708 14776
rect 19760 14764 19766 14816
rect 1104 14714 22816 14736
rect 1104 14662 8982 14714
rect 9034 14662 9046 14714
rect 9098 14662 9110 14714
rect 9162 14662 9174 14714
rect 9226 14662 16982 14714
rect 17034 14662 17046 14714
rect 17098 14662 17110 14714
rect 17162 14662 17174 14714
rect 17226 14662 22816 14714
rect 1104 14640 22816 14662
rect 2682 14600 2688 14612
rect 2643 14572 2688 14600
rect 2682 14560 2688 14572
rect 2740 14560 2746 14612
rect 3145 14603 3203 14609
rect 3145 14569 3157 14603
rect 3191 14600 3203 14603
rect 4246 14600 4252 14612
rect 3191 14572 4252 14600
rect 3191 14569 3203 14572
rect 3145 14563 3203 14569
rect 1854 14532 1860 14544
rect 1815 14504 1860 14532
rect 1854 14492 1860 14504
rect 1912 14492 1918 14544
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 3160 14396 3188 14563
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 4338 14560 4344 14612
rect 4396 14600 4402 14612
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 4396 14572 4445 14600
rect 4396 14560 4402 14572
rect 4433 14569 4445 14572
rect 4479 14569 4491 14603
rect 4982 14600 4988 14612
rect 4943 14572 4988 14600
rect 4433 14563 4491 14569
rect 4982 14560 4988 14572
rect 5040 14560 5046 14612
rect 10318 14600 10324 14612
rect 10279 14572 10324 14600
rect 10318 14560 10324 14572
rect 10376 14560 10382 14612
rect 14458 14600 14464 14612
rect 14419 14572 14464 14600
rect 14458 14560 14464 14572
rect 14516 14560 14522 14612
rect 19886 14600 19892 14612
rect 19847 14572 19892 14600
rect 19886 14560 19892 14572
rect 19944 14560 19950 14612
rect 3881 14535 3939 14541
rect 3881 14501 3893 14535
rect 3927 14532 3939 14535
rect 4062 14532 4068 14544
rect 3927 14504 4068 14532
rect 3927 14501 3939 14504
rect 3881 14495 3939 14501
rect 4062 14492 4068 14504
rect 4120 14492 4126 14544
rect 6267 14535 6325 14541
rect 6267 14501 6279 14535
rect 6313 14532 6325 14535
rect 6362 14532 6368 14544
rect 6313 14504 6368 14532
rect 6313 14501 6325 14504
rect 6267 14495 6325 14501
rect 6362 14492 6368 14504
rect 6420 14492 6426 14544
rect 12342 14532 12348 14544
rect 12303 14504 12348 14532
rect 12342 14492 12348 14504
rect 12400 14492 12406 14544
rect 14090 14532 14096 14544
rect 14051 14504 14096 14532
rect 14090 14492 14096 14504
rect 14148 14492 14154 14544
rect 16758 14532 16764 14544
rect 16719 14504 16764 14532
rect 16758 14492 16764 14504
rect 16816 14492 16822 14544
rect 10134 14464 10140 14476
rect 10095 14436 10140 14464
rect 10134 14424 10140 14436
rect 10192 14424 10198 14476
rect 10505 14467 10563 14473
rect 10505 14464 10517 14467
rect 10336 14436 10517 14464
rect 4062 14396 4068 14408
rect 1811 14368 3188 14396
rect 4023 14368 4068 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 5902 14396 5908 14408
rect 5863 14368 5908 14396
rect 5902 14356 5908 14368
rect 5960 14356 5966 14408
rect 8110 14356 8116 14408
rect 8168 14396 8174 14408
rect 8389 14399 8447 14405
rect 8389 14396 8401 14399
rect 8168 14368 8401 14396
rect 8168 14356 8174 14368
rect 8389 14365 8401 14368
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 9953 14399 10011 14405
rect 9953 14365 9965 14399
rect 9999 14396 10011 14399
rect 10226 14396 10232 14408
rect 9999 14368 10232 14396
rect 9999 14365 10011 14368
rect 9953 14359 10011 14365
rect 10226 14356 10232 14368
rect 10284 14396 10290 14408
rect 10336 14396 10364 14436
rect 10505 14433 10517 14436
rect 10551 14433 10563 14467
rect 11882 14464 11888 14476
rect 11843 14436 11888 14464
rect 10505 14427 10563 14433
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 12158 14464 12164 14476
rect 12119 14436 12164 14464
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 13722 14464 13728 14476
rect 13683 14436 13728 14464
rect 13722 14424 13728 14436
rect 13780 14424 13786 14476
rect 18782 14464 18788 14476
rect 18743 14436 18788 14464
rect 18782 14424 18788 14436
rect 18840 14424 18846 14476
rect 19702 14464 19708 14476
rect 19663 14436 19708 14464
rect 19702 14424 19708 14436
rect 19760 14424 19766 14476
rect 16666 14396 16672 14408
rect 10284 14368 10364 14396
rect 16627 14368 16672 14396
rect 10284 14356 10290 14368
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 17310 14396 17316 14408
rect 17271 14368 17316 14396
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 2314 14328 2320 14340
rect 2275 14300 2320 14328
rect 2314 14288 2320 14300
rect 2372 14288 2378 14340
rect 2590 14288 2596 14340
rect 2648 14328 2654 14340
rect 6825 14331 6883 14337
rect 6825 14328 6837 14331
rect 2648 14300 6837 14328
rect 2648 14288 2654 14300
rect 6825 14297 6837 14300
rect 6871 14297 6883 14331
rect 6825 14291 6883 14297
rect 10778 14288 10784 14340
rect 10836 14328 10842 14340
rect 11425 14331 11483 14337
rect 11425 14328 11437 14331
rect 10836 14300 11437 14328
rect 10836 14288 10842 14300
rect 11425 14297 11437 14300
rect 11471 14297 11483 14331
rect 11425 14291 11483 14297
rect 11054 14260 11060 14272
rect 11015 14232 11060 14260
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 12802 14260 12808 14272
rect 12763 14232 12808 14260
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 15470 14260 15476 14272
rect 15431 14232 15476 14260
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 18414 14260 18420 14272
rect 18375 14232 18420 14260
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 1104 14170 22816 14192
rect 1104 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 12982 14170
rect 13034 14118 13046 14170
rect 13098 14118 13110 14170
rect 13162 14118 13174 14170
rect 13226 14118 20982 14170
rect 21034 14118 21046 14170
rect 21098 14118 21110 14170
rect 21162 14118 21174 14170
rect 21226 14118 22816 14170
rect 1104 14096 22816 14118
rect 1854 14056 1860 14068
rect 1815 14028 1860 14056
rect 1854 14016 1860 14028
rect 1912 14016 1918 14068
rect 2590 14056 2596 14068
rect 2551 14028 2596 14056
rect 2590 14016 2596 14028
rect 2648 14016 2654 14068
rect 3694 14056 3700 14068
rect 3655 14028 3700 14056
rect 3694 14016 3700 14028
rect 3752 14016 3758 14068
rect 5902 14016 5908 14068
rect 5960 14056 5966 14068
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 5960 14028 6561 14056
rect 5960 14016 5966 14028
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 11054 14056 11060 14068
rect 11015 14028 11060 14056
rect 6549 14019 6607 14025
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 12158 14056 12164 14068
rect 12119 14028 12164 14056
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 13722 14056 13728 14068
rect 13683 14028 13728 14056
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 16758 14056 16764 14068
rect 16719 14028 16764 14056
rect 16758 14016 16764 14028
rect 16816 14016 16822 14068
rect 18046 14016 18052 14068
rect 18104 14056 18110 14068
rect 18782 14056 18788 14068
rect 18104 14028 18788 14056
rect 18104 14016 18110 14028
rect 18782 14016 18788 14028
rect 18840 14056 18846 14068
rect 19061 14059 19119 14065
rect 19061 14056 19073 14059
rect 18840 14028 19073 14056
rect 18840 14016 18846 14028
rect 19061 14025 19073 14028
rect 19107 14025 19119 14059
rect 19061 14019 19119 14025
rect 19702 14016 19708 14068
rect 19760 14056 19766 14068
rect 20073 14059 20131 14065
rect 20073 14056 20085 14059
rect 19760 14028 20085 14056
rect 19760 14016 19766 14028
rect 20073 14025 20085 14028
rect 20119 14025 20131 14059
rect 20073 14019 20131 14025
rect 2682 13948 2688 14000
rect 2740 13988 2746 14000
rect 5491 13991 5549 13997
rect 5491 13988 5503 13991
rect 2740 13960 5503 13988
rect 2740 13948 2746 13960
rect 5491 13957 5503 13960
rect 5537 13957 5549 13991
rect 5491 13951 5549 13957
rect 10134 13948 10140 14000
rect 10192 13988 10198 14000
rect 10321 13991 10379 13997
rect 10321 13988 10333 13991
rect 10192 13960 10333 13988
rect 10192 13948 10198 13960
rect 10321 13957 10333 13960
rect 10367 13988 10379 13991
rect 10367 13960 11928 13988
rect 10367 13957 10379 13960
rect 10321 13951 10379 13957
rect 11900 13932 11928 13960
rect 16666 13948 16672 14000
rect 16724 13988 16730 14000
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 16724 13960 17049 13988
rect 16724 13948 16730 13960
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 2314 13880 2320 13932
rect 2372 13920 2378 13932
rect 9306 13920 9312 13932
rect 2372 13892 9312 13920
rect 2372 13880 2378 13892
rect 9306 13880 9312 13892
rect 9364 13880 9370 13932
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13920 10747 13923
rect 11146 13920 11152 13932
rect 10735 13892 11152 13920
rect 10735 13889 10747 13892
rect 10689 13883 10747 13889
rect 11146 13880 11152 13892
rect 11204 13880 11210 13932
rect 11882 13920 11888 13932
rect 11795 13892 11888 13920
rect 11882 13880 11888 13892
rect 11940 13920 11946 13932
rect 15194 13920 15200 13932
rect 11940 13892 15200 13920
rect 11940 13880 11946 13892
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 15470 13920 15476 13932
rect 15431 13892 15476 13920
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 17972 13892 18920 13920
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13852 2283 13855
rect 2590 13852 2596 13864
rect 2271 13824 2596 13852
rect 2271 13821 2283 13824
rect 2225 13815 2283 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 3694 13812 3700 13864
rect 3752 13852 3758 13864
rect 3789 13855 3847 13861
rect 3789 13852 3801 13855
rect 3752 13824 3801 13852
rect 3752 13812 3758 13824
rect 3789 13821 3801 13824
rect 3835 13821 3847 13855
rect 3789 13815 3847 13821
rect 4341 13855 4399 13861
rect 4341 13821 4353 13855
rect 4387 13852 4399 13855
rect 4522 13852 4528 13864
rect 4387 13824 4528 13852
rect 4387 13821 4399 13824
rect 4341 13815 4399 13821
rect 4522 13812 4528 13824
rect 4580 13812 4586 13864
rect 5420 13855 5478 13861
rect 5420 13821 5432 13855
rect 5466 13852 5478 13855
rect 5718 13852 5724 13864
rect 5466 13824 5724 13852
rect 5466 13821 5478 13824
rect 5420 13815 5478 13821
rect 5718 13812 5724 13824
rect 5776 13852 5782 13864
rect 5813 13855 5871 13861
rect 5813 13852 5825 13855
rect 5776 13824 5825 13852
rect 5776 13812 5782 13824
rect 5813 13821 5825 13824
rect 5859 13821 5871 13855
rect 7466 13852 7472 13864
rect 7427 13824 7472 13852
rect 5813 13815 5871 13821
rect 7466 13812 7472 13824
rect 7524 13812 7530 13864
rect 10778 13852 10784 13864
rect 10739 13824 10784 13852
rect 10778 13812 10784 13824
rect 10836 13812 10842 13864
rect 10928 13855 10986 13861
rect 10928 13821 10940 13855
rect 10974 13852 10986 13855
rect 11514 13852 11520 13864
rect 10974 13824 11520 13852
rect 10974 13821 10986 13824
rect 10928 13815 10986 13821
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 12802 13852 12808 13864
rect 12763 13824 12808 13852
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 2038 13744 2044 13796
rect 2096 13784 2102 13796
rect 3970 13784 3976 13796
rect 2096 13756 3976 13784
rect 2096 13744 2102 13756
rect 3970 13744 3976 13756
rect 4028 13744 4034 13796
rect 9401 13787 9459 13793
rect 9401 13784 9413 13787
rect 9048 13756 9413 13784
rect 3329 13719 3387 13725
rect 3329 13685 3341 13719
rect 3375 13716 3387 13719
rect 4062 13716 4068 13728
rect 3375 13688 4068 13716
rect 3375 13685 3387 13688
rect 3329 13679 3387 13685
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 4154 13676 4160 13728
rect 4212 13716 4218 13728
rect 4338 13716 4344 13728
rect 4212 13688 4344 13716
rect 4212 13676 4218 13688
rect 4338 13676 4344 13688
rect 4396 13716 4402 13728
rect 4893 13719 4951 13725
rect 4893 13716 4905 13719
rect 4396 13688 4905 13716
rect 4396 13676 4402 13688
rect 4893 13685 4905 13688
rect 4939 13716 4951 13719
rect 6273 13719 6331 13725
rect 6273 13716 6285 13719
rect 4939 13688 6285 13716
rect 4939 13685 4951 13688
rect 4893 13679 4951 13685
rect 6273 13685 6285 13688
rect 6319 13716 6331 13719
rect 6362 13716 6368 13728
rect 6319 13688 6368 13716
rect 6319 13685 6331 13688
rect 6273 13679 6331 13685
rect 6362 13676 6368 13688
rect 6420 13716 6426 13728
rect 7377 13719 7435 13725
rect 7377 13716 7389 13719
rect 6420 13688 7389 13716
rect 6420 13676 6426 13688
rect 7377 13685 7389 13688
rect 7423 13716 7435 13719
rect 7837 13719 7895 13725
rect 7837 13716 7849 13719
rect 7423 13688 7849 13716
rect 7423 13685 7435 13688
rect 7377 13679 7435 13685
rect 7837 13685 7849 13688
rect 7883 13685 7895 13719
rect 7837 13679 7895 13685
rect 7926 13676 7932 13728
rect 7984 13716 7990 13728
rect 9048 13725 9076 13756
rect 9401 13753 9413 13756
rect 9447 13753 9459 13787
rect 9950 13784 9956 13796
rect 9911 13756 9956 13784
rect 9401 13747 9459 13753
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 14734 13784 14740 13796
rect 11440 13756 14740 13784
rect 8389 13719 8447 13725
rect 8389 13716 8401 13719
rect 7984 13688 8401 13716
rect 7984 13676 7990 13688
rect 8389 13685 8401 13688
rect 8435 13716 8447 13719
rect 9033 13719 9091 13725
rect 9033 13716 9045 13719
rect 8435 13688 9045 13716
rect 8435 13685 8447 13688
rect 8389 13679 8447 13685
rect 9033 13685 9045 13688
rect 9079 13685 9091 13719
rect 9033 13679 9091 13685
rect 10226 13676 10232 13728
rect 10284 13716 10290 13728
rect 10594 13716 10600 13728
rect 10284 13688 10600 13716
rect 10284 13676 10290 13688
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 11440 13725 11468 13756
rect 14734 13744 14740 13756
rect 14792 13744 14798 13796
rect 15794 13787 15852 13793
rect 15794 13753 15806 13787
rect 15840 13753 15852 13787
rect 15794 13747 15852 13753
rect 17497 13787 17555 13793
rect 17497 13753 17509 13787
rect 17543 13784 17555 13787
rect 17972 13784 18000 13892
rect 18141 13787 18199 13793
rect 18141 13784 18153 13787
rect 17543 13756 18153 13784
rect 17543 13753 17555 13756
rect 17497 13747 17555 13753
rect 18141 13753 18153 13756
rect 18187 13753 18199 13787
rect 18141 13747 18199 13753
rect 18233 13787 18291 13793
rect 18233 13753 18245 13787
rect 18279 13784 18291 13787
rect 18414 13784 18420 13796
rect 18279 13756 18420 13784
rect 18279 13753 18291 13756
rect 18233 13747 18291 13753
rect 11425 13719 11483 13725
rect 11425 13685 11437 13719
rect 11471 13685 11483 13719
rect 11425 13679 11483 13685
rect 13173 13719 13231 13725
rect 13173 13685 13185 13719
rect 13219 13716 13231 13719
rect 13262 13716 13268 13728
rect 13219 13688 13268 13716
rect 13219 13685 13231 13688
rect 13173 13679 13231 13685
rect 13262 13676 13268 13688
rect 13320 13676 13326 13728
rect 15381 13719 15439 13725
rect 15381 13685 15393 13719
rect 15427 13716 15439 13719
rect 15809 13716 15837 13747
rect 15930 13716 15936 13728
rect 15427 13688 15936 13716
rect 15427 13685 15439 13688
rect 15381 13679 15439 13685
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 16393 13719 16451 13725
rect 16393 13685 16405 13719
rect 16439 13716 16451 13719
rect 17402 13716 17408 13728
rect 16439 13688 17408 13716
rect 16439 13685 16451 13688
rect 16393 13679 16451 13685
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 17865 13719 17923 13725
rect 17865 13685 17877 13719
rect 17911 13716 17923 13719
rect 18248 13716 18276 13747
rect 18414 13744 18420 13756
rect 18472 13744 18478 13796
rect 18506 13744 18512 13796
rect 18564 13784 18570 13796
rect 18782 13784 18788 13796
rect 18564 13756 18788 13784
rect 18564 13744 18570 13756
rect 18782 13744 18788 13756
rect 18840 13744 18846 13796
rect 18892 13784 18920 13892
rect 19613 13787 19671 13793
rect 19613 13784 19625 13787
rect 18892 13756 19625 13784
rect 19613 13753 19625 13756
rect 19659 13753 19671 13787
rect 19613 13747 19671 13753
rect 17911 13688 18276 13716
rect 17911 13685 17923 13688
rect 17865 13679 17923 13685
rect 1104 13626 22816 13648
rect 1104 13574 8982 13626
rect 9034 13574 9046 13626
rect 9098 13574 9110 13626
rect 9162 13574 9174 13626
rect 9226 13574 16982 13626
rect 17034 13574 17046 13626
rect 17098 13574 17110 13626
rect 17162 13574 17174 13626
rect 17226 13574 22816 13626
rect 1104 13552 22816 13574
rect 1765 13515 1823 13521
rect 1765 13481 1777 13515
rect 1811 13512 1823 13515
rect 1854 13512 1860 13524
rect 1811 13484 1860 13512
rect 1811 13481 1823 13484
rect 1765 13475 1823 13481
rect 1854 13472 1860 13484
rect 1912 13472 1918 13524
rect 3234 13512 3240 13524
rect 2240 13484 3240 13512
rect 2240 13453 2268 13484
rect 3234 13472 3240 13484
rect 3292 13472 3298 13524
rect 3418 13472 3424 13524
rect 3476 13512 3482 13524
rect 4157 13515 4215 13521
rect 4157 13512 4169 13515
rect 3476 13484 4169 13512
rect 3476 13472 3482 13484
rect 4157 13481 4169 13484
rect 4203 13481 4215 13515
rect 4157 13475 4215 13481
rect 5902 13472 5908 13524
rect 5960 13512 5966 13524
rect 6089 13515 6147 13521
rect 6089 13512 6101 13515
rect 5960 13484 6101 13512
rect 5960 13472 5966 13484
rect 6089 13481 6101 13484
rect 6135 13481 6147 13515
rect 7466 13512 7472 13524
rect 7427 13484 7472 13512
rect 6089 13475 6147 13481
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 9306 13512 9312 13524
rect 9267 13484 9312 13512
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 10778 13512 10784 13524
rect 10192 13484 10784 13512
rect 10192 13472 10198 13484
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 11514 13512 11520 13524
rect 11475 13484 11520 13512
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 12989 13515 13047 13521
rect 12989 13512 13001 13515
rect 12860 13484 13001 13512
rect 12860 13472 12866 13484
rect 12989 13481 13001 13484
rect 13035 13481 13047 13515
rect 12989 13475 13047 13481
rect 13357 13515 13415 13521
rect 13357 13481 13369 13515
rect 13403 13512 13415 13515
rect 13446 13512 13452 13524
rect 13403 13484 13452 13512
rect 13403 13481 13415 13484
rect 13357 13475 13415 13481
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 16393 13515 16451 13521
rect 16393 13481 16405 13515
rect 16439 13512 16451 13515
rect 16758 13512 16764 13524
rect 16439 13484 16764 13512
rect 16439 13481 16451 13484
rect 16393 13475 16451 13481
rect 16758 13472 16764 13484
rect 16816 13472 16822 13524
rect 2225 13447 2283 13453
rect 2225 13413 2237 13447
rect 2271 13413 2283 13447
rect 2225 13407 2283 13413
rect 2317 13447 2375 13453
rect 2317 13413 2329 13447
rect 2363 13444 2375 13447
rect 2682 13444 2688 13456
rect 2363 13416 2688 13444
rect 2363 13413 2375 13416
rect 2317 13407 2375 13413
rect 2682 13404 2688 13416
rect 2740 13404 2746 13456
rect 3694 13404 3700 13456
rect 3752 13444 3758 13456
rect 10870 13444 10876 13456
rect 3752 13416 6132 13444
rect 3752 13404 3758 13416
rect 6104 13388 6132 13416
rect 10520 13416 10876 13444
rect 10520 13388 10548 13416
rect 10870 13404 10876 13416
rect 10928 13404 10934 13456
rect 12066 13404 12072 13456
rect 12124 13444 12130 13456
rect 12390 13447 12448 13453
rect 12390 13444 12402 13447
rect 12124 13416 12402 13444
rect 12124 13404 12130 13416
rect 12390 13413 12402 13416
rect 12436 13413 12448 13447
rect 12390 13407 12448 13413
rect 15835 13447 15893 13453
rect 15835 13413 15847 13447
rect 15881 13444 15893 13447
rect 15930 13444 15936 13456
rect 15881 13416 15936 13444
rect 15881 13413 15893 13416
rect 15835 13407 15893 13413
rect 15930 13404 15936 13416
rect 15988 13404 15994 13456
rect 17402 13404 17408 13456
rect 17460 13444 17466 13456
rect 17957 13447 18015 13453
rect 17957 13444 17969 13447
rect 17460 13416 17969 13444
rect 17460 13404 17466 13416
rect 17957 13413 17969 13416
rect 18003 13444 18015 13447
rect 18046 13444 18052 13456
rect 18003 13416 18052 13444
rect 18003 13413 18015 13416
rect 17957 13407 18015 13413
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 18509 13447 18567 13453
rect 18509 13413 18521 13447
rect 18555 13444 18567 13447
rect 18782 13444 18788 13456
rect 18555 13416 18788 13444
rect 18555 13413 18567 13416
rect 18509 13407 18567 13413
rect 18782 13404 18788 13416
rect 18840 13404 18846 13456
rect 4341 13379 4399 13385
rect 4341 13345 4353 13379
rect 4387 13345 4399 13379
rect 4614 13376 4620 13388
rect 4575 13348 4620 13376
rect 4341 13339 4399 13345
rect 2314 13268 2320 13320
rect 2372 13308 2378 13320
rect 2501 13311 2559 13317
rect 2501 13308 2513 13311
rect 2372 13280 2513 13308
rect 2372 13268 2378 13280
rect 2501 13277 2513 13280
rect 2547 13277 2559 13311
rect 2501 13271 2559 13277
rect 3326 13268 3332 13320
rect 3384 13308 3390 13320
rect 3878 13308 3884 13320
rect 3384 13280 3884 13308
rect 3384 13268 3390 13280
rect 3878 13268 3884 13280
rect 3936 13308 3942 13320
rect 4356 13308 4384 13339
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 6086 13376 6092 13388
rect 6047 13348 6092 13376
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 6549 13379 6607 13385
rect 6549 13345 6561 13379
rect 6595 13376 6607 13379
rect 6595 13348 7144 13376
rect 6595 13345 6607 13348
rect 6549 13339 6607 13345
rect 6454 13308 6460 13320
rect 3936 13280 6460 13308
rect 3936 13268 3942 13280
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 3878 13172 3884 13184
rect 3839 13144 3884 13172
rect 3878 13132 3884 13144
rect 3936 13132 3942 13184
rect 7116 13181 7144 13348
rect 7926 13336 7932 13388
rect 7984 13376 7990 13388
rect 8113 13379 8171 13385
rect 8113 13376 8125 13379
rect 7984 13348 8125 13376
rect 7984 13336 7990 13348
rect 8113 13345 8125 13348
rect 8159 13345 8171 13379
rect 10502 13376 10508 13388
rect 10463 13348 10508 13376
rect 8113 13339 8171 13345
rect 10502 13336 10508 13348
rect 10560 13336 10566 13388
rect 10778 13336 10784 13388
rect 10836 13376 10842 13388
rect 11057 13379 11115 13385
rect 11057 13376 11069 13379
rect 10836 13348 11069 13376
rect 10836 13336 10842 13348
rect 11057 13345 11069 13348
rect 11103 13376 11115 13379
rect 12158 13376 12164 13388
rect 11103 13348 12164 13376
rect 11103 13345 11115 13348
rect 11057 13339 11115 13345
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13308 11299 13311
rect 12069 13311 12127 13317
rect 12069 13308 12081 13311
rect 11287 13280 12081 13308
rect 11287 13277 11299 13280
rect 11241 13271 11299 13277
rect 12069 13277 12081 13280
rect 12115 13308 12127 13311
rect 12618 13308 12624 13320
rect 12115 13280 12624 13308
rect 12115 13277 12127 13280
rect 12069 13271 12127 13277
rect 12618 13268 12624 13280
rect 12676 13268 12682 13320
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 15470 13308 15476 13320
rect 13872 13280 13917 13308
rect 15431 13280 15476 13308
rect 13872 13268 13878 13280
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 17310 13268 17316 13320
rect 17368 13308 17374 13320
rect 17865 13311 17923 13317
rect 17865 13308 17877 13311
rect 17368 13280 17877 13308
rect 17368 13268 17374 13280
rect 17865 13277 17877 13280
rect 17911 13308 17923 13311
rect 18690 13308 18696 13320
rect 17911 13280 18696 13308
rect 17911 13277 17923 13280
rect 17865 13271 17923 13277
rect 18690 13268 18696 13280
rect 18748 13268 18754 13320
rect 7101 13175 7159 13181
rect 7101 13141 7113 13175
rect 7147 13172 7159 13175
rect 7282 13172 7288 13184
rect 7147 13144 7288 13172
rect 7147 13141 7159 13144
rect 7101 13135 7159 13141
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 8478 13172 8484 13184
rect 8439 13144 8484 13172
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 10229 13175 10287 13181
rect 10229 13141 10241 13175
rect 10275 13172 10287 13175
rect 10410 13172 10416 13184
rect 10275 13144 10416 13172
rect 10275 13141 10287 13144
rect 10229 13135 10287 13141
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 1104 13082 22816 13104
rect 1104 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 12982 13082
rect 13034 13030 13046 13082
rect 13098 13030 13110 13082
rect 13162 13030 13174 13082
rect 13226 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 22816 13082
rect 1104 13008 22816 13030
rect 3326 12968 3332 12980
rect 3287 12940 3332 12968
rect 3326 12928 3332 12940
rect 3384 12928 3390 12980
rect 3878 12928 3884 12980
rect 3936 12968 3942 12980
rect 4614 12968 4620 12980
rect 3936 12940 4620 12968
rect 3936 12928 3942 12940
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 8110 12968 8116 12980
rect 8071 12940 8116 12968
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 8478 12968 8484 12980
rect 8439 12940 8484 12968
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 8570 12928 8576 12980
rect 8628 12968 8634 12980
rect 10302 12971 10360 12977
rect 10302 12968 10314 12971
rect 8628 12940 10314 12968
rect 8628 12928 8634 12940
rect 10302 12937 10314 12940
rect 10348 12968 10360 12971
rect 10778 12968 10784 12980
rect 10348 12940 10548 12968
rect 10739 12940 10784 12968
rect 10348 12937 10360 12940
rect 10302 12931 10360 12937
rect 4065 12903 4123 12909
rect 4065 12869 4077 12903
rect 4111 12900 4123 12903
rect 4338 12900 4344 12912
rect 4111 12872 4344 12900
rect 4111 12869 4123 12872
rect 4065 12863 4123 12869
rect 4338 12860 4344 12872
rect 4396 12900 4402 12912
rect 4433 12903 4491 12909
rect 4433 12900 4445 12903
rect 4396 12872 4445 12900
rect 4396 12860 4402 12872
rect 4433 12869 4445 12872
rect 4479 12900 4491 12903
rect 6270 12900 6276 12912
rect 4479 12872 6276 12900
rect 4479 12869 4491 12872
rect 4433 12863 4491 12869
rect 6270 12860 6276 12872
rect 6328 12860 6334 12912
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 4522 12832 4528 12844
rect 3743 12804 4528 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 7466 12832 7472 12844
rect 7427 12804 7472 12832
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 8128 12832 8156 12928
rect 10413 12903 10471 12909
rect 10413 12869 10425 12903
rect 10459 12869 10471 12903
rect 10520 12900 10548 12940
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 11514 12968 11520 12980
rect 11475 12940 11520 12968
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 12066 12968 12072 12980
rect 12027 12940 12072 12968
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 12618 12968 12624 12980
rect 12579 12940 12624 12968
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 12802 12928 12808 12980
rect 12860 12968 12866 12980
rect 12989 12971 13047 12977
rect 12989 12968 13001 12971
rect 12860 12940 13001 12968
rect 12860 12928 12866 12940
rect 12989 12937 13001 12940
rect 13035 12937 13047 12971
rect 12989 12931 13047 12937
rect 16301 12971 16359 12977
rect 16301 12937 16313 12971
rect 16347 12968 16359 12971
rect 16758 12968 16764 12980
rect 16347 12940 16764 12968
rect 16347 12937 16359 12940
rect 16301 12931 16359 12937
rect 11532 12900 11560 12928
rect 10520 12872 11560 12900
rect 10413 12863 10471 12869
rect 8665 12835 8723 12841
rect 8665 12832 8677 12835
rect 8128 12804 8677 12832
rect 8665 12801 8677 12804
rect 8711 12801 8723 12835
rect 10428 12832 10456 12863
rect 8665 12795 8723 12801
rect 10336 12804 10456 12832
rect 10505 12835 10563 12841
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12764 1915 12767
rect 3418 12764 3424 12776
rect 1903 12736 3424 12764
rect 1903 12733 1915 12736
rect 1857 12727 1915 12733
rect 3418 12724 3424 12736
rect 3476 12724 3482 12776
rect 4304 12767 4362 12773
rect 4304 12733 4316 12767
rect 4350 12764 4362 12767
rect 5629 12767 5687 12773
rect 4350 12736 5304 12764
rect 4350 12733 4362 12736
rect 4304 12727 4362 12733
rect 1765 12699 1823 12705
rect 1765 12665 1777 12699
rect 1811 12696 1823 12699
rect 2038 12696 2044 12708
rect 1811 12668 2044 12696
rect 1811 12665 1823 12668
rect 1765 12659 1823 12665
rect 2038 12656 2044 12668
rect 2096 12696 2102 12708
rect 2178 12699 2236 12705
rect 2178 12696 2190 12699
rect 2096 12668 2190 12696
rect 2096 12656 2102 12668
rect 2178 12665 2190 12668
rect 2224 12696 2236 12699
rect 2406 12696 2412 12708
rect 2224 12668 2412 12696
rect 2224 12665 2236 12668
rect 2178 12659 2236 12665
rect 2406 12656 2412 12668
rect 2464 12656 2470 12708
rect 4154 12656 4160 12708
rect 4212 12696 4218 12708
rect 4212 12668 4257 12696
rect 4212 12656 4218 12668
rect 2774 12628 2780 12640
rect 2735 12600 2780 12628
rect 2774 12588 2780 12600
rect 2832 12588 2838 12640
rect 5276 12637 5304 12736
rect 5629 12733 5641 12767
rect 5675 12764 5687 12767
rect 6178 12764 6184 12776
rect 5675 12736 6184 12764
rect 5675 12733 5687 12736
rect 5629 12727 5687 12733
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6564 12736 6837 12764
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5350 12628 5356 12640
rect 5307 12600 5356 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 5718 12628 5724 12640
rect 5679 12600 5724 12628
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 6086 12588 6092 12640
rect 6144 12628 6150 12640
rect 6181 12631 6239 12637
rect 6181 12628 6193 12631
rect 6144 12600 6193 12628
rect 6144 12588 6150 12600
rect 6181 12597 6193 12600
rect 6227 12597 6239 12631
rect 6181 12591 6239 12597
rect 6454 12588 6460 12640
rect 6512 12628 6518 12640
rect 6564 12637 6592 12736
rect 6825 12733 6837 12736
rect 6871 12733 6883 12767
rect 7282 12764 7288 12776
rect 7243 12736 7288 12764
rect 6825 12727 6883 12733
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12764 9367 12767
rect 9950 12764 9956 12776
rect 9355 12736 9956 12764
rect 9355 12733 9367 12736
rect 9309 12727 9367 12733
rect 9950 12724 9956 12736
rect 10008 12764 10014 12776
rect 10226 12764 10232 12776
rect 10008 12736 10232 12764
rect 10008 12724 10014 12736
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 8757 12699 8815 12705
rect 8757 12665 8769 12699
rect 8803 12665 8815 12699
rect 10134 12696 10140 12708
rect 8757 12659 8815 12665
rect 9600 12668 10140 12696
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 6512 12600 6561 12628
rect 6512 12588 6518 12600
rect 6549 12597 6561 12600
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 8478 12588 8484 12640
rect 8536 12628 8542 12640
rect 8772 12628 8800 12659
rect 9600 12640 9628 12668
rect 10134 12656 10140 12668
rect 10192 12656 10198 12708
rect 10336 12640 10364 12804
rect 10505 12801 10517 12835
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 10410 12724 10416 12776
rect 10468 12764 10474 12776
rect 10520 12764 10548 12795
rect 10468 12736 10548 12764
rect 10468 12724 10474 12736
rect 13004 12696 13032 12931
rect 16758 12928 16764 12940
rect 16816 12928 16822 12980
rect 17402 12968 17408 12980
rect 17363 12940 17408 12968
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 18690 12900 18696 12912
rect 18651 12872 18696 12900
rect 18690 12860 18696 12872
rect 18748 12900 18754 12912
rect 19429 12903 19487 12909
rect 19429 12900 19441 12903
rect 18748 12872 19441 12900
rect 18748 12860 18754 12872
rect 19429 12869 19441 12872
rect 19475 12869 19487 12903
rect 19429 12863 19487 12869
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12832 13323 12835
rect 13446 12832 13452 12844
rect 13311 12804 13452 12832
rect 13311 12801 13323 12804
rect 13265 12795 13323 12801
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 13722 12832 13728 12844
rect 13683 12804 13728 12832
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 15378 12832 15384 12844
rect 15339 12804 15384 12832
rect 15378 12792 15384 12804
rect 15436 12792 15442 12844
rect 18138 12832 18144 12844
rect 18051 12804 18144 12832
rect 18138 12792 18144 12804
rect 18196 12832 18202 12844
rect 19061 12835 19119 12841
rect 19061 12832 19073 12835
rect 18196 12804 19073 12832
rect 18196 12792 18202 12804
rect 19061 12801 19073 12804
rect 19107 12801 19119 12835
rect 19061 12795 19119 12801
rect 14645 12767 14703 12773
rect 14645 12733 14657 12767
rect 14691 12764 14703 12767
rect 14737 12767 14795 12773
rect 14737 12764 14749 12767
rect 14691 12736 14749 12764
rect 14691 12733 14703 12736
rect 14645 12727 14703 12733
rect 14737 12733 14749 12736
rect 14783 12733 14795 12767
rect 14737 12727 14795 12733
rect 13357 12699 13415 12705
rect 13357 12696 13369 12699
rect 13004 12668 13369 12696
rect 13357 12665 13369 12668
rect 13403 12665 13415 12699
rect 13357 12659 13415 12665
rect 9582 12628 9588 12640
rect 8536 12600 8800 12628
rect 9543 12600 9588 12628
rect 8536 12588 8542 12600
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 10045 12631 10103 12637
rect 10045 12597 10057 12631
rect 10091 12628 10103 12631
rect 10318 12628 10324 12640
rect 10091 12600 10324 12628
rect 10091 12597 10103 12600
rect 10045 12591 10103 12597
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 10502 12588 10508 12640
rect 10560 12628 10566 12640
rect 11149 12631 11207 12637
rect 11149 12628 11161 12631
rect 10560 12600 11161 12628
rect 10560 12588 10566 12600
rect 11149 12597 11161 12600
rect 11195 12597 11207 12631
rect 11149 12591 11207 12597
rect 13446 12588 13452 12640
rect 13504 12628 13510 12640
rect 14660 12628 14688 12727
rect 14826 12724 14832 12776
rect 14884 12764 14890 12776
rect 15197 12767 15255 12773
rect 15197 12764 15209 12767
rect 14884 12736 15209 12764
rect 14884 12724 14890 12736
rect 15197 12733 15209 12736
rect 15243 12733 15255 12767
rect 16758 12764 16764 12776
rect 16719 12736 16764 12764
rect 15197 12727 15255 12733
rect 16758 12724 16764 12736
rect 16816 12724 16822 12776
rect 17129 12699 17187 12705
rect 17129 12665 17141 12699
rect 17175 12696 17187 12699
rect 17773 12699 17831 12705
rect 17773 12696 17785 12699
rect 17175 12668 17785 12696
rect 17175 12665 17187 12668
rect 17129 12659 17187 12665
rect 17773 12665 17785 12668
rect 17819 12665 17831 12699
rect 17773 12659 17831 12665
rect 18233 12699 18291 12705
rect 18233 12665 18245 12699
rect 18279 12665 18291 12699
rect 18233 12659 18291 12665
rect 13504 12600 14688 12628
rect 15841 12631 15899 12637
rect 13504 12588 13510 12600
rect 15841 12597 15853 12631
rect 15887 12628 15899 12631
rect 15930 12628 15936 12640
rect 15887 12600 15936 12628
rect 15887 12597 15899 12600
rect 15841 12591 15899 12597
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 17788 12628 17816 12659
rect 18248 12628 18276 12659
rect 17788 12600 18276 12628
rect 1104 12538 22816 12560
rect 1104 12486 8982 12538
rect 9034 12486 9046 12538
rect 9098 12486 9110 12538
rect 9162 12486 9174 12538
rect 9226 12486 16982 12538
rect 17034 12486 17046 12538
rect 17098 12486 17110 12538
rect 17162 12486 17174 12538
rect 17226 12486 22816 12538
rect 1104 12464 22816 12486
rect 3145 12427 3203 12433
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 3418 12424 3424 12436
rect 3191 12396 3424 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 3878 12424 3884 12436
rect 3839 12396 3884 12424
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 7926 12424 7932 12436
rect 7887 12396 7932 12424
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 8662 12424 8668 12436
rect 8623 12396 8668 12424
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 10686 12424 10692 12436
rect 10647 12396 10692 12424
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 10778 12384 10784 12436
rect 10836 12424 10842 12436
rect 11057 12427 11115 12433
rect 11057 12424 11069 12427
rect 10836 12396 11069 12424
rect 10836 12384 10842 12396
rect 11057 12393 11069 12396
rect 11103 12393 11115 12427
rect 11057 12387 11115 12393
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 12492 12396 12633 12424
rect 12492 12384 12498 12396
rect 12621 12393 12633 12396
rect 12667 12424 12679 12427
rect 14734 12424 14740 12436
rect 12667 12396 13676 12424
rect 14695 12396 14740 12424
rect 12667 12393 12679 12396
rect 12621 12387 12679 12393
rect 1857 12359 1915 12365
rect 1857 12325 1869 12359
rect 1903 12356 1915 12359
rect 2038 12356 2044 12368
rect 1903 12328 2044 12356
rect 1903 12325 1915 12328
rect 1857 12319 1915 12325
rect 2038 12316 2044 12328
rect 2096 12356 2102 12368
rect 4065 12359 4123 12365
rect 4065 12356 4077 12359
rect 2096 12328 4077 12356
rect 2096 12316 2102 12328
rect 4065 12325 4077 12328
rect 4111 12325 4123 12359
rect 8021 12359 8079 12365
rect 8021 12356 8033 12359
rect 4065 12319 4123 12325
rect 6380 12328 8033 12356
rect 2774 12288 2780 12300
rect 2687 12260 2780 12288
rect 2774 12248 2780 12260
rect 2832 12288 2838 12300
rect 4614 12288 4620 12300
rect 2832 12260 4620 12288
rect 2832 12248 2838 12260
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 6178 12248 6184 12300
rect 6236 12288 6242 12300
rect 6380 12297 6408 12328
rect 8021 12325 8033 12328
rect 8067 12356 8079 12359
rect 9582 12356 9588 12368
rect 8067 12328 9588 12356
rect 8067 12325 8079 12328
rect 8021 12319 8079 12325
rect 9582 12316 9588 12328
rect 9640 12316 9646 12368
rect 13081 12359 13139 12365
rect 13081 12325 13093 12359
rect 13127 12356 13139 12359
rect 13262 12356 13268 12368
rect 13127 12328 13268 12356
rect 13127 12325 13139 12328
rect 13081 12319 13139 12325
rect 13262 12316 13268 12328
rect 13320 12316 13326 12368
rect 13648 12365 13676 12396
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 15565 12427 15623 12433
rect 15565 12424 15577 12427
rect 15528 12396 15577 12424
rect 15528 12384 15534 12396
rect 15565 12393 15577 12396
rect 15611 12424 15623 12427
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 15611 12396 16313 12424
rect 15611 12393 15623 12396
rect 15565 12387 15623 12393
rect 16301 12393 16313 12396
rect 16347 12393 16359 12427
rect 16301 12387 16359 12393
rect 17727 12427 17785 12433
rect 17727 12393 17739 12427
rect 17773 12424 17785 12427
rect 18138 12424 18144 12436
rect 17773 12396 18144 12424
rect 17773 12393 17785 12396
rect 17727 12387 17785 12393
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 21082 12424 21088 12436
rect 21043 12396 21088 12424
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 13633 12359 13691 12365
rect 13633 12325 13645 12359
rect 13679 12356 13691 12359
rect 13722 12356 13728 12368
rect 13679 12328 13728 12356
rect 13679 12325 13691 12328
rect 13633 12319 13691 12325
rect 13722 12316 13728 12328
rect 13780 12316 13786 12368
rect 14752 12356 14780 12384
rect 18785 12359 18843 12365
rect 14752 12328 15792 12356
rect 6365 12291 6423 12297
rect 6365 12288 6377 12291
rect 6236 12260 6377 12288
rect 6236 12248 6242 12260
rect 6365 12257 6377 12260
rect 6411 12257 6423 12291
rect 6365 12251 6423 12257
rect 6546 12248 6552 12300
rect 6604 12288 6610 12300
rect 6604 12260 7833 12288
rect 6604 12248 6610 12260
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12220 1823 12223
rect 1946 12220 1952 12232
rect 1811 12192 1952 12220
rect 1811 12189 1823 12192
rect 1765 12183 1823 12189
rect 1946 12180 1952 12192
rect 2004 12220 2010 12232
rect 5718 12220 5724 12232
rect 2004 12192 5724 12220
rect 2004 12180 2010 12192
rect 5718 12180 5724 12192
rect 5776 12180 5782 12232
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 6733 12223 6791 12229
rect 6733 12220 6745 12223
rect 6696 12192 6745 12220
rect 6696 12180 6702 12192
rect 6733 12189 6745 12192
rect 6779 12189 6791 12223
rect 7805 12220 7833 12260
rect 9490 12248 9496 12300
rect 9548 12288 9554 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 9548 12260 10057 12288
rect 9548 12248 9554 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 10045 12251 10103 12257
rect 10226 12248 10232 12300
rect 10284 12288 10290 12300
rect 11676 12291 11734 12297
rect 11676 12288 11688 12291
rect 10284 12260 11688 12288
rect 10284 12248 10290 12260
rect 11676 12257 11688 12260
rect 11722 12288 11734 12291
rect 12069 12291 12127 12297
rect 12069 12288 12081 12291
rect 11722 12260 12081 12288
rect 11722 12257 11734 12260
rect 11676 12251 11734 12257
rect 12069 12257 12081 12260
rect 12115 12257 12127 12291
rect 12069 12251 12127 12257
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 15764 12297 15792 12328
rect 18785 12325 18797 12359
rect 18831 12356 18843 12359
rect 19426 12356 19432 12368
rect 18831 12328 19432 12356
rect 18831 12325 18843 12328
rect 18785 12319 18843 12325
rect 19426 12316 19432 12328
rect 19484 12316 19490 12368
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 15252 12260 15301 12288
rect 15252 12248 15258 12260
rect 15289 12257 15301 12260
rect 15335 12257 15347 12291
rect 15289 12251 15347 12257
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 16666 12288 16672 12300
rect 15795 12260 16672 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 17589 12291 17647 12297
rect 17589 12257 17601 12291
rect 17635 12288 17647 12291
rect 17678 12288 17684 12300
rect 17635 12260 17684 12288
rect 17635 12257 17647 12260
rect 17589 12251 17647 12257
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 20806 12248 20812 12300
rect 20864 12288 20870 12300
rect 20901 12291 20959 12297
rect 20901 12288 20913 12291
rect 20864 12260 20913 12288
rect 20864 12248 20870 12260
rect 20901 12257 20913 12260
rect 20947 12257 20959 12291
rect 20901 12251 20959 12257
rect 8110 12220 8116 12232
rect 7805 12192 8116 12220
rect 6733 12183 6791 12189
rect 8110 12180 8116 12192
rect 8168 12229 8174 12232
rect 8168 12223 8226 12229
rect 8168 12189 8180 12223
rect 8214 12189 8226 12223
rect 8386 12220 8392 12232
rect 8347 12192 8392 12220
rect 8168 12183 8226 12189
rect 8168 12180 8174 12183
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 10410 12220 10416 12232
rect 10371 12192 10416 12220
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12220 13047 12223
rect 13354 12220 13360 12232
rect 13035 12192 13360 12220
rect 13035 12189 13047 12192
rect 12989 12183 13047 12189
rect 13354 12180 13360 12192
rect 13412 12220 13418 12232
rect 13814 12220 13820 12232
rect 13412 12192 13820 12220
rect 13412 12180 13418 12192
rect 13814 12180 13820 12192
rect 13872 12180 13878 12232
rect 18690 12220 18696 12232
rect 18651 12192 18696 12220
rect 18690 12180 18696 12192
rect 18748 12180 18754 12232
rect 18966 12220 18972 12232
rect 18927 12192 18972 12220
rect 18966 12180 18972 12192
rect 19024 12180 19030 12232
rect 2314 12152 2320 12164
rect 2275 12124 2320 12152
rect 2314 12112 2320 12124
rect 2372 12112 2378 12164
rect 5350 12112 5356 12164
rect 5408 12152 5414 12164
rect 5905 12155 5963 12161
rect 5408 12124 5764 12152
rect 5408 12112 5414 12124
rect 5736 12096 5764 12124
rect 5905 12121 5917 12155
rect 5951 12152 5963 12155
rect 6825 12155 6883 12161
rect 6825 12152 6837 12155
rect 5951 12124 6837 12152
rect 5951 12121 5963 12124
rect 5905 12115 5963 12121
rect 6825 12121 6837 12124
rect 6871 12152 6883 12155
rect 7282 12152 7288 12164
rect 6871 12124 7288 12152
rect 6871 12121 6883 12124
rect 6825 12115 6883 12121
rect 7282 12112 7288 12124
rect 7340 12112 7346 12164
rect 11514 12152 11520 12164
rect 10198 12124 11520 12152
rect 10198 12096 10226 12124
rect 11514 12112 11520 12124
rect 11572 12112 11578 12164
rect 11747 12155 11805 12161
rect 11747 12121 11759 12155
rect 11793 12152 11805 12155
rect 20714 12152 20720 12164
rect 11793 12124 12801 12152
rect 11793 12121 11805 12124
rect 11747 12115 11805 12121
rect 5261 12087 5319 12093
rect 5261 12053 5273 12087
rect 5307 12084 5319 12087
rect 5626 12084 5632 12096
rect 5307 12056 5632 12084
rect 5307 12053 5319 12056
rect 5261 12047 5319 12053
rect 5626 12044 5632 12056
rect 5684 12044 5690 12096
rect 5718 12044 5724 12096
rect 5776 12084 5782 12096
rect 6546 12093 6552 12096
rect 6181 12087 6239 12093
rect 6181 12084 6193 12087
rect 5776 12056 6193 12084
rect 5776 12044 5782 12056
rect 6181 12053 6193 12056
rect 6227 12084 6239 12087
rect 6503 12087 6552 12093
rect 6503 12084 6515 12087
rect 6227 12056 6515 12084
rect 6227 12053 6239 12056
rect 6181 12047 6239 12053
rect 6503 12053 6515 12056
rect 6549 12053 6552 12087
rect 6503 12047 6552 12053
rect 6546 12044 6552 12047
rect 6604 12044 6610 12096
rect 6641 12087 6699 12093
rect 6641 12053 6653 12087
rect 6687 12084 6699 12087
rect 7098 12084 7104 12096
rect 6687 12056 7104 12084
rect 6687 12053 6699 12056
rect 6641 12047 6699 12053
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 7374 12084 7380 12096
rect 7335 12056 7380 12084
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 8294 12084 8300 12096
rect 8255 12056 8300 12084
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 9122 12084 9128 12096
rect 9083 12056 9128 12084
rect 9122 12044 9128 12056
rect 9180 12044 9186 12096
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 10198 12093 10232 12096
rect 9861 12087 9919 12093
rect 9861 12084 9873 12087
rect 9456 12056 9873 12084
rect 9456 12044 9462 12056
rect 9861 12053 9873 12056
rect 9907 12084 9919 12087
rect 10183 12087 10232 12093
rect 10183 12084 10195 12087
rect 9907 12056 10195 12084
rect 9907 12053 9919 12056
rect 9861 12047 9919 12053
rect 10183 12053 10195 12056
rect 10229 12053 10232 12087
rect 10183 12047 10232 12053
rect 10226 12044 10232 12047
rect 10284 12044 10290 12096
rect 10318 12044 10324 12096
rect 10376 12084 10382 12096
rect 12773 12084 12801 12124
rect 13786 12124 20720 12152
rect 13786 12084 13814 12124
rect 20714 12112 20720 12124
rect 20772 12112 20778 12164
rect 13998 12084 14004 12096
rect 10376 12056 10421 12084
rect 12773 12056 13814 12084
rect 13959 12056 14004 12084
rect 10376 12044 10382 12056
rect 13998 12044 14004 12056
rect 14056 12044 14062 12096
rect 18325 12087 18383 12093
rect 18325 12053 18337 12087
rect 18371 12084 18383 12087
rect 18414 12084 18420 12096
rect 18371 12056 18420 12084
rect 18371 12053 18383 12056
rect 18325 12047 18383 12053
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 1104 11994 22816 12016
rect 1104 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 12982 11994
rect 13034 11942 13046 11994
rect 13098 11942 13110 11994
rect 13162 11942 13174 11994
rect 13226 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 22816 11994
rect 1104 11920 22816 11942
rect 2038 11880 2044 11892
rect 1999 11852 2044 11880
rect 2038 11840 2044 11852
rect 2096 11840 2102 11892
rect 4614 11880 4620 11892
rect 4575 11852 4620 11880
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 10413 11883 10471 11889
rect 10413 11880 10425 11883
rect 10100 11852 10425 11880
rect 10100 11840 10106 11852
rect 10413 11849 10425 11852
rect 10459 11849 10471 11883
rect 10594 11880 10600 11892
rect 10555 11852 10600 11880
rect 10413 11843 10471 11849
rect 10594 11840 10600 11852
rect 10652 11840 10658 11892
rect 11146 11880 11152 11892
rect 11107 11852 11152 11880
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 11514 11880 11520 11892
rect 11475 11852 11520 11880
rect 11514 11840 11520 11852
rect 11572 11840 11578 11892
rect 13354 11880 13360 11892
rect 13315 11852 13360 11880
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15289 11883 15347 11889
rect 15289 11880 15301 11883
rect 15252 11852 15301 11880
rect 15252 11840 15258 11852
rect 15289 11849 15301 11852
rect 15335 11849 15347 11883
rect 16666 11880 16672 11892
rect 16627 11852 16672 11880
rect 15289 11843 15347 11849
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 106 11772 112 11824
rect 164 11812 170 11824
rect 1581 11815 1639 11821
rect 1581 11812 1593 11815
rect 164 11784 1593 11812
rect 164 11772 170 11784
rect 1581 11781 1593 11784
rect 1627 11781 1639 11815
rect 1581 11775 1639 11781
rect 2682 11772 2688 11824
rect 2740 11812 2746 11824
rect 3605 11815 3663 11821
rect 3605 11812 3617 11815
rect 2740 11784 3617 11812
rect 2740 11772 2746 11784
rect 3605 11781 3617 11784
rect 3651 11781 3663 11815
rect 3605 11775 3663 11781
rect 4522 11772 4528 11824
rect 4580 11812 4586 11824
rect 6365 11815 6423 11821
rect 6365 11812 6377 11815
rect 4580 11784 6377 11812
rect 4580 11772 4586 11784
rect 6365 11781 6377 11784
rect 6411 11812 6423 11815
rect 6638 11812 6644 11824
rect 6411 11784 6644 11812
rect 6411 11781 6423 11784
rect 6365 11775 6423 11781
rect 6638 11772 6644 11784
rect 6696 11812 6702 11824
rect 8481 11815 8539 11821
rect 8481 11812 8493 11815
rect 6696 11784 8493 11812
rect 6696 11772 6702 11784
rect 3970 11744 3976 11756
rect 2240 11716 3976 11744
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 2240 11676 2268 11716
rect 3970 11704 3976 11716
rect 4028 11704 4034 11756
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 4126 11716 7205 11744
rect 1443 11648 2268 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 2682 11608 2688 11620
rect 2643 11580 2688 11608
rect 2682 11568 2688 11580
rect 2740 11568 2746 11620
rect 2777 11611 2835 11617
rect 2777 11577 2789 11611
rect 2823 11608 2835 11611
rect 3142 11608 3148 11620
rect 2823 11580 3148 11608
rect 2823 11577 2835 11580
rect 2777 11571 2835 11577
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 2792 11540 2820 11571
rect 3142 11568 3148 11580
rect 3200 11568 3206 11620
rect 3329 11611 3387 11617
rect 3329 11577 3341 11611
rect 3375 11608 3387 11611
rect 4126 11608 4154 11716
rect 7193 11713 7205 11716
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 5445 11679 5503 11685
rect 5445 11645 5457 11679
rect 5491 11645 5503 11679
rect 5626 11676 5632 11688
rect 5587 11648 5632 11676
rect 5445 11639 5503 11645
rect 3375 11580 4154 11608
rect 3375 11577 3387 11580
rect 3329 11571 3387 11577
rect 2547 11512 2820 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 2866 11500 2872 11552
rect 2924 11540 2930 11552
rect 3344 11540 3372 11571
rect 2924 11512 3372 11540
rect 2924 11500 2930 11512
rect 3510 11500 3516 11552
rect 3568 11540 3574 11552
rect 4157 11543 4215 11549
rect 4157 11540 4169 11543
rect 3568 11512 4169 11540
rect 3568 11500 3574 11512
rect 4157 11509 4169 11512
rect 4203 11509 4215 11543
rect 4157 11503 4215 11509
rect 5077 11543 5135 11549
rect 5077 11509 5089 11543
rect 5123 11540 5135 11543
rect 5460 11540 5488 11639
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 8312 11676 8340 11784
rect 8481 11781 8493 11784
rect 8527 11781 8539 11815
rect 8481 11775 8539 11781
rect 10226 11772 10232 11824
rect 10284 11821 10290 11824
rect 10284 11815 10333 11821
rect 10284 11781 10287 11815
rect 10321 11781 10333 11815
rect 11164 11812 11192 11840
rect 10284 11775 10333 11781
rect 10520 11784 11192 11812
rect 10284 11772 10290 11775
rect 8386 11704 8392 11756
rect 8444 11744 8450 11756
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 8444 11716 9321 11744
rect 8444 11704 8450 11716
rect 9309 11713 9321 11716
rect 9355 11744 9367 11747
rect 10134 11744 10140 11756
rect 9355 11716 10140 11744
rect 9355 11713 9367 11716
rect 9309 11707 9367 11713
rect 10134 11704 10140 11716
rect 10192 11744 10198 11756
rect 10520 11753 10548 11784
rect 12066 11772 12072 11824
rect 12124 11812 12130 11824
rect 13081 11815 13139 11821
rect 12124 11784 12801 11812
rect 12124 11772 12130 11784
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 10192 11716 10517 11744
rect 10192 11704 10198 11716
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 12667 11747 12725 11753
rect 12667 11744 12679 11747
rect 10836 11716 12679 11744
rect 10836 11704 10842 11716
rect 12667 11713 12679 11716
rect 12713 11713 12725 11747
rect 12773 11744 12801 11784
rect 13081 11781 13093 11815
rect 13127 11812 13139 11815
rect 13262 11812 13268 11824
rect 13127 11784 13268 11812
rect 13127 11781 13139 11784
rect 13081 11775 13139 11781
rect 13262 11772 13268 11784
rect 13320 11772 13326 11824
rect 16393 11815 16451 11821
rect 16393 11781 16405 11815
rect 16439 11812 16451 11815
rect 18414 11812 18420 11824
rect 16439 11784 18420 11812
rect 16439 11781 16451 11784
rect 16393 11775 16451 11781
rect 18414 11772 18420 11784
rect 18472 11772 18478 11824
rect 20806 11772 20812 11824
rect 20864 11812 20870 11824
rect 20947 11815 21005 11821
rect 20947 11812 20959 11815
rect 20864 11784 20959 11812
rect 20864 11772 20870 11784
rect 20947 11781 20959 11784
rect 20993 11812 21005 11815
rect 21637 11815 21695 11821
rect 21637 11812 21649 11815
rect 20993 11784 21649 11812
rect 20993 11781 21005 11784
rect 20947 11775 21005 11781
rect 21637 11781 21649 11784
rect 21683 11781 21695 11815
rect 21637 11775 21695 11781
rect 14921 11747 14979 11753
rect 14921 11744 14933 11747
rect 12773 11716 14933 11744
rect 12667 11707 12725 11713
rect 14921 11713 14933 11716
rect 14967 11744 14979 11747
rect 15197 11747 15255 11753
rect 15197 11744 15209 11747
rect 14967 11716 15209 11744
rect 14967 11713 14979 11716
rect 14921 11707 14979 11713
rect 15197 11713 15209 11716
rect 15243 11713 15255 11747
rect 18966 11744 18972 11756
rect 18927 11716 18972 11744
rect 15197 11707 15255 11713
rect 18966 11704 18972 11716
rect 19024 11744 19030 11756
rect 21269 11747 21327 11753
rect 21269 11744 21281 11747
rect 19024 11716 21281 11744
rect 19024 11704 19030 11716
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 8312 11648 8677 11676
rect 8665 11645 8677 11648
rect 8711 11676 8723 11679
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 8711 11648 9597 11676
rect 8711 11645 8723 11648
rect 8665 11639 8723 11645
rect 9585 11645 9597 11648
rect 9631 11676 9643 11679
rect 10410 11676 10416 11688
rect 9631 11648 10416 11676
rect 9631 11645 9643 11648
rect 9585 11639 9643 11645
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 12434 11676 12440 11688
rect 12395 11648 12440 11676
rect 12434 11636 12440 11648
rect 12492 11636 12498 11688
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11645 13967 11679
rect 13909 11639 13967 11645
rect 5902 11608 5908 11620
rect 5863 11580 5908 11608
rect 5902 11568 5908 11580
rect 5960 11568 5966 11620
rect 6917 11611 6975 11617
rect 6917 11577 6929 11611
rect 6963 11577 6975 11611
rect 6917 11571 6975 11577
rect 6086 11540 6092 11552
rect 5123 11512 6092 11540
rect 5123 11509 5135 11512
rect 5077 11503 5135 11509
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 6932 11540 6960 11571
rect 7006 11568 7012 11620
rect 7064 11608 7070 11620
rect 7374 11608 7380 11620
rect 7064 11580 7380 11608
rect 7064 11568 7070 11580
rect 7374 11568 7380 11580
rect 7432 11568 7438 11620
rect 9122 11608 9128 11620
rect 7806 11580 9128 11608
rect 7806 11540 7834 11580
rect 9122 11568 9128 11580
rect 9180 11568 9186 11620
rect 9490 11568 9496 11620
rect 9548 11608 9554 11620
rect 10137 11611 10195 11617
rect 10137 11608 10149 11611
rect 9548 11580 10149 11608
rect 9548 11568 9554 11580
rect 10137 11577 10149 11580
rect 10183 11608 10195 11611
rect 11885 11611 11943 11617
rect 11885 11608 11897 11611
rect 10183 11580 11897 11608
rect 10183 11577 10195 11580
rect 10137 11571 10195 11577
rect 11885 11577 11897 11580
rect 11931 11577 11943 11611
rect 11885 11571 11943 11577
rect 6932 11512 7834 11540
rect 8113 11543 8171 11549
rect 8113 11509 8125 11543
rect 8159 11540 8171 11543
rect 8294 11540 8300 11552
rect 8159 11512 8300 11540
rect 8159 11509 8171 11512
rect 8113 11503 8171 11509
rect 8294 11500 8300 11512
rect 8352 11540 8358 11552
rect 9674 11540 9680 11552
rect 8352 11512 9680 11540
rect 8352 11500 8358 11512
rect 9674 11500 9680 11512
rect 9732 11540 9738 11552
rect 9953 11543 10011 11549
rect 9953 11540 9965 11543
rect 9732 11512 9965 11540
rect 9732 11500 9738 11512
rect 9953 11509 9965 11512
rect 9999 11540 10011 11543
rect 10318 11540 10324 11552
rect 9999 11512 10324 11540
rect 9999 11509 10011 11512
rect 9953 11503 10011 11509
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 13446 11500 13452 11552
rect 13504 11540 13510 11552
rect 13725 11543 13783 11549
rect 13725 11540 13737 11543
rect 13504 11512 13737 11540
rect 13504 11500 13510 11512
rect 13725 11509 13737 11512
rect 13771 11540 13783 11543
rect 13924 11540 13952 11639
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 20859 11685 20887 11716
rect 21269 11713 21281 11716
rect 21315 11713 21327 11747
rect 21269 11707 21327 11713
rect 14369 11679 14427 11685
rect 14369 11676 14381 11679
rect 14056 11648 14381 11676
rect 14056 11636 14062 11648
rect 14369 11645 14381 11648
rect 14415 11645 14427 11679
rect 14369 11639 14427 11645
rect 14645 11679 14703 11685
rect 14645 11645 14657 11679
rect 14691 11676 14703 11679
rect 15473 11679 15531 11685
rect 15473 11676 15485 11679
rect 14691 11648 15485 11676
rect 14691 11645 14703 11648
rect 14645 11639 14703 11645
rect 15473 11645 15485 11648
rect 15519 11676 15531 11679
rect 17037 11679 17095 11685
rect 17037 11676 17049 11679
rect 15519 11648 17049 11676
rect 15519 11645 15531 11648
rect 15473 11639 15531 11645
rect 17037 11645 17049 11648
rect 17083 11645 17095 11679
rect 17037 11639 17095 11645
rect 20844 11679 20902 11685
rect 20844 11645 20856 11679
rect 20890 11645 20902 11679
rect 20844 11639 20902 11645
rect 15197 11611 15255 11617
rect 15197 11577 15209 11611
rect 15243 11608 15255 11611
rect 15794 11611 15852 11617
rect 15794 11608 15806 11611
rect 15243 11580 15806 11608
rect 15243 11577 15255 11580
rect 15197 11571 15255 11577
rect 15794 11577 15806 11580
rect 15840 11608 15852 11611
rect 15930 11608 15936 11620
rect 15840 11580 15936 11608
rect 15840 11577 15852 11580
rect 15794 11571 15852 11577
rect 15930 11568 15936 11580
rect 15988 11568 15994 11620
rect 18322 11608 18328 11620
rect 18283 11580 18328 11608
rect 18322 11568 18328 11580
rect 18380 11568 18386 11620
rect 18414 11568 18420 11620
rect 18472 11608 18478 11620
rect 18472 11580 18517 11608
rect 18472 11568 18478 11580
rect 18690 11568 18696 11620
rect 18748 11608 18754 11620
rect 19797 11611 19855 11617
rect 19797 11608 19809 11611
rect 18748 11580 19809 11608
rect 18748 11568 18754 11580
rect 19797 11577 19809 11580
rect 19843 11577 19855 11611
rect 19797 11571 19855 11577
rect 17678 11540 17684 11552
rect 13771 11512 13952 11540
rect 17639 11512 17684 11540
rect 13771 11509 13783 11512
rect 13725 11503 13783 11509
rect 17678 11500 17684 11512
rect 17736 11500 17742 11552
rect 19337 11543 19395 11549
rect 19337 11509 19349 11543
rect 19383 11540 19395 11543
rect 19426 11540 19432 11552
rect 19383 11512 19432 11540
rect 19383 11509 19395 11512
rect 19337 11503 19395 11509
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 1104 11450 22816 11472
rect 1104 11398 8982 11450
rect 9034 11398 9046 11450
rect 9098 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 16982 11450
rect 17034 11398 17046 11450
rect 17098 11398 17110 11450
rect 17162 11398 17174 11450
rect 17226 11398 22816 11450
rect 1104 11376 22816 11398
rect 1535 11339 1593 11345
rect 1535 11305 1547 11339
rect 1581 11336 1593 11339
rect 2682 11336 2688 11348
rect 1581 11308 2688 11336
rect 1581 11305 1593 11308
rect 1535 11299 1593 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 4985 11339 5043 11345
rect 4985 11336 4997 11339
rect 4764 11308 4997 11336
rect 4764 11296 4770 11308
rect 4985 11305 4997 11308
rect 5031 11305 5043 11339
rect 4985 11299 5043 11305
rect 6825 11339 6883 11345
rect 6825 11305 6837 11339
rect 6871 11336 6883 11339
rect 7006 11336 7012 11348
rect 6871 11308 7012 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 8205 11339 8263 11345
rect 8205 11305 8217 11339
rect 8251 11336 8263 11339
rect 8386 11336 8392 11348
rect 8251 11308 8392 11336
rect 8251 11305 8263 11308
rect 8205 11299 8263 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 10413 11339 10471 11345
rect 10413 11305 10425 11339
rect 10459 11336 10471 11339
rect 13998 11336 14004 11348
rect 10459 11308 14004 11336
rect 10459 11305 10471 11308
rect 10413 11299 10471 11305
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 15930 11336 15936 11348
rect 15891 11308 15936 11336
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 19426 11336 19432 11348
rect 19387 11308 19432 11336
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 1946 11268 1952 11280
rect 1907 11240 1952 11268
rect 1946 11228 1952 11240
rect 2004 11228 2010 11280
rect 2590 11268 2596 11280
rect 2551 11240 2596 11268
rect 2590 11228 2596 11240
rect 2648 11228 2654 11280
rect 5994 11228 6000 11280
rect 6052 11268 6058 11280
rect 6226 11271 6284 11277
rect 6226 11268 6238 11271
rect 6052 11240 6238 11268
rect 6052 11228 6058 11240
rect 6226 11237 6238 11240
rect 6272 11237 6284 11271
rect 6226 11231 6284 11237
rect 8110 11228 8116 11280
rect 8168 11268 8174 11280
rect 8481 11271 8539 11277
rect 8481 11268 8493 11271
rect 8168 11240 8493 11268
rect 8168 11228 8174 11240
rect 8481 11237 8493 11240
rect 8527 11268 8539 11271
rect 9398 11268 9404 11280
rect 8527 11240 9404 11268
rect 8527 11237 8539 11240
rect 8481 11231 8539 11237
rect 9398 11228 9404 11240
rect 9456 11268 9462 11280
rect 9456 11240 9959 11268
rect 9456 11228 9462 11240
rect 1461 11200 1467 11212
rect 1422 11172 1467 11200
rect 1461 11160 1467 11172
rect 1519 11160 1525 11212
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4341 11203 4399 11209
rect 4341 11200 4353 11203
rect 4212 11172 4353 11200
rect 4212 11160 4218 11172
rect 4341 11169 4353 11172
rect 4387 11169 4399 11203
rect 4341 11163 4399 11169
rect 4430 11160 4436 11212
rect 4488 11200 4494 11212
rect 5718 11200 5724 11212
rect 4488 11172 5724 11200
rect 4488 11160 4494 11172
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 7688 11203 7746 11209
rect 7688 11200 7700 11203
rect 7484 11172 7700 11200
rect 2130 11092 2136 11144
rect 2188 11132 2194 11144
rect 2501 11135 2559 11141
rect 2501 11132 2513 11135
rect 2188 11104 2513 11132
rect 2188 11092 2194 11104
rect 2501 11101 2513 11104
rect 2547 11132 2559 11135
rect 2774 11132 2780 11144
rect 2547 11104 2780 11132
rect 2547 11101 2559 11104
rect 2501 11095 2559 11101
rect 2774 11092 2780 11104
rect 2832 11092 2838 11144
rect 2958 11132 2964 11144
rect 2919 11104 2964 11132
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 5442 11132 5448 11144
rect 4755 11104 5448 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 5442 11092 5448 11104
rect 5500 11092 5506 11144
rect 5902 11132 5908 11144
rect 5815 11104 5908 11132
rect 5902 11092 5908 11104
rect 5960 11132 5966 11144
rect 7374 11132 7380 11144
rect 5960 11104 7380 11132
rect 5960 11092 5966 11104
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 2314 11024 2320 11076
rect 2372 11064 2378 11076
rect 7484 11073 7512 11172
rect 7688 11169 7700 11172
rect 7734 11169 7746 11203
rect 7688 11163 7746 11169
rect 9490 11160 9496 11212
rect 9548 11200 9554 11212
rect 9769 11203 9827 11209
rect 9769 11200 9781 11203
rect 9548 11172 9781 11200
rect 9548 11160 9554 11172
rect 9769 11169 9781 11172
rect 9815 11169 9827 11203
rect 9769 11163 9827 11169
rect 9931 11141 9959 11240
rect 10042 11228 10048 11280
rect 10100 11268 10106 11280
rect 10781 11271 10839 11277
rect 10781 11268 10793 11271
rect 10100 11240 10793 11268
rect 10100 11228 10106 11240
rect 10781 11237 10793 11240
rect 10827 11268 10839 11271
rect 11054 11268 11060 11280
rect 10827 11240 11060 11268
rect 10827 11237 10839 11240
rect 10781 11231 10839 11237
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 11514 11228 11520 11280
rect 11572 11268 11578 11280
rect 11695 11271 11753 11277
rect 11695 11268 11707 11271
rect 11572 11240 11707 11268
rect 11572 11228 11578 11240
rect 11695 11237 11707 11240
rect 11741 11268 11753 11271
rect 12066 11268 12072 11280
rect 11741 11240 12072 11268
rect 11741 11237 11753 11240
rect 11695 11231 11753 11237
rect 12066 11228 12072 11240
rect 12124 11228 12130 11280
rect 12250 11228 12256 11280
rect 12308 11268 12314 11280
rect 13265 11271 13323 11277
rect 13265 11268 13277 11271
rect 12308 11240 13277 11268
rect 12308 11228 12314 11240
rect 13265 11237 13277 11240
rect 13311 11268 13323 11271
rect 13538 11268 13544 11280
rect 13311 11240 13544 11268
rect 13311 11237 13323 11240
rect 13265 11231 13323 11237
rect 13538 11228 13544 11240
rect 13596 11228 13602 11280
rect 17402 11228 17408 11280
rect 17460 11268 17466 11280
rect 17773 11271 17831 11277
rect 17773 11268 17785 11271
rect 17460 11240 17785 11268
rect 17460 11228 17466 11240
rect 17773 11237 17785 11240
rect 17819 11237 17831 11271
rect 18322 11268 18328 11280
rect 18283 11240 18328 11268
rect 17773 11231 17831 11237
rect 18322 11228 18328 11240
rect 18380 11268 18386 11280
rect 18969 11271 19027 11277
rect 18969 11268 18981 11271
rect 18380 11240 18981 11268
rect 18380 11228 18386 11240
rect 18969 11237 18981 11240
rect 19015 11237 19027 11271
rect 18969 11231 19027 11237
rect 18414 11160 18420 11212
rect 18472 11200 18478 11212
rect 19150 11200 19156 11212
rect 18472 11172 19156 11200
rect 18472 11160 18478 11172
rect 19150 11160 19156 11172
rect 19208 11200 19214 11212
rect 19245 11203 19303 11209
rect 19245 11200 19257 11203
rect 19208 11172 19257 11200
rect 19208 11160 19214 11172
rect 19245 11169 19257 11172
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 20714 11160 20720 11212
rect 20772 11200 20778 11212
rect 20901 11203 20959 11209
rect 20901 11200 20913 11203
rect 20772 11172 20913 11200
rect 20772 11160 20778 11172
rect 20901 11169 20913 11172
rect 20947 11169 20959 11203
rect 20901 11163 20959 11169
rect 9916 11135 9974 11141
rect 9916 11101 9928 11135
rect 9962 11101 9974 11135
rect 10134 11132 10140 11144
rect 10095 11104 10140 11132
rect 9916 11095 9974 11101
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 11330 11132 11336 11144
rect 11291 11104 11336 11132
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 12710 11092 12716 11144
rect 12768 11132 12774 11144
rect 13173 11135 13231 11141
rect 13173 11132 13185 11135
rect 12768 11104 13185 11132
rect 12768 11092 12774 11104
rect 13173 11101 13185 11104
rect 13219 11132 13231 11135
rect 13262 11132 13268 11144
rect 13219 11104 13268 11132
rect 13219 11101 13231 11104
rect 13173 11095 13231 11101
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 13449 11135 13507 11141
rect 13449 11132 13461 11135
rect 13412 11104 13461 11132
rect 13412 11092 13418 11104
rect 13449 11101 13461 11104
rect 13495 11101 13507 11135
rect 15562 11132 15568 11144
rect 15523 11104 15568 11132
rect 13449 11095 13507 11101
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 17681 11135 17739 11141
rect 17681 11101 17693 11135
rect 17727 11132 17739 11135
rect 17862 11132 17868 11144
rect 17727 11104 17868 11132
rect 17727 11101 17739 11104
rect 17681 11095 17739 11101
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 7469 11067 7527 11073
rect 7469 11064 7481 11067
rect 2372 11036 7481 11064
rect 2372 11024 2378 11036
rect 7469 11033 7481 11036
rect 7515 11033 7527 11067
rect 7469 11027 7527 11033
rect 2222 10996 2228 11008
rect 2183 10968 2228 10996
rect 2222 10956 2228 10968
rect 2280 10956 2286 11008
rect 4522 11005 4528 11008
rect 4506 10999 4528 11005
rect 4506 10965 4518 10999
rect 4506 10959 4528 10965
rect 4522 10956 4528 10959
rect 4580 10956 4586 11008
rect 4617 10999 4675 11005
rect 4617 10965 4629 10999
rect 4663 10996 4675 10999
rect 4706 10996 4712 11008
rect 4663 10968 4712 10996
rect 4663 10965 4675 10968
rect 4617 10959 4675 10965
rect 4706 10956 4712 10968
rect 4764 10956 4770 11008
rect 5442 10996 5448 11008
rect 5403 10968 5448 10996
rect 5442 10956 5448 10968
rect 5500 10956 5506 11008
rect 7098 10996 7104 11008
rect 7059 10968 7104 10996
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 7791 10999 7849 11005
rect 7791 10996 7803 10999
rect 7248 10968 7803 10996
rect 7248 10956 7254 10968
rect 7791 10965 7803 10968
rect 7837 10965 7849 10999
rect 7791 10959 7849 10965
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 8849 10999 8907 11005
rect 8849 10996 8861 10999
rect 8352 10968 8861 10996
rect 8352 10956 8358 10968
rect 8849 10965 8861 10968
rect 8895 10965 8907 10999
rect 9490 10996 9496 11008
rect 9451 10968 9496 10996
rect 8849 10959 8907 10965
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 10045 10999 10103 11005
rect 10045 10996 10057 10999
rect 9732 10968 10057 10996
rect 9732 10956 9738 10968
rect 10045 10965 10057 10968
rect 10091 10965 10103 10999
rect 12250 10996 12256 11008
rect 12211 10968 12256 10996
rect 10045 10959 10103 10965
rect 12250 10956 12256 10968
rect 12308 10956 12314 11008
rect 12710 10996 12716 11008
rect 12671 10968 12716 10996
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 16485 10999 16543 11005
rect 16485 10965 16497 10999
rect 16531 10996 16543 10999
rect 17402 10996 17408 11008
rect 16531 10968 17408 10996
rect 16531 10965 16543 10968
rect 16485 10959 16543 10965
rect 17402 10956 17408 10968
rect 17460 10956 17466 11008
rect 21085 10999 21143 11005
rect 21085 10965 21097 10999
rect 21131 10996 21143 10999
rect 23566 10996 23572 11008
rect 21131 10968 23572 10996
rect 21131 10965 21143 10968
rect 21085 10959 21143 10965
rect 23566 10956 23572 10968
rect 23624 10956 23630 11008
rect 1104 10906 22816 10928
rect 1104 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 12982 10906
rect 13034 10854 13046 10906
rect 13098 10854 13110 10906
rect 13162 10854 13174 10906
rect 13226 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 22816 10906
rect 1104 10832 22816 10854
rect 1486 10752 1492 10804
rect 1544 10792 1550 10804
rect 1949 10795 2007 10801
rect 1949 10792 1961 10795
rect 1544 10764 1961 10792
rect 1544 10752 1550 10764
rect 1949 10761 1961 10764
rect 1995 10761 2007 10795
rect 1949 10755 2007 10761
rect 2406 10752 2412 10804
rect 2464 10792 2470 10804
rect 2961 10795 3019 10801
rect 2961 10792 2973 10795
rect 2464 10764 2973 10792
rect 2464 10752 2470 10764
rect 2961 10761 2973 10764
rect 3007 10792 3019 10795
rect 3418 10792 3424 10804
rect 3007 10764 3424 10792
rect 3007 10761 3019 10764
rect 2961 10755 3019 10761
rect 3418 10752 3424 10764
rect 3476 10752 3482 10804
rect 4338 10792 4344 10804
rect 4299 10764 4344 10792
rect 4338 10752 4344 10764
rect 4396 10792 4402 10804
rect 4706 10792 4712 10804
rect 4396 10764 4712 10792
rect 4396 10752 4402 10764
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 4893 10795 4951 10801
rect 4893 10761 4905 10795
rect 4939 10792 4951 10795
rect 5994 10792 6000 10804
rect 4939 10764 6000 10792
rect 4939 10761 4951 10764
rect 4893 10755 4951 10761
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7929 10795 7987 10801
rect 7929 10792 7941 10795
rect 7156 10764 7941 10792
rect 7156 10752 7162 10764
rect 7929 10761 7941 10764
rect 7975 10792 7987 10795
rect 9398 10792 9404 10804
rect 7975 10764 8708 10792
rect 9359 10764 9404 10792
rect 7975 10761 7987 10764
rect 7929 10755 7987 10761
rect 106 10684 112 10736
rect 164 10724 170 10736
rect 1581 10727 1639 10733
rect 1581 10724 1593 10727
rect 164 10696 1593 10724
rect 164 10684 170 10696
rect 1581 10693 1593 10696
rect 1627 10693 1639 10727
rect 1581 10687 1639 10693
rect 2501 10727 2559 10733
rect 2501 10693 2513 10727
rect 2547 10724 2559 10727
rect 2590 10724 2596 10736
rect 2547 10696 2596 10724
rect 2547 10693 2559 10696
rect 2501 10687 2559 10693
rect 2590 10684 2596 10696
rect 2648 10724 2654 10736
rect 2866 10724 2872 10736
rect 2648 10696 2872 10724
rect 2648 10684 2654 10696
rect 2866 10684 2872 10696
rect 2924 10724 2930 10736
rect 3973 10727 4031 10733
rect 3973 10724 3985 10727
rect 2924 10696 3985 10724
rect 2924 10684 2930 10696
rect 3973 10693 3985 10696
rect 4019 10693 4031 10727
rect 3973 10687 4031 10693
rect 4430 10684 4436 10736
rect 4488 10724 4494 10736
rect 5123 10727 5181 10733
rect 5123 10724 5135 10727
rect 4488 10696 5135 10724
rect 4488 10684 4494 10696
rect 5123 10693 5135 10696
rect 5169 10693 5181 10727
rect 5123 10687 5181 10693
rect 5261 10727 5319 10733
rect 5261 10693 5273 10727
rect 5307 10724 5319 10727
rect 5534 10724 5540 10736
rect 5307 10696 5540 10724
rect 5307 10693 5319 10696
rect 5261 10687 5319 10693
rect 5534 10684 5540 10696
rect 5592 10724 5598 10736
rect 7116 10724 7144 10752
rect 8570 10733 8576 10736
rect 5592 10696 7144 10724
rect 8554 10727 8576 10733
rect 5592 10684 5598 10696
rect 8554 10693 8566 10727
rect 8554 10687 8576 10693
rect 8570 10684 8576 10687
rect 8628 10684 8634 10736
rect 8680 10733 8708 10764
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 10134 10792 10140 10804
rect 10095 10764 10140 10792
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 11514 10792 11520 10804
rect 11475 10764 11520 10792
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 13538 10752 13544 10804
rect 13596 10792 13602 10804
rect 13633 10795 13691 10801
rect 13633 10792 13645 10795
rect 13596 10764 13645 10792
rect 13596 10752 13602 10764
rect 13633 10761 13645 10764
rect 13679 10761 13691 10795
rect 13633 10755 13691 10761
rect 15749 10795 15807 10801
rect 15749 10761 15761 10795
rect 15795 10792 15807 10795
rect 15930 10792 15936 10804
rect 15795 10764 15936 10792
rect 15795 10761 15807 10764
rect 15749 10755 15807 10761
rect 15930 10752 15936 10764
rect 15988 10752 15994 10804
rect 17402 10792 17408 10804
rect 17363 10764 17408 10792
rect 17402 10752 17408 10764
rect 17460 10752 17466 10804
rect 19150 10792 19156 10804
rect 19111 10764 19156 10792
rect 19150 10752 19156 10764
rect 19208 10752 19214 10804
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 20901 10795 20959 10801
rect 20901 10792 20913 10795
rect 20772 10764 20913 10792
rect 20772 10752 20778 10764
rect 20901 10761 20913 10764
rect 20947 10761 20959 10795
rect 20901 10755 20959 10761
rect 8665 10727 8723 10733
rect 8665 10693 8677 10727
rect 8711 10724 8723 10727
rect 10042 10724 10048 10736
rect 8711 10696 10048 10724
rect 8711 10693 8723 10696
rect 8665 10687 8723 10693
rect 10042 10684 10048 10696
rect 10100 10684 10106 10736
rect 4801 10659 4859 10665
rect 4801 10625 4813 10659
rect 4847 10656 4859 10659
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 4847 10628 5365 10656
rect 4847 10625 4859 10628
rect 4801 10619 4859 10625
rect 5353 10625 5365 10628
rect 5399 10656 5411 10659
rect 5442 10656 5448 10668
rect 5399 10628 5448 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 5442 10616 5448 10628
rect 5500 10656 5506 10668
rect 6362 10656 6368 10668
rect 5500 10628 6368 10656
rect 5500 10616 5506 10628
rect 6362 10616 6368 10628
rect 6420 10656 6426 10668
rect 8297 10659 8355 10665
rect 8297 10656 8309 10659
rect 6420 10628 8309 10656
rect 6420 10616 6426 10628
rect 8297 10625 8309 10628
rect 8343 10656 8355 10659
rect 8757 10659 8815 10665
rect 8757 10656 8769 10659
rect 8343 10628 8769 10656
rect 8343 10625 8355 10628
rect 8297 10619 8355 10625
rect 8757 10625 8769 10628
rect 8803 10656 8815 10659
rect 10152 10656 10180 10752
rect 17129 10727 17187 10733
rect 17129 10693 17141 10727
rect 17175 10724 17187 10727
rect 17862 10724 17868 10736
rect 17175 10696 17868 10724
rect 17175 10693 17187 10696
rect 17129 10687 17187 10693
rect 17862 10684 17868 10696
rect 17920 10684 17926 10736
rect 8803 10628 10180 10656
rect 11149 10659 11207 10665
rect 8803 10625 8815 10628
rect 8757 10619 8815 10625
rect 11149 10625 11161 10659
rect 11195 10656 11207 10659
rect 11330 10656 11336 10668
rect 11195 10628 11336 10656
rect 11195 10625 11207 10628
rect 11149 10619 11207 10625
rect 11330 10616 11336 10628
rect 11388 10656 11394 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11388 10628 11805 10656
rect 11388 10616 11394 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 12710 10656 12716 10668
rect 12671 10628 12716 10656
rect 11793 10619 11851 10625
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 13354 10656 13360 10668
rect 13315 10628 13360 10656
rect 13354 10616 13360 10628
rect 13412 10616 13418 10668
rect 14458 10616 14464 10668
rect 14516 10656 14522 10668
rect 14553 10659 14611 10665
rect 14553 10656 14565 10659
rect 14516 10628 14565 10656
rect 14516 10616 14522 10628
rect 14553 10625 14565 10628
rect 14599 10656 14611 10659
rect 15194 10656 15200 10668
rect 14599 10628 15200 10656
rect 14599 10625 14611 10628
rect 14553 10619 14611 10625
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1670 10588 1676 10600
rect 1443 10560 1676 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 1670 10548 1676 10560
rect 1728 10588 1734 10600
rect 2222 10588 2228 10600
rect 1728 10560 2228 10588
rect 1728 10548 1734 10560
rect 2222 10548 2228 10560
rect 2280 10548 2286 10600
rect 3050 10588 3056 10600
rect 3011 10560 3056 10588
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 3142 10548 3148 10600
rect 3200 10588 3206 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 3200 10560 6837 10588
rect 3200 10548 3206 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 7006 10588 7012 10600
rect 6967 10560 7012 10588
rect 6825 10551 6883 10557
rect 7006 10548 7012 10560
rect 7064 10548 7070 10600
rect 10502 10588 10508 10600
rect 10463 10560 10508 10588
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 10594 10548 10600 10600
rect 10652 10588 10658 10600
rect 14936 10597 14964 10628
rect 15194 10616 15200 10628
rect 15252 10616 15258 10668
rect 15381 10659 15439 10665
rect 15381 10625 15393 10659
rect 15427 10656 15439 10659
rect 15562 10656 15568 10668
rect 15427 10628 15568 10656
rect 15427 10625 15439 10628
rect 15381 10619 15439 10625
rect 15562 10616 15568 10628
rect 15620 10656 15626 10668
rect 16025 10659 16083 10665
rect 16025 10656 16037 10659
rect 15620 10628 16037 10656
rect 15620 10616 15626 10628
rect 16025 10625 16037 10628
rect 16071 10625 16083 10659
rect 16025 10619 16083 10625
rect 18322 10616 18328 10668
rect 18380 10656 18386 10668
rect 18417 10659 18475 10665
rect 18417 10656 18429 10659
rect 18380 10628 18429 10656
rect 18380 10616 18386 10628
rect 18417 10625 18429 10628
rect 18463 10625 18475 10659
rect 18417 10619 18475 10625
rect 10873 10591 10931 10597
rect 10873 10588 10885 10591
rect 10652 10560 10885 10588
rect 10652 10548 10658 10560
rect 10873 10557 10885 10560
rect 10919 10557 10931 10591
rect 10873 10551 10931 10557
rect 14921 10591 14979 10597
rect 14921 10557 14933 10591
rect 14967 10557 14979 10591
rect 15102 10588 15108 10600
rect 15063 10560 15108 10588
rect 14921 10551 14979 10557
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 4893 10523 4951 10529
rect 4893 10520 4905 10523
rect 4126 10492 4905 10520
rect 3418 10452 3424 10464
rect 3379 10424 3424 10452
rect 3418 10412 3424 10424
rect 3476 10452 3482 10464
rect 4126 10452 4154 10492
rect 4893 10489 4905 10492
rect 4939 10489 4951 10523
rect 4893 10483 4951 10489
rect 4982 10480 4988 10532
rect 5040 10520 5046 10532
rect 5442 10520 5448 10532
rect 5040 10492 5448 10520
rect 5040 10480 5046 10492
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 5718 10480 5724 10532
rect 5776 10520 5782 10532
rect 8386 10520 8392 10532
rect 5776 10492 8392 10520
rect 5776 10480 5782 10492
rect 8386 10480 8392 10492
rect 8444 10480 8450 10532
rect 12253 10523 12311 10529
rect 12253 10489 12265 10523
rect 12299 10520 12311 10523
rect 12526 10520 12532 10532
rect 12299 10492 12532 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 12526 10480 12532 10492
rect 12584 10520 12590 10532
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 12584 10492 12817 10520
rect 12584 10480 12590 10492
rect 12805 10489 12817 10492
rect 12851 10489 12863 10523
rect 18138 10520 18144 10532
rect 18099 10492 18144 10520
rect 12805 10483 12863 10489
rect 18138 10480 18144 10492
rect 18196 10480 18202 10532
rect 18233 10523 18291 10529
rect 18233 10489 18245 10523
rect 18279 10489 18291 10523
rect 18233 10483 18291 10489
rect 3476 10424 4154 10452
rect 3476 10412 3482 10424
rect 4798 10412 4804 10464
rect 4856 10452 4862 10464
rect 5626 10452 5632 10464
rect 4856 10424 5632 10452
rect 4856 10412 4862 10424
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 6178 10452 6184 10464
rect 6052 10424 6184 10452
rect 6052 10412 6058 10424
rect 6178 10412 6184 10424
rect 6236 10452 6242 10464
rect 6365 10455 6423 10461
rect 6365 10452 6377 10455
rect 6236 10424 6377 10452
rect 6236 10412 6242 10424
rect 6365 10421 6377 10424
rect 6411 10452 6423 10455
rect 8294 10452 8300 10464
rect 6411 10424 8300 10452
rect 6411 10421 6423 10424
rect 6365 10415 6423 10421
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8478 10412 8484 10464
rect 8536 10452 8542 10464
rect 9033 10455 9091 10461
rect 9033 10452 9045 10455
rect 8536 10424 9045 10452
rect 8536 10412 8542 10424
rect 9033 10421 9045 10424
rect 9079 10421 9091 10455
rect 9033 10415 9091 10421
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 9769 10455 9827 10461
rect 9769 10452 9781 10455
rect 9732 10424 9781 10452
rect 9732 10412 9738 10424
rect 9769 10421 9781 10424
rect 9815 10421 9827 10455
rect 17770 10452 17776 10464
rect 17731 10424 17776 10452
rect 9769 10415 9827 10421
rect 17770 10412 17776 10424
rect 17828 10452 17834 10464
rect 18248 10452 18276 10483
rect 17828 10424 18276 10452
rect 17828 10412 17834 10424
rect 1104 10362 22816 10384
rect 1104 10310 8982 10362
rect 9034 10310 9046 10362
rect 9098 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 16982 10362
rect 17034 10310 17046 10362
rect 17098 10310 17110 10362
rect 17162 10310 17174 10362
rect 17226 10310 22816 10362
rect 1104 10288 22816 10310
rect 1670 10248 1676 10260
rect 1631 10220 1676 10248
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 2130 10208 2136 10260
rect 2188 10248 2194 10260
rect 2225 10251 2283 10257
rect 2225 10248 2237 10251
rect 2188 10220 2237 10248
rect 2188 10208 2194 10220
rect 2225 10217 2237 10220
rect 2271 10217 2283 10251
rect 2225 10211 2283 10217
rect 2332 10220 3004 10248
rect 1464 10115 1522 10121
rect 1464 10081 1476 10115
rect 1510 10112 1522 10115
rect 2332 10112 2360 10220
rect 2976 10192 3004 10220
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 3421 10251 3479 10257
rect 3421 10248 3433 10251
rect 3108 10220 3433 10248
rect 3108 10208 3114 10220
rect 3421 10217 3433 10220
rect 3467 10248 3479 10251
rect 4525 10251 4583 10257
rect 4525 10248 4537 10251
rect 3467 10220 4537 10248
rect 3467 10217 3479 10220
rect 3421 10211 3479 10217
rect 4525 10217 4537 10220
rect 4571 10217 4583 10251
rect 4982 10248 4988 10260
rect 4525 10211 4583 10217
rect 4632 10220 4988 10248
rect 2590 10180 2596 10192
rect 2551 10152 2596 10180
rect 2590 10140 2596 10152
rect 2648 10140 2654 10192
rect 2958 10140 2964 10192
rect 3016 10180 3022 10192
rect 3145 10183 3203 10189
rect 3145 10180 3157 10183
rect 3016 10152 3157 10180
rect 3016 10140 3022 10152
rect 3145 10149 3157 10152
rect 3191 10149 3203 10183
rect 3145 10143 3203 10149
rect 4154 10140 4160 10192
rect 4212 10180 4218 10192
rect 4249 10183 4307 10189
rect 4249 10180 4261 10183
rect 4212 10152 4261 10180
rect 4212 10140 4218 10152
rect 4249 10149 4261 10152
rect 4295 10180 4307 10183
rect 4632 10180 4660 10220
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 5534 10248 5540 10260
rect 5495 10220 5540 10248
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 7006 10248 7012 10260
rect 6967 10220 7012 10248
rect 7006 10208 7012 10220
rect 7064 10208 7070 10260
rect 7374 10248 7380 10260
rect 7335 10220 7380 10248
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 9033 10251 9091 10257
rect 9033 10248 9045 10251
rect 8444 10220 9045 10248
rect 8444 10208 8450 10220
rect 9033 10217 9045 10220
rect 9079 10248 9091 10251
rect 9401 10251 9459 10257
rect 9401 10248 9413 10251
rect 9079 10220 9413 10248
rect 9079 10217 9091 10220
rect 9033 10211 9091 10217
rect 9401 10217 9413 10220
rect 9447 10248 9459 10251
rect 9490 10248 9496 10260
rect 9447 10220 9496 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 9953 10251 10011 10257
rect 9953 10217 9965 10251
rect 9999 10248 10011 10251
rect 10042 10248 10048 10260
rect 9999 10220 10048 10248
rect 9999 10217 10011 10220
rect 9953 10211 10011 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10594 10208 10600 10260
rect 10652 10248 10658 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 10652 10220 11069 10248
rect 10652 10208 10658 10220
rect 11057 10217 11069 10220
rect 11103 10217 11115 10251
rect 12526 10248 12532 10260
rect 12487 10220 12532 10248
rect 11057 10211 11115 10217
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 13262 10248 13268 10260
rect 13223 10220 13268 10248
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 14645 10251 14703 10257
rect 14645 10248 14657 10251
rect 14056 10220 14657 10248
rect 14056 10208 14062 10220
rect 14645 10217 14657 10220
rect 14691 10248 14703 10251
rect 15102 10248 15108 10260
rect 14691 10220 15108 10248
rect 14691 10217 14703 10220
rect 14645 10211 14703 10217
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 6546 10180 6552 10192
rect 4295 10152 4660 10180
rect 4724 10152 6552 10180
rect 4295 10149 4307 10152
rect 4249 10143 4307 10149
rect 1510 10084 2360 10112
rect 1510 10081 1522 10084
rect 1464 10075 1522 10081
rect 4338 10072 4344 10124
rect 4396 10112 4402 10124
rect 4724 10121 4752 10152
rect 6546 10140 6552 10152
rect 6604 10140 6610 10192
rect 6730 10180 6736 10192
rect 6691 10152 6736 10180
rect 6730 10140 6736 10152
rect 6788 10140 6794 10192
rect 6825 10183 6883 10189
rect 6825 10149 6837 10183
rect 6871 10180 6883 10183
rect 7929 10183 7987 10189
rect 7929 10180 7941 10183
rect 6871 10152 7941 10180
rect 6871 10149 6883 10152
rect 6825 10143 6883 10149
rect 7929 10149 7941 10152
rect 7975 10180 7987 10183
rect 8570 10180 8576 10192
rect 7975 10152 8576 10180
rect 7975 10149 7987 10152
rect 7929 10143 7987 10149
rect 8570 10140 8576 10152
rect 8628 10140 8634 10192
rect 17770 10180 17776 10192
rect 17731 10152 17776 10180
rect 17770 10140 17776 10152
rect 17828 10140 17834 10192
rect 4709 10115 4767 10121
rect 4709 10112 4721 10115
rect 4396 10084 4721 10112
rect 4396 10072 4402 10084
rect 4709 10081 4721 10084
rect 4755 10081 4767 10115
rect 4709 10075 4767 10081
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 4893 10115 4951 10121
rect 4893 10112 4905 10115
rect 4856 10084 4905 10112
rect 4856 10072 4862 10084
rect 4893 10081 4905 10084
rect 4939 10081 4951 10115
rect 4893 10075 4951 10081
rect 5718 10072 5724 10124
rect 5776 10112 5782 10124
rect 5997 10115 6055 10121
rect 5997 10112 6009 10115
rect 5776 10084 6009 10112
rect 5776 10072 5782 10084
rect 5997 10081 6009 10084
rect 6043 10081 6055 10115
rect 7190 10112 7196 10124
rect 5997 10075 6055 10081
rect 6159 10084 7196 10112
rect 2130 10004 2136 10056
rect 2188 10044 2194 10056
rect 2501 10047 2559 10053
rect 2501 10044 2513 10047
rect 2188 10016 2513 10044
rect 2188 10004 2194 10016
rect 2501 10013 2513 10016
rect 2547 10044 2559 10047
rect 3510 10044 3516 10056
rect 2547 10016 3516 10044
rect 2547 10013 2559 10016
rect 2501 10007 2559 10013
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 6159 10044 6187 10084
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 8294 10112 8300 10124
rect 8255 10084 8300 10112
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 8478 10112 8484 10124
rect 8439 10084 8484 10112
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 9769 10115 9827 10121
rect 9769 10112 9781 10115
rect 9732 10084 9781 10112
rect 9732 10072 9738 10084
rect 9769 10081 9781 10084
rect 9815 10081 9827 10115
rect 9769 10075 9827 10081
rect 12250 10072 12256 10124
rect 12308 10112 12314 10124
rect 12345 10115 12403 10121
rect 12345 10112 12357 10115
rect 12308 10084 12357 10112
rect 12308 10072 12314 10084
rect 12345 10081 12357 10084
rect 12391 10081 12403 10115
rect 12345 10075 12403 10081
rect 13354 10072 13360 10124
rect 13412 10112 13418 10124
rect 13814 10112 13820 10124
rect 13872 10121 13878 10124
rect 13872 10115 13910 10121
rect 13412 10084 13820 10112
rect 13412 10072 13418 10084
rect 13814 10072 13820 10084
rect 13898 10112 13910 10115
rect 17402 10112 17408 10124
rect 13898 10084 13965 10112
rect 17363 10084 17408 10112
rect 13898 10081 13910 10084
rect 13872 10075 13910 10081
rect 13872 10072 13878 10075
rect 17402 10072 17408 10084
rect 17460 10072 17466 10124
rect 6362 10044 6368 10056
rect 4126 10016 6187 10044
rect 6323 10016 6368 10044
rect 1394 9936 1400 9988
rect 1452 9976 1458 9988
rect 1949 9979 2007 9985
rect 1949 9976 1961 9979
rect 1452 9948 1961 9976
rect 1452 9936 1458 9948
rect 1949 9945 1961 9948
rect 1995 9976 2007 9979
rect 4126 9976 4154 10016
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 6546 10004 6552 10056
rect 6604 10044 6610 10056
rect 8312 10044 8340 10072
rect 8754 10044 8760 10056
rect 6604 10016 8340 10044
rect 8715 10016 8760 10044
rect 6604 10004 6610 10016
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 1995 9948 2452 9976
rect 1995 9945 2007 9948
rect 1949 9939 2007 9945
rect 2424 9908 2452 9948
rect 3160 9948 4154 9976
rect 6162 9979 6220 9985
rect 3160 9908 3188 9948
rect 6162 9945 6174 9979
rect 6208 9976 6220 9979
rect 6454 9976 6460 9988
rect 6208 9948 6460 9976
rect 6208 9945 6220 9948
rect 6162 9939 6220 9945
rect 6454 9936 6460 9948
rect 6512 9976 6518 9988
rect 6825 9979 6883 9985
rect 6825 9976 6837 9979
rect 6512 9948 6837 9976
rect 6512 9936 6518 9948
rect 6825 9945 6837 9948
rect 6871 9945 6883 9979
rect 9674 9976 9680 9988
rect 6825 9939 6883 9945
rect 7576 9948 9680 9976
rect 2424 9880 3188 9908
rect 3881 9911 3939 9917
rect 3881 9877 3893 9911
rect 3927 9908 3939 9911
rect 4154 9908 4160 9920
rect 3927 9880 4160 9908
rect 3927 9877 3939 9880
rect 3881 9871 3939 9877
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 5813 9911 5871 9917
rect 5813 9908 5825 9911
rect 5592 9880 5825 9908
rect 5592 9868 5598 9880
rect 5813 9877 5825 9880
rect 5859 9908 5871 9911
rect 5994 9908 6000 9920
rect 5859 9880 6000 9908
rect 5859 9877 5871 9880
rect 5813 9871 5871 9877
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 6270 9868 6276 9920
rect 6328 9908 6334 9920
rect 7576 9908 7604 9948
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 6328 9880 7604 9908
rect 6328 9868 6334 9880
rect 10502 9868 10508 9920
rect 10560 9908 10566 9920
rect 10781 9911 10839 9917
rect 10781 9908 10793 9911
rect 10560 9880 10793 9908
rect 10560 9868 10566 9880
rect 10781 9877 10793 9880
rect 10827 9908 10839 9911
rect 11698 9908 11704 9920
rect 10827 9880 11704 9908
rect 10827 9877 10839 9880
rect 10781 9871 10839 9877
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 13955 9911 14013 9917
rect 13955 9877 13967 9911
rect 14001 9908 14013 9911
rect 14090 9908 14096 9920
rect 14001 9880 14096 9908
rect 14001 9877 14013 9880
rect 13955 9871 14013 9877
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 18046 9908 18052 9920
rect 18007 9880 18052 9908
rect 18046 9868 18052 9880
rect 18104 9868 18110 9920
rect 1104 9818 22816 9840
rect 1104 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 12982 9818
rect 13034 9766 13046 9818
rect 13098 9766 13110 9818
rect 13162 9766 13174 9818
rect 13226 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 22816 9818
rect 1104 9744 22816 9766
rect 2130 9704 2136 9716
rect 2091 9676 2136 9704
rect 2130 9664 2136 9676
rect 2188 9664 2194 9716
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 4338 9704 4344 9716
rect 4120 9676 4344 9704
rect 4120 9664 4126 9676
rect 4338 9664 4344 9676
rect 4396 9704 4402 9716
rect 4433 9707 4491 9713
rect 4433 9704 4445 9707
rect 4396 9676 4445 9704
rect 4396 9664 4402 9676
rect 4433 9673 4445 9676
rect 4479 9673 4491 9707
rect 4798 9704 4804 9716
rect 4759 9676 4804 9704
rect 4433 9667 4491 9673
rect 4798 9664 4804 9676
rect 4856 9664 4862 9716
rect 6181 9707 6239 9713
rect 6181 9673 6193 9707
rect 6227 9704 6239 9707
rect 6270 9704 6276 9716
rect 6227 9676 6276 9704
rect 6227 9673 6239 9676
rect 6181 9667 6239 9673
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 6457 9707 6515 9713
rect 6457 9704 6469 9707
rect 6420 9676 6469 9704
rect 6420 9664 6426 9676
rect 6457 9673 6469 9676
rect 6503 9673 6515 9707
rect 6457 9667 6515 9673
rect 8294 9664 8300 9716
rect 8352 9704 8358 9716
rect 8481 9707 8539 9713
rect 8481 9704 8493 9707
rect 8352 9676 8493 9704
rect 8352 9664 8358 9676
rect 8481 9673 8493 9676
rect 8527 9704 8539 9707
rect 10502 9704 10508 9716
rect 8527 9676 10508 9704
rect 8527 9673 8539 9676
rect 8481 9667 8539 9673
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 12250 9664 12256 9716
rect 12308 9704 12314 9716
rect 12897 9707 12955 9713
rect 12897 9704 12909 9707
rect 12308 9676 12909 9704
rect 12308 9664 12314 9676
rect 12897 9673 12909 9676
rect 12943 9673 12955 9707
rect 12897 9667 12955 9673
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 16991 9707 17049 9713
rect 13872 9676 13917 9704
rect 13872 9664 13878 9676
rect 16991 9673 17003 9707
rect 17037 9704 17049 9707
rect 18046 9704 18052 9716
rect 17037 9676 18052 9704
rect 17037 9673 17049 9676
rect 16991 9667 17049 9673
rect 18046 9664 18052 9676
rect 18104 9664 18110 9716
rect 106 9596 112 9648
rect 164 9636 170 9648
rect 1581 9639 1639 9645
rect 1581 9636 1593 9639
rect 164 9608 1593 9636
rect 164 9596 170 9608
rect 1581 9605 1593 9608
rect 1627 9605 1639 9639
rect 8113 9639 8171 9645
rect 8113 9636 8125 9639
rect 1581 9599 1639 9605
rect 6012 9608 8125 9636
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2590 9568 2596 9580
rect 2547 9540 2596 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2590 9528 2596 9540
rect 2648 9568 2654 9580
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2648 9540 2697 9568
rect 2648 9528 2654 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 2866 9500 2872 9512
rect 2827 9472 2872 9500
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 4982 9460 4988 9512
rect 5040 9500 5046 9512
rect 5442 9500 5448 9512
rect 5040 9472 5448 9500
rect 5040 9460 5046 9472
rect 5442 9460 5448 9472
rect 5500 9500 5506 9512
rect 5721 9503 5779 9509
rect 5721 9500 5733 9503
rect 5500 9472 5733 9500
rect 5500 9460 5506 9472
rect 5721 9469 5733 9472
rect 5767 9500 5779 9503
rect 6012 9500 6040 9608
rect 8113 9605 8125 9608
rect 8159 9605 8171 9639
rect 8113 9599 8171 9605
rect 9950 9596 9956 9648
rect 10008 9636 10014 9648
rect 11514 9636 11520 9648
rect 10008 9608 11520 9636
rect 10008 9596 10014 9608
rect 11514 9596 11520 9608
rect 11572 9596 11578 9648
rect 17402 9596 17408 9648
rect 17460 9636 17466 9648
rect 17681 9639 17739 9645
rect 17681 9636 17693 9639
rect 17460 9608 17693 9636
rect 17460 9596 17466 9608
rect 17681 9605 17693 9608
rect 17727 9605 17739 9639
rect 17681 9599 17739 9605
rect 9401 9571 9459 9577
rect 9401 9537 9413 9571
rect 9447 9568 9459 9571
rect 10226 9568 10232 9580
rect 9447 9540 10232 9568
rect 9447 9537 9459 9540
rect 9401 9531 9459 9537
rect 10226 9528 10232 9540
rect 10284 9528 10290 9580
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9568 12495 9571
rect 12710 9568 12716 9580
rect 12483 9540 12716 9568
rect 12483 9537 12495 9540
rect 12437 9531 12495 9537
rect 12710 9528 12716 9540
rect 12768 9528 12774 9580
rect 7190 9500 7196 9512
rect 5767 9472 6040 9500
rect 7151 9472 7196 9500
rect 5767 9469 5779 9472
rect 5721 9463 5779 9469
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 9950 9500 9956 9512
rect 7570 9472 9956 9500
rect 4154 9392 4160 9444
rect 4212 9432 4218 9444
rect 4522 9432 4528 9444
rect 4212 9404 4528 9432
rect 4212 9392 4218 9404
rect 4522 9392 4528 9404
rect 4580 9432 4586 9444
rect 6454 9432 6460 9444
rect 4580 9404 6460 9432
rect 4580 9392 4586 9404
rect 6454 9392 6460 9404
rect 6512 9392 6518 9444
rect 7570 9441 7598 9472
rect 9950 9460 9956 9472
rect 10008 9460 10014 9512
rect 16920 9503 16978 9509
rect 16920 9469 16932 9503
rect 16966 9500 16978 9503
rect 16966 9472 17448 9500
rect 16966 9469 16978 9472
rect 16920 9463 16978 9469
rect 7101 9435 7159 9441
rect 7101 9401 7113 9435
rect 7147 9432 7159 9435
rect 7555 9435 7613 9441
rect 7555 9432 7567 9435
rect 7147 9404 7567 9432
rect 7147 9401 7159 9404
rect 7101 9395 7159 9401
rect 7555 9401 7567 9404
rect 7601 9401 7613 9435
rect 7555 9395 7613 9401
rect 7834 9392 7840 9444
rect 7892 9432 7898 9444
rect 8478 9432 8484 9444
rect 7892 9404 8484 9432
rect 7892 9392 7898 9404
rect 8478 9392 8484 9404
rect 8536 9432 8542 9444
rect 8757 9435 8815 9441
rect 8757 9432 8769 9435
rect 8536 9404 8769 9432
rect 8536 9392 8542 9404
rect 8757 9401 8769 9404
rect 8803 9401 8815 9435
rect 8757 9395 8815 9401
rect 10137 9435 10195 9441
rect 10137 9401 10149 9435
rect 10183 9401 10195 9435
rect 10137 9395 10195 9401
rect 5350 9364 5356 9376
rect 5311 9336 5356 9364
rect 5350 9324 5356 9336
rect 5408 9324 5414 9376
rect 9674 9364 9680 9376
rect 9635 9336 9680 9364
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 10152 9364 10180 9395
rect 10226 9392 10232 9444
rect 10284 9432 10290 9444
rect 10781 9435 10839 9441
rect 10284 9404 10329 9432
rect 10284 9392 10290 9404
rect 10781 9401 10793 9435
rect 10827 9432 10839 9435
rect 11146 9432 11152 9444
rect 10827 9404 11152 9432
rect 10827 9401 10839 9404
rect 10781 9395 10839 9401
rect 11146 9392 11152 9404
rect 11204 9392 11210 9444
rect 17420 9376 17448 9472
rect 11057 9367 11115 9373
rect 11057 9364 11069 9367
rect 9824 9336 11069 9364
rect 9824 9324 9830 9336
rect 11057 9333 11069 9336
rect 11103 9333 11115 9367
rect 17402 9364 17408 9376
rect 17363 9336 17408 9364
rect 11057 9327 11115 9333
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 1104 9274 22816 9296
rect 1104 9222 8982 9274
rect 9034 9222 9046 9274
rect 9098 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 16982 9274
rect 17034 9222 17046 9274
rect 17098 9222 17110 9274
rect 17162 9222 17174 9274
rect 17226 9222 22816 9274
rect 1104 9200 22816 9222
rect 2777 9163 2835 9169
rect 2777 9129 2789 9163
rect 2823 9160 2835 9163
rect 2866 9160 2872 9172
rect 2823 9132 2872 9160
rect 2823 9129 2835 9132
rect 2777 9123 2835 9129
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 3053 9163 3111 9169
rect 3053 9160 3065 9163
rect 3016 9132 3065 9160
rect 3016 9120 3022 9132
rect 3053 9129 3065 9132
rect 3099 9129 3111 9163
rect 3053 9123 3111 9129
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 4203 9163 4261 9169
rect 4203 9160 4215 9163
rect 3660 9132 4215 9160
rect 3660 9120 3666 9132
rect 4203 9129 4215 9132
rect 4249 9129 4261 9163
rect 4982 9160 4988 9172
rect 4943 9132 4988 9160
rect 4203 9123 4261 9129
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 6454 9160 6460 9172
rect 6415 9132 6460 9160
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 7190 9160 7196 9172
rect 7151 9132 7196 9160
rect 7190 9120 7196 9132
rect 7248 9160 7254 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 7248 9132 7481 9160
rect 7248 9120 7254 9132
rect 7469 9129 7481 9132
rect 7515 9129 7527 9163
rect 7469 9123 7527 9129
rect 9950 9120 9956 9172
rect 10008 9160 10014 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 10008 9132 10057 9160
rect 10008 9120 10014 9132
rect 10045 9129 10057 9132
rect 10091 9129 10103 9163
rect 10045 9123 10103 9129
rect 10226 9120 10232 9172
rect 10284 9160 10290 9172
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 10284 9132 10609 9160
rect 10284 9120 10290 9132
rect 10597 9129 10609 9132
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 3786 9052 3792 9104
rect 3844 9092 3850 9104
rect 5261 9095 5319 9101
rect 3844 9064 5028 9092
rect 3844 9052 3850 9064
rect 1946 9024 1952 9036
rect 1907 8996 1952 9024
rect 1946 8984 1952 8996
rect 2004 8984 2010 9036
rect 2222 8984 2228 9036
rect 2280 9024 2286 9036
rect 4132 9027 4190 9033
rect 4132 9024 4144 9027
rect 2280 8996 4144 9024
rect 2280 8984 2286 8996
rect 4132 8993 4144 8996
rect 4178 9024 4190 9027
rect 4525 9027 4583 9033
rect 4525 9024 4537 9027
rect 4178 8996 4537 9024
rect 4178 8993 4190 8996
rect 4132 8987 4190 8993
rect 4525 8993 4537 8996
rect 4571 8993 4583 9027
rect 4525 8987 4583 8993
rect 5000 8956 5028 9064
rect 5261 9061 5273 9095
rect 5307 9092 5319 9095
rect 5350 9092 5356 9104
rect 5307 9064 5356 9092
rect 5307 9061 5319 9064
rect 5261 9055 5319 9061
rect 5350 9052 5356 9064
rect 5408 9052 5414 9104
rect 5813 9095 5871 9101
rect 5813 9061 5825 9095
rect 5859 9092 5871 9095
rect 5902 9092 5908 9104
rect 5859 9064 5908 9092
rect 5859 9061 5871 9064
rect 5813 9055 5871 9061
rect 5902 9052 5908 9064
rect 5960 9092 5966 9104
rect 9766 9092 9772 9104
rect 5960 9064 9772 9092
rect 5960 9052 5966 9064
rect 9766 9052 9772 9064
rect 9824 9052 9830 9104
rect 6086 8984 6092 9036
rect 6144 9024 6150 9036
rect 7653 9027 7711 9033
rect 7653 9024 7665 9027
rect 6144 8996 7665 9024
rect 6144 8984 6150 8996
rect 7653 8993 7665 8996
rect 7699 8993 7711 9027
rect 7834 9024 7840 9036
rect 7795 8996 7840 9024
rect 7653 8987 7711 8993
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 5000 8928 5181 8956
rect 5169 8925 5181 8928
rect 5215 8956 5227 8959
rect 5626 8956 5632 8968
rect 5215 8928 5632 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 7668 8956 7696 8987
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 8754 8984 8760 9036
rect 8812 9024 8818 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 8812 8996 9689 9024
rect 8812 8984 8818 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 13722 9024 13728 9036
rect 13683 8996 13728 9024
rect 9677 8987 9735 8993
rect 13722 8984 13728 8996
rect 13780 9024 13786 9036
rect 14458 9024 14464 9036
rect 13780 8996 14464 9024
rect 13780 8984 13786 8996
rect 14458 8984 14464 8996
rect 14516 8984 14522 9036
rect 8110 8956 8116 8968
rect 7668 8928 8116 8956
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 13633 8959 13691 8965
rect 13633 8956 13645 8959
rect 13596 8928 13645 8956
rect 13596 8916 13602 8928
rect 13633 8925 13645 8928
rect 13679 8925 13691 8959
rect 13633 8919 13691 8925
rect 1762 8820 1768 8832
rect 1723 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 5718 8780 5724 8832
rect 5776 8820 5782 8832
rect 6089 8823 6147 8829
rect 6089 8820 6101 8823
rect 5776 8792 6101 8820
rect 5776 8780 5782 8792
rect 6089 8789 6101 8792
rect 6135 8789 6147 8823
rect 10870 8820 10876 8832
rect 10831 8792 10876 8820
rect 6089 8783 6147 8789
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 1104 8730 22816 8752
rect 1104 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 12982 8730
rect 13034 8678 13046 8730
rect 13098 8678 13110 8730
rect 13162 8678 13174 8730
rect 13226 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 22816 8730
rect 1104 8656 22816 8678
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5350 8616 5356 8628
rect 5123 8588 5356 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 6641 8619 6699 8625
rect 6641 8585 6653 8619
rect 6687 8616 6699 8619
rect 7834 8616 7840 8628
rect 6687 8588 7840 8616
rect 6687 8585 6699 8588
rect 6641 8579 6699 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8754 8576 8760 8628
rect 8812 8616 8818 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 8812 8588 9229 8616
rect 8812 8576 8818 8588
rect 9217 8585 9229 8588
rect 9263 8585 9275 8619
rect 9950 8616 9956 8628
rect 9911 8588 9956 8616
rect 9217 8579 9275 8585
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 2222 8480 2228 8492
rect 2183 8452 2228 8480
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 4062 8480 4068 8492
rect 3804 8452 4068 8480
rect 3804 8421 3832 8452
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 5261 8483 5319 8489
rect 5261 8480 5273 8483
rect 4764 8452 5273 8480
rect 4764 8440 4770 8452
rect 5261 8449 5273 8452
rect 5307 8449 5319 8483
rect 5902 8480 5908 8492
rect 5863 8452 5908 8480
rect 5261 8443 5319 8449
rect 5902 8440 5908 8452
rect 5960 8440 5966 8492
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 10505 8483 10563 8489
rect 10505 8480 10517 8483
rect 9447 8452 10517 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 10505 8449 10517 8452
rect 10551 8480 10563 8483
rect 10870 8480 10876 8492
rect 10551 8452 10876 8480
rect 10551 8449 10563 8452
rect 10505 8443 10563 8449
rect 10870 8440 10876 8452
rect 10928 8440 10934 8492
rect 3421 8415 3479 8421
rect 3421 8381 3433 8415
rect 3467 8412 3479 8415
rect 3789 8415 3847 8421
rect 3789 8412 3801 8415
rect 3467 8384 3801 8412
rect 3467 8381 3479 8384
rect 3421 8375 3479 8381
rect 3789 8381 3801 8384
rect 3835 8381 3847 8415
rect 3970 8412 3976 8424
rect 3931 8384 3976 8412
rect 3789 8375 3847 8381
rect 3970 8372 3976 8384
rect 4028 8372 4034 8424
rect 6273 8415 6331 8421
rect 6273 8381 6285 8415
rect 6319 8412 6331 8415
rect 7101 8415 7159 8421
rect 7101 8412 7113 8415
rect 6319 8384 7113 8412
rect 6319 8381 6331 8384
rect 6273 8375 6331 8381
rect 7101 8381 7113 8384
rect 7147 8412 7159 8415
rect 7742 8412 7748 8424
rect 7147 8384 7748 8412
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8313 1639 8347
rect 1581 8307 1639 8313
rect 1673 8347 1731 8353
rect 1673 8313 1685 8347
rect 1719 8344 1731 8347
rect 1762 8344 1768 8356
rect 1719 8316 1768 8344
rect 1719 8313 1731 8316
rect 1673 8307 1731 8313
rect 1596 8276 1624 8307
rect 1762 8304 1768 8316
rect 1820 8304 1826 8356
rect 5353 8347 5411 8353
rect 5353 8313 5365 8347
rect 5399 8344 5411 8347
rect 5442 8344 5448 8356
rect 5399 8316 5448 8344
rect 5399 8313 5411 8316
rect 5353 8307 5411 8313
rect 2590 8276 2596 8288
rect 1596 8248 2596 8276
rect 2590 8236 2596 8248
rect 2648 8236 2654 8288
rect 2866 8276 2872 8288
rect 2827 8248 2872 8276
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 3786 8276 3792 8288
rect 3747 8248 3792 8276
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 4709 8279 4767 8285
rect 4709 8245 4721 8279
rect 4755 8276 4767 8279
rect 5368 8276 5396 8307
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 10597 8347 10655 8353
rect 10597 8313 10609 8347
rect 10643 8313 10655 8347
rect 11146 8344 11152 8356
rect 11107 8316 11152 8344
rect 10597 8307 10655 8313
rect 7282 8276 7288 8288
rect 4755 8248 5396 8276
rect 7243 8248 7288 8276
rect 4755 8245 4767 8248
rect 4709 8239 4767 8245
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 8110 8276 8116 8288
rect 8071 8248 8116 8276
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 10318 8276 10324 8288
rect 10231 8248 10324 8276
rect 10318 8236 10324 8248
rect 10376 8276 10382 8288
rect 10612 8276 10640 8307
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 13722 8276 13728 8288
rect 10376 8248 10640 8276
rect 13683 8248 13728 8276
rect 10376 8236 10382 8248
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 1104 8186 22816 8208
rect 1104 8134 8982 8186
rect 9034 8134 9046 8186
rect 9098 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 16982 8186
rect 17034 8134 17046 8186
rect 17098 8134 17110 8186
rect 17162 8134 17174 8186
rect 17226 8134 22816 8186
rect 1104 8112 22816 8134
rect 1673 8075 1731 8081
rect 1673 8041 1685 8075
rect 1719 8072 1731 8075
rect 1762 8072 1768 8084
rect 1719 8044 1768 8072
rect 1719 8041 1731 8044
rect 1673 8035 1731 8041
rect 1762 8032 1768 8044
rect 1820 8032 1826 8084
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 1964 8044 2789 8072
rect 1964 8016 1992 8044
rect 2777 8041 2789 8044
rect 2823 8072 2835 8075
rect 2866 8072 2872 8084
rect 2823 8044 2872 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 3605 8075 3663 8081
rect 3605 8041 3617 8075
rect 3651 8072 3663 8075
rect 3970 8072 3976 8084
rect 3651 8044 3976 8072
rect 3651 8041 3663 8044
rect 3605 8035 3663 8041
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 4985 8075 5043 8081
rect 4985 8072 4997 8075
rect 4126 8044 4997 8072
rect 1946 8004 1952 8016
rect 1907 7976 1952 8004
rect 1946 7964 1952 7976
rect 2004 7964 2010 8016
rect 2222 7964 2228 8016
rect 2280 8004 2286 8016
rect 2501 8007 2559 8013
rect 2501 8004 2513 8007
rect 2280 7976 2513 8004
rect 2280 7964 2286 7976
rect 2501 7973 2513 7976
rect 2547 7973 2559 8007
rect 2884 8004 2912 8032
rect 4126 8004 4154 8044
rect 4985 8041 4997 8044
rect 5031 8041 5043 8075
rect 5626 8072 5632 8084
rect 5587 8044 5632 8072
rect 4985 8035 5043 8041
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 10318 8072 10324 8084
rect 10279 8044 10324 8072
rect 10318 8032 10324 8044
rect 10376 8032 10382 8084
rect 4338 8004 4344 8016
rect 2884 7976 4154 8004
rect 4299 7976 4344 8004
rect 2501 7967 2559 7973
rect 4338 7964 4344 7976
rect 4396 7964 4402 8016
rect 7282 8004 7288 8016
rect 7243 7976 7288 8004
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 11146 7964 11152 8016
rect 11204 8004 11210 8016
rect 11204 7976 19323 8004
rect 11204 7964 11210 7976
rect 19295 7948 19323 7976
rect 3786 7896 3792 7948
rect 3844 7936 3850 7948
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 3844 7908 4077 7936
rect 3844 7896 3850 7908
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 10226 7936 10232 7948
rect 10187 7908 10232 7936
rect 4065 7899 4123 7905
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7905 11943 7939
rect 12066 7936 12072 7948
rect 12027 7908 12072 7936
rect 11885 7899 11943 7905
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7868 1915 7871
rect 2130 7868 2136 7880
rect 1903 7840 2136 7868
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 2130 7828 2136 7840
rect 2188 7868 2194 7880
rect 3145 7871 3203 7877
rect 3145 7868 3157 7871
rect 2188 7840 3157 7868
rect 2188 7828 2194 7840
rect 3145 7837 3157 7840
rect 3191 7837 3203 7871
rect 3145 7831 3203 7837
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7868 6147 7871
rect 6270 7868 6276 7880
rect 6135 7840 6276 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 6270 7828 6276 7840
rect 6328 7868 6334 7880
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 6328 7840 7205 7868
rect 6328 7828 6334 7840
rect 7193 7837 7205 7840
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7868 7895 7871
rect 8202 7868 8208 7880
rect 7883 7840 8208 7868
rect 7883 7837 7895 7840
rect 7837 7831 7895 7837
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 11698 7828 11704 7880
rect 11756 7868 11762 7880
rect 11900 7868 11928 7899
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 19242 7936 19248 7948
rect 19300 7945 19323 7948
rect 19300 7939 19338 7945
rect 19190 7908 19248 7936
rect 19242 7896 19248 7908
rect 19326 7905 19338 7939
rect 19300 7899 19338 7905
rect 19300 7896 19306 7899
rect 12342 7868 12348 7880
rect 11756 7840 12112 7868
rect 12303 7840 12348 7868
rect 11756 7828 11762 7840
rect 1302 7760 1308 7812
rect 1360 7800 1366 7812
rect 5718 7800 5724 7812
rect 1360 7772 5724 7800
rect 1360 7760 1366 7772
rect 5718 7760 5724 7772
rect 5776 7760 5782 7812
rect 12084 7800 12112 7840
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 13538 7800 13544 7812
rect 12084 7772 13544 7800
rect 13538 7760 13544 7772
rect 13596 7760 13602 7812
rect 3970 7692 3976 7744
rect 4028 7732 4034 7744
rect 4522 7732 4528 7744
rect 4028 7704 4528 7732
rect 4028 7692 4034 7704
rect 4522 7692 4528 7704
rect 4580 7692 4586 7744
rect 4706 7692 4712 7744
rect 4764 7732 4770 7744
rect 5261 7735 5319 7741
rect 5261 7732 5273 7735
rect 4764 7704 5273 7732
rect 4764 7692 4770 7704
rect 5261 7701 5273 7704
rect 5307 7701 5319 7735
rect 6822 7732 6828 7744
rect 6783 7704 6828 7732
rect 5261 7695 5319 7701
rect 6822 7692 6828 7704
rect 6880 7692 6886 7744
rect 8665 7735 8723 7741
rect 8665 7701 8677 7735
rect 8711 7732 8723 7735
rect 8754 7732 8760 7744
rect 8711 7704 8760 7732
rect 8711 7701 8723 7704
rect 8665 7695 8723 7701
rect 8754 7692 8760 7704
rect 8812 7692 8818 7744
rect 12710 7692 12716 7744
rect 12768 7732 12774 7744
rect 12897 7735 12955 7741
rect 12897 7732 12909 7735
rect 12768 7704 12909 7732
rect 12768 7692 12774 7704
rect 12897 7701 12909 7704
rect 12943 7701 12955 7735
rect 12897 7695 12955 7701
rect 19383 7735 19441 7741
rect 19383 7701 19395 7735
rect 19429 7732 19441 7735
rect 19978 7732 19984 7744
rect 19429 7704 19984 7732
rect 19429 7701 19441 7704
rect 19383 7695 19441 7701
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 1104 7642 22816 7664
rect 1104 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 12982 7642
rect 13034 7590 13046 7642
rect 13098 7590 13110 7642
rect 13162 7590 13174 7642
rect 13226 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 22816 7642
rect 1104 7568 22816 7590
rect 106 7488 112 7540
rect 164 7528 170 7540
rect 2869 7531 2927 7537
rect 2869 7528 2881 7531
rect 164 7500 2881 7528
rect 164 7488 170 7500
rect 2869 7497 2881 7500
rect 2915 7497 2927 7531
rect 2869 7491 2927 7497
rect 4065 7531 4123 7537
rect 4065 7497 4077 7531
rect 4111 7528 4123 7531
rect 4111 7500 4476 7528
rect 4111 7497 4123 7500
rect 4065 7491 4123 7497
rect 2130 7460 2136 7472
rect 2091 7432 2136 7460
rect 2130 7420 2136 7432
rect 2188 7420 2194 7472
rect 2884 7324 2912 7491
rect 3878 7420 3884 7472
rect 3936 7460 3942 7472
rect 4448 7469 4476 7500
rect 5718 7488 5724 7540
rect 5776 7528 5782 7540
rect 5859 7531 5917 7537
rect 5859 7528 5871 7531
rect 5776 7500 5871 7528
rect 5776 7488 5782 7500
rect 5859 7497 5871 7500
rect 5905 7497 5917 7531
rect 6270 7528 6276 7540
rect 6231 7500 6276 7528
rect 5859 7491 5917 7497
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 7742 7528 7748 7540
rect 7703 7500 7748 7528
rect 7742 7488 7748 7500
rect 7800 7528 7806 7540
rect 8018 7528 8024 7540
rect 7800 7500 8024 7528
rect 7800 7488 7806 7500
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 10045 7531 10103 7537
rect 10045 7497 10057 7531
rect 10091 7528 10103 7531
rect 10226 7528 10232 7540
rect 10091 7500 10232 7528
rect 10091 7497 10103 7500
rect 10045 7491 10103 7497
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 11698 7528 11704 7540
rect 11659 7500 11704 7528
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 12066 7528 12072 7540
rect 12027 7500 12072 7528
rect 12066 7488 12072 7500
rect 12124 7488 12130 7540
rect 14550 7488 14556 7540
rect 14608 7528 14614 7540
rect 14737 7531 14795 7537
rect 14737 7528 14749 7531
rect 14608 7500 14749 7528
rect 14608 7488 14614 7500
rect 14737 7497 14749 7500
rect 14783 7497 14795 7531
rect 19242 7528 19248 7540
rect 19203 7500 19248 7528
rect 14737 7491 14795 7497
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 21450 7528 21456 7540
rect 21411 7500 21456 7528
rect 21450 7488 21456 7500
rect 21508 7488 21514 7540
rect 4295 7463 4353 7469
rect 4295 7460 4307 7463
rect 3936 7432 4307 7460
rect 3936 7420 3942 7432
rect 4295 7429 4307 7432
rect 4341 7429 4353 7463
rect 4295 7423 4353 7429
rect 4433 7463 4491 7469
rect 4433 7429 4445 7463
rect 4479 7460 4491 7463
rect 4798 7460 4804 7472
rect 4479 7432 4804 7460
rect 4479 7429 4491 7432
rect 4433 7423 4491 7429
rect 4798 7420 4804 7432
rect 4856 7460 4862 7472
rect 6178 7460 6184 7472
rect 4856 7432 6184 7460
rect 4856 7420 4862 7432
rect 6178 7420 6184 7432
rect 6236 7420 6242 7472
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4525 7395 4583 7401
rect 4525 7392 4537 7395
rect 4028 7364 4537 7392
rect 4028 7352 4034 7364
rect 4525 7361 4537 7364
rect 4571 7392 4583 7395
rect 4614 7392 4620 7404
rect 4571 7364 4620 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 8665 7395 8723 7401
rect 8665 7361 8677 7395
rect 8711 7392 8723 7395
rect 8754 7392 8760 7404
rect 8711 7364 8760 7392
rect 8711 7361 8723 7364
rect 8665 7355 8723 7361
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 13446 7392 13452 7404
rect 13407 7364 13452 7392
rect 13446 7352 13452 7364
rect 13504 7392 13510 7404
rect 13504 7364 13814 7392
rect 13504 7352 13510 7364
rect 3088 7327 3146 7333
rect 3088 7324 3100 7327
rect 2884 7296 3100 7324
rect 3088 7293 3100 7296
rect 3134 7293 3146 7327
rect 3088 7287 3146 7293
rect 5788 7327 5846 7333
rect 5788 7293 5800 7327
rect 5834 7324 5846 7327
rect 5994 7324 6000 7336
rect 5834 7296 6000 7324
rect 5834 7293 5846 7296
rect 5788 7287 5846 7293
rect 5994 7284 6000 7296
rect 6052 7284 6058 7336
rect 6822 7324 6828 7336
rect 6783 7296 6828 7324
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 9677 7327 9735 7333
rect 9677 7293 9689 7327
rect 9723 7324 9735 7327
rect 9858 7324 9864 7336
rect 9723 7296 9864 7324
rect 9723 7293 9735 7296
rect 9677 7287 9735 7293
rect 9858 7284 9864 7296
rect 9916 7324 9922 7336
rect 10229 7327 10287 7333
rect 10229 7324 10241 7327
rect 9916 7296 10241 7324
rect 9916 7284 9922 7296
rect 10229 7293 10241 7296
rect 10275 7293 10287 7327
rect 13786 7324 13814 7364
rect 14528 7327 14586 7333
rect 14528 7324 14540 7327
rect 13786 7296 14540 7324
rect 10229 7287 10287 7293
rect 14528 7293 14540 7296
rect 14574 7324 14586 7327
rect 14921 7327 14979 7333
rect 14921 7324 14933 7327
rect 14574 7296 14933 7324
rect 14574 7293 14586 7296
rect 14528 7287 14586 7293
rect 14921 7293 14933 7296
rect 14967 7293 14979 7327
rect 14921 7287 14979 7293
rect 20968 7327 21026 7333
rect 20968 7293 20980 7327
rect 21014 7324 21026 7327
rect 21450 7324 21456 7336
rect 21014 7296 21456 7324
rect 21014 7293 21026 7296
rect 20968 7287 21026 7293
rect 21450 7284 21456 7296
rect 21508 7284 21514 7336
rect 1578 7256 1584 7268
rect 1539 7228 1584 7256
rect 1578 7216 1584 7228
rect 1636 7216 1642 7268
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7256 1731 7259
rect 4154 7256 4160 7268
rect 1719 7228 2544 7256
rect 4115 7228 4160 7256
rect 1719 7225 1731 7228
rect 1673 7219 1731 7225
rect 2516 7200 2544 7228
rect 4154 7216 4160 7228
rect 4212 7216 4218 7268
rect 4430 7216 4436 7268
rect 4488 7256 4494 7268
rect 4614 7256 4620 7268
rect 4488 7228 4620 7256
rect 4488 7216 4494 7228
rect 4614 7216 4620 7228
rect 4672 7216 4678 7268
rect 6549 7259 6607 7265
rect 6549 7256 6561 7259
rect 5460 7228 6561 7256
rect 2498 7188 2504 7200
rect 2459 7160 2504 7188
rect 2498 7148 2504 7160
rect 2556 7148 2562 7200
rect 2866 7148 2872 7200
rect 2924 7188 2930 7200
rect 3191 7191 3249 7197
rect 3191 7188 3203 7191
rect 2924 7160 3203 7188
rect 2924 7148 2930 7160
rect 3191 7157 3203 7160
rect 3237 7157 3249 7191
rect 3191 7151 3249 7157
rect 3697 7191 3755 7197
rect 3697 7157 3709 7191
rect 3743 7188 3755 7191
rect 3970 7188 3976 7200
rect 3743 7160 3976 7188
rect 3743 7157 3755 7160
rect 3697 7151 3755 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 4801 7191 4859 7197
rect 4801 7188 4813 7191
rect 4580 7160 4813 7188
rect 4580 7148 4586 7160
rect 4801 7157 4813 7160
rect 4847 7157 4859 7191
rect 5166 7188 5172 7200
rect 5127 7160 5172 7188
rect 4801 7151 4859 7157
rect 5166 7148 5172 7160
rect 5224 7188 5230 7200
rect 5460 7188 5488 7228
rect 6549 7225 6561 7228
rect 6595 7256 6607 7259
rect 7146 7259 7204 7265
rect 7146 7256 7158 7259
rect 6595 7228 7158 7256
rect 6595 7225 6607 7228
rect 6549 7219 6607 7225
rect 7146 7225 7158 7228
rect 7192 7225 7204 7259
rect 7146 7219 7204 7225
rect 8757 7259 8815 7265
rect 8757 7225 8769 7259
rect 8803 7225 8815 7259
rect 9306 7256 9312 7268
rect 9267 7228 9312 7256
rect 8757 7219 8815 7225
rect 5626 7188 5632 7200
rect 5224 7160 5488 7188
rect 5587 7160 5632 7188
rect 5224 7148 5230 7160
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 8481 7191 8539 7197
rect 8481 7157 8493 7191
rect 8527 7188 8539 7191
rect 8772 7188 8800 7219
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 10137 7259 10195 7265
rect 10137 7256 10149 7259
rect 9416 7228 10149 7256
rect 9416 7188 9444 7228
rect 10137 7225 10149 7228
rect 10183 7225 10195 7259
rect 10137 7219 10195 7225
rect 11698 7216 11704 7268
rect 11756 7256 11762 7268
rect 12710 7256 12716 7268
rect 11756 7228 12716 7256
rect 11756 7216 11762 7228
rect 12710 7216 12716 7228
rect 12768 7256 12774 7268
rect 12989 7259 13047 7265
rect 12989 7256 13001 7259
rect 12768 7228 13001 7256
rect 12768 7216 12774 7228
rect 12989 7225 13001 7228
rect 13035 7225 13047 7259
rect 12989 7219 13047 7225
rect 13081 7259 13139 7265
rect 13081 7225 13093 7259
rect 13127 7225 13139 7259
rect 13081 7219 13139 7225
rect 12802 7188 12808 7200
rect 8527 7160 9444 7188
rect 12763 7160 12808 7188
rect 8527 7157 8539 7160
rect 8481 7151 8539 7157
rect 12802 7148 12808 7160
rect 12860 7188 12866 7200
rect 13096 7188 13124 7219
rect 12860 7160 13124 7188
rect 12860 7148 12866 7160
rect 17310 7148 17316 7200
rect 17368 7188 17374 7200
rect 21039 7191 21097 7197
rect 21039 7188 21051 7191
rect 17368 7160 21051 7188
rect 17368 7148 17374 7160
rect 21039 7157 21051 7160
rect 21085 7157 21097 7191
rect 21039 7151 21097 7157
rect 1104 7098 22816 7120
rect 1104 7046 8982 7098
rect 9034 7046 9046 7098
rect 9098 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 17174 7098
rect 17226 7046 22816 7098
rect 1104 7024 22816 7046
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 2866 6984 2872 6996
rect 1636 6956 2872 6984
rect 1636 6944 1642 6956
rect 2866 6944 2872 6956
rect 2924 6944 2930 6996
rect 3513 6987 3571 6993
rect 3513 6953 3525 6987
rect 3559 6984 3571 6987
rect 3786 6984 3792 6996
rect 3559 6956 3792 6984
rect 3559 6953 3571 6956
rect 3513 6947 3571 6953
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 4157 6987 4215 6993
rect 4157 6953 4169 6987
rect 4203 6953 4215 6987
rect 6086 6984 6092 6996
rect 4157 6947 4215 6953
rect 5000 6956 6092 6984
rect 1926 6919 1984 6925
rect 1926 6885 1938 6919
rect 1972 6916 1984 6919
rect 2038 6916 2044 6928
rect 1972 6888 2044 6916
rect 1972 6885 1984 6888
rect 1926 6879 1984 6885
rect 2038 6876 2044 6888
rect 2096 6876 2102 6928
rect 4172 6916 4200 6947
rect 5000 6916 5028 6956
rect 6086 6944 6092 6956
rect 6144 6944 6150 6996
rect 6822 6984 6828 6996
rect 6783 6956 6828 6984
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 7282 6984 7288 6996
rect 7243 6956 7288 6984
rect 7282 6944 7288 6956
rect 7340 6944 7346 6996
rect 9306 6984 9312 6996
rect 7944 6956 9312 6984
rect 2700 6888 4200 6916
rect 4356 6888 5028 6916
rect 5813 6919 5871 6925
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 2406 6848 2412 6860
rect 1719 6820 2412 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 2406 6808 2412 6820
rect 2464 6848 2470 6860
rect 2700 6848 2728 6888
rect 2464 6820 2728 6848
rect 2464 6808 2470 6820
rect 3786 6808 3792 6860
rect 3844 6848 3850 6860
rect 4356 6857 4384 6888
rect 5813 6885 5825 6919
rect 5859 6916 5871 6919
rect 5994 6916 6000 6928
rect 5859 6888 6000 6916
rect 5859 6885 5871 6888
rect 5813 6879 5871 6885
rect 5994 6876 6000 6888
rect 6052 6916 6058 6928
rect 7944 6925 7972 6956
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 11698 6984 11704 6996
rect 11659 6956 11704 6984
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 12437 6987 12495 6993
rect 12437 6984 12449 6987
rect 12400 6956 12449 6984
rect 12400 6944 12406 6956
rect 12437 6953 12449 6956
rect 12483 6953 12495 6987
rect 12437 6947 12495 6953
rect 7929 6919 7987 6925
rect 6052 6888 7052 6916
rect 6052 6876 6058 6888
rect 4341 6851 4399 6857
rect 4341 6848 4353 6851
rect 3844 6820 4353 6848
rect 3844 6808 3850 6820
rect 4341 6817 4353 6820
rect 4387 6817 4399 6851
rect 4522 6848 4528 6860
rect 4483 6820 4528 6848
rect 4341 6811 4399 6817
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 6178 6848 6184 6860
rect 6139 6820 6184 6848
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6733 6851 6791 6857
rect 6733 6817 6745 6851
rect 6779 6817 6791 6851
rect 6914 6848 6920 6860
rect 6875 6820 6920 6848
rect 6733 6811 6791 6817
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 6362 6780 6368 6792
rect 4212 6752 6368 6780
rect 4212 6740 4218 6752
rect 6362 6740 6368 6752
rect 6420 6780 6426 6792
rect 6748 6780 6776 6811
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 6420 6752 6776 6780
rect 6420 6740 6426 6752
rect 2038 6672 2044 6724
rect 2096 6712 2102 6724
rect 4338 6712 4344 6724
rect 2096 6684 4344 6712
rect 2096 6672 2102 6684
rect 4338 6672 4344 6684
rect 4396 6712 4402 6724
rect 5166 6712 5172 6724
rect 4396 6684 5172 6712
rect 4396 6672 4402 6684
rect 5166 6672 5172 6684
rect 5224 6672 5230 6724
rect 7024 6712 7052 6888
rect 7929 6885 7941 6919
rect 7975 6885 7987 6919
rect 7929 6879 7987 6885
rect 8018 6876 8024 6928
rect 8076 6916 8082 6928
rect 9858 6916 9864 6928
rect 8076 6888 8121 6916
rect 9819 6888 9864 6916
rect 8076 6876 8082 6888
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 12250 6876 12256 6928
rect 12308 6916 12314 6928
rect 12897 6919 12955 6925
rect 12897 6916 12909 6919
rect 12308 6888 12909 6916
rect 12308 6876 12314 6888
rect 12897 6885 12909 6888
rect 12943 6885 12955 6919
rect 13446 6916 13452 6928
rect 13407 6888 13452 6916
rect 12897 6879 12955 6885
rect 13446 6876 13452 6888
rect 13504 6876 13510 6928
rect 8202 6780 8208 6792
rect 8163 6752 8208 6780
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6780 9827 6783
rect 11238 6780 11244 6792
rect 9815 6752 11244 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6749 12863 6783
rect 12805 6743 12863 6749
rect 8220 6712 8248 6740
rect 7024 6684 8248 6712
rect 9306 6672 9312 6724
rect 9364 6712 9370 6724
rect 10321 6715 10379 6721
rect 10321 6712 10333 6715
rect 9364 6684 10333 6712
rect 9364 6672 9370 6684
rect 10321 6681 10333 6684
rect 10367 6681 10379 6715
rect 10321 6675 10379 6681
rect 12710 6672 12716 6724
rect 12768 6712 12774 6724
rect 12820 6712 12848 6743
rect 12768 6684 12848 6712
rect 12768 6672 12774 6684
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 2498 6644 2504 6656
rect 2004 6616 2504 6644
rect 2004 6604 2010 6616
rect 2498 6604 2504 6616
rect 2556 6644 2562 6656
rect 2593 6647 2651 6653
rect 2593 6644 2605 6647
rect 2556 6616 2605 6644
rect 2556 6604 2562 6616
rect 2593 6613 2605 6616
rect 2639 6613 2651 6647
rect 3878 6644 3884 6656
rect 3839 6616 3884 6644
rect 2593 6607 2651 6613
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 7006 6604 7012 6656
rect 7064 6644 7070 6656
rect 7653 6647 7711 6653
rect 7653 6644 7665 6647
rect 7064 6616 7665 6644
rect 7064 6604 7070 6616
rect 7653 6613 7665 6616
rect 7699 6613 7711 6647
rect 7653 6607 7711 6613
rect 1104 6554 22816 6576
rect 1104 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 12982 6554
rect 13034 6502 13046 6554
rect 13098 6502 13110 6554
rect 13162 6502 13174 6554
rect 13226 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 22816 6554
rect 1104 6480 22816 6502
rect 14 6400 20 6452
rect 72 6440 78 6452
rect 3421 6443 3479 6449
rect 3421 6440 3433 6443
rect 72 6412 3433 6440
rect 72 6400 78 6412
rect 3421 6409 3433 6412
rect 3467 6409 3479 6443
rect 3786 6440 3792 6452
rect 3747 6412 3792 6440
rect 3421 6403 3479 6409
rect 2130 6372 2136 6384
rect 2091 6344 2136 6372
rect 2130 6332 2136 6344
rect 2188 6332 2194 6384
rect 3436 6304 3464 6403
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 5261 6443 5319 6449
rect 5261 6409 5273 6443
rect 5307 6440 5319 6443
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 5307 6412 5457 6440
rect 5307 6409 5319 6412
rect 5261 6403 5319 6409
rect 5445 6409 5457 6412
rect 5491 6440 5503 6443
rect 5534 6440 5540 6452
rect 5491 6412 5540 6440
rect 5491 6409 5503 6412
rect 5445 6403 5503 6409
rect 5534 6400 5540 6412
rect 5592 6440 5598 6452
rect 6178 6440 6184 6452
rect 5592 6412 6184 6440
rect 5592 6400 5598 6412
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 6362 6440 6368 6452
rect 6323 6412 6368 6440
rect 6362 6400 6368 6412
rect 6420 6400 6426 6452
rect 9125 6443 9183 6449
rect 9125 6409 9137 6443
rect 9171 6440 9183 6443
rect 9858 6440 9864 6452
rect 9171 6412 9864 6440
rect 9171 6409 9183 6412
rect 9125 6403 9183 6409
rect 9858 6400 9864 6412
rect 9916 6440 9922 6452
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 9916 6412 10517 6440
rect 9916 6400 9922 6412
rect 10505 6409 10517 6412
rect 10551 6409 10563 6443
rect 10505 6403 10563 6409
rect 3878 6332 3884 6384
rect 3936 6372 3942 6384
rect 4065 6375 4123 6381
rect 4065 6372 4077 6375
rect 3936 6344 4077 6372
rect 3936 6332 3942 6344
rect 4065 6341 4077 6344
rect 4111 6372 4123 6375
rect 6454 6372 6460 6384
rect 4111 6344 6460 6372
rect 4111 6341 4123 6344
rect 4065 6335 4123 6341
rect 6454 6332 6460 6344
rect 6512 6332 6518 6384
rect 3786 6304 3792 6316
rect 3436 6276 3792 6304
rect 3786 6264 3792 6276
rect 3844 6304 3850 6316
rect 5813 6307 5871 6313
rect 3844 6276 4384 6304
rect 3844 6264 3850 6276
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6205 4307 6239
rect 4356 6236 4384 6276
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 11054 6304 11060 6316
rect 5859 6276 11060 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 11054 6264 11060 6276
rect 11112 6264 11118 6316
rect 11238 6304 11244 6316
rect 11199 6276 11244 6304
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 12342 6264 12348 6316
rect 12400 6304 12406 6316
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 12400 6276 12449 6304
rect 12400 6264 12406 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 12710 6264 12716 6316
rect 12768 6304 12774 6316
rect 13633 6307 13691 6313
rect 13633 6304 13645 6307
rect 12768 6276 13645 6304
rect 12768 6264 12774 6276
rect 13633 6273 13645 6276
rect 13679 6273 13691 6307
rect 13633 6267 13691 6273
rect 4525 6239 4583 6245
rect 4525 6236 4537 6239
rect 4356 6208 4537 6236
rect 4249 6199 4307 6205
rect 4525 6205 4537 6208
rect 4571 6205 4583 6239
rect 4525 6199 4583 6205
rect 5604 6239 5662 6245
rect 5604 6205 5616 6239
rect 5650 6236 5662 6239
rect 5718 6236 5724 6248
rect 5650 6208 5724 6236
rect 5650 6205 5662 6208
rect 5604 6199 5662 6205
rect 1394 6128 1400 6180
rect 1452 6168 1458 6180
rect 1581 6171 1639 6177
rect 1581 6168 1593 6171
rect 1452 6140 1593 6168
rect 1452 6128 1458 6140
rect 1581 6137 1593 6140
rect 1627 6137 1639 6171
rect 1581 6131 1639 6137
rect 1670 6128 1676 6180
rect 1728 6168 1734 6180
rect 4264 6168 4292 6199
rect 5718 6196 5724 6208
rect 5776 6236 5782 6248
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 5776 6208 6009 6236
rect 5776 6196 5782 6208
rect 5997 6205 6009 6208
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 6178 6196 6184 6248
rect 6236 6236 6242 6248
rect 7742 6236 7748 6248
rect 6236 6208 7748 6236
rect 6236 6196 6242 6208
rect 7742 6196 7748 6208
rect 7800 6196 7806 6248
rect 8113 6239 8171 6245
rect 8113 6205 8125 6239
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 8757 6239 8815 6245
rect 8757 6205 8769 6239
rect 8803 6236 8815 6239
rect 9585 6239 9643 6245
rect 9585 6236 9597 6239
rect 8803 6208 9597 6236
rect 8803 6205 8815 6208
rect 8757 6199 8815 6205
rect 9585 6205 9597 6208
rect 9631 6236 9643 6239
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 9631 6208 10793 6236
rect 9631 6205 9643 6208
rect 9585 6199 9643 6205
rect 10781 6205 10793 6208
rect 10827 6205 10839 6239
rect 10781 6199 10839 6205
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6236 12127 6239
rect 12115 6208 12801 6236
rect 12115 6205 12127 6208
rect 12069 6199 12127 6205
rect 5077 6171 5135 6177
rect 5077 6168 5089 6171
rect 1728 6140 1773 6168
rect 4264 6140 5089 6168
rect 1728 6128 1734 6140
rect 5077 6137 5089 6140
rect 5123 6168 5135 6171
rect 5442 6168 5448 6180
rect 5123 6140 5448 6168
rect 5123 6137 5135 6140
rect 5077 6131 5135 6137
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 8128 6168 8156 6199
rect 7024 6140 8156 6168
rect 7024 6112 7052 6140
rect 2038 6060 2044 6112
rect 2096 6100 2102 6112
rect 2498 6100 2504 6112
rect 2096 6072 2504 6100
rect 2096 6060 2102 6072
rect 2498 6060 2504 6072
rect 2556 6060 2562 6112
rect 2866 6100 2872 6112
rect 2827 6072 2872 6100
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 3878 6060 3884 6112
rect 3936 6100 3942 6112
rect 5261 6103 5319 6109
rect 5261 6100 5273 6103
rect 3936 6072 5273 6100
rect 3936 6060 3942 6072
rect 5261 6069 5273 6072
rect 5307 6069 5319 6103
rect 7006 6100 7012 6112
rect 6967 6072 7012 6100
rect 5261 6063 5319 6069
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 7466 6100 7472 6112
rect 7427 6072 7472 6100
rect 7466 6060 7472 6072
rect 7524 6100 7530 6112
rect 8110 6100 8116 6112
rect 7524 6072 8116 6100
rect 7524 6060 7530 6072
rect 8110 6060 8116 6072
rect 8168 6100 8174 6112
rect 8496 6100 8524 6199
rect 9950 6177 9956 6180
rect 9493 6171 9551 6177
rect 9493 6137 9505 6171
rect 9539 6168 9551 6171
rect 9947 6168 9956 6177
rect 9539 6140 9956 6168
rect 9539 6137 9551 6140
rect 9493 6131 9551 6137
rect 9947 6131 9956 6140
rect 9950 6128 9956 6131
rect 10008 6128 10014 6180
rect 11885 6171 11943 6177
rect 11885 6137 11897 6171
rect 11931 6168 11943 6171
rect 12250 6168 12256 6180
rect 11931 6140 12256 6168
rect 11931 6137 11943 6140
rect 11885 6131 11943 6137
rect 12250 6128 12256 6140
rect 12308 6128 12314 6180
rect 12773 6177 12801 6208
rect 13722 6196 13728 6248
rect 13780 6236 13786 6248
rect 13814 6236 13820 6248
rect 13780 6208 13820 6236
rect 13780 6196 13786 6208
rect 13814 6196 13820 6208
rect 13872 6236 13878 6248
rect 14185 6239 14243 6245
rect 14185 6236 14197 6239
rect 13872 6208 14197 6236
rect 13872 6196 13878 6208
rect 14185 6205 14197 6208
rect 14231 6236 14243 6239
rect 14369 6239 14427 6245
rect 14369 6236 14381 6239
rect 14231 6208 14381 6236
rect 14231 6205 14243 6208
rect 14185 6199 14243 6205
rect 14369 6205 14381 6208
rect 14415 6205 14427 6239
rect 14369 6199 14427 6205
rect 14458 6196 14464 6248
rect 14516 6236 14522 6248
rect 14829 6239 14887 6245
rect 14829 6236 14841 6239
rect 14516 6208 14841 6236
rect 14516 6196 14522 6208
rect 14829 6205 14841 6208
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 12758 6171 12816 6177
rect 12758 6137 12770 6171
rect 12804 6137 12816 6171
rect 15102 6168 15108 6180
rect 15063 6140 15108 6168
rect 12758 6131 12816 6137
rect 15102 6128 15108 6140
rect 15160 6128 15166 6180
rect 8168 6072 8524 6100
rect 9968 6100 9996 6128
rect 11790 6100 11796 6112
rect 9968 6072 11796 6100
rect 8168 6060 8174 6072
rect 11790 6060 11796 6072
rect 11848 6100 11854 6112
rect 12069 6103 12127 6109
rect 12069 6100 12081 6103
rect 11848 6072 12081 6100
rect 11848 6060 11854 6072
rect 12069 6069 12081 6072
rect 12115 6100 12127 6103
rect 12161 6103 12219 6109
rect 12161 6100 12173 6103
rect 12115 6072 12173 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12161 6069 12173 6072
rect 12207 6069 12219 6103
rect 12268 6100 12296 6128
rect 13357 6103 13415 6109
rect 13357 6100 13369 6103
rect 12268 6072 13369 6100
rect 12161 6063 12219 6069
rect 13357 6069 13369 6072
rect 13403 6069 13415 6103
rect 13357 6063 13415 6069
rect 1104 6010 22816 6032
rect 1104 5958 8982 6010
rect 9034 5958 9046 6010
rect 9098 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 17174 6010
rect 17226 5958 22816 6010
rect 1104 5936 22816 5958
rect 2406 5896 2412 5908
rect 2367 5868 2412 5896
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 2590 5856 2596 5908
rect 2648 5896 2654 5908
rect 2961 5899 3019 5905
rect 2961 5896 2973 5899
rect 2648 5868 2973 5896
rect 2648 5856 2654 5868
rect 2961 5865 2973 5868
rect 3007 5865 3019 5899
rect 2961 5859 3019 5865
rect 3881 5899 3939 5905
rect 3881 5865 3893 5899
rect 3927 5896 3939 5899
rect 4522 5896 4528 5908
rect 3927 5868 4528 5896
rect 3927 5865 3939 5868
rect 3881 5859 3939 5865
rect 4522 5856 4528 5868
rect 4580 5856 4586 5908
rect 8018 5896 8024 5908
rect 7979 5868 8024 5896
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 8757 5899 8815 5905
rect 8757 5865 8769 5899
rect 8803 5896 8815 5899
rect 9306 5896 9312 5908
rect 8803 5868 9312 5896
rect 8803 5865 8815 5868
rect 8757 5859 8815 5865
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 12802 5896 12808 5908
rect 12763 5868 12808 5896
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 14458 5896 14464 5908
rect 14419 5868 14464 5896
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 15102 5856 15108 5908
rect 15160 5896 15166 5908
rect 15562 5896 15568 5908
rect 15160 5868 15568 5896
rect 15160 5856 15166 5868
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 1670 5788 1676 5840
rect 1728 5828 1734 5840
rect 2133 5831 2191 5837
rect 2133 5828 2145 5831
rect 1728 5800 2145 5828
rect 1728 5788 1734 5800
rect 2133 5797 2145 5800
rect 2179 5828 2191 5831
rect 2866 5828 2872 5840
rect 2179 5800 2872 5828
rect 2179 5797 2191 5800
rect 2133 5791 2191 5797
rect 2866 5788 2872 5800
rect 2924 5788 2930 5840
rect 5077 5831 5135 5837
rect 5077 5797 5089 5831
rect 5123 5828 5135 5831
rect 7006 5828 7012 5840
rect 5123 5800 7012 5828
rect 5123 5797 5135 5800
rect 5077 5791 5135 5797
rect 7006 5788 7012 5800
rect 7064 5788 7070 5840
rect 9398 5788 9404 5840
rect 9456 5828 9462 5840
rect 9456 5800 10235 5828
rect 9456 5788 9462 5800
rect 1946 5760 1952 5772
rect 1907 5732 1952 5760
rect 1946 5720 1952 5732
rect 2004 5720 2010 5772
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4341 5763 4399 5769
rect 4341 5760 4353 5763
rect 4212 5732 4353 5760
rect 4212 5720 4218 5732
rect 4341 5729 4353 5732
rect 4387 5760 4399 5763
rect 5442 5760 5448 5772
rect 4387 5732 5448 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 5442 5720 5448 5732
rect 5500 5720 5506 5772
rect 5994 5760 6000 5772
rect 5955 5732 6000 5760
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 8202 5760 8208 5772
rect 8163 5732 8208 5760
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 10207 5769 10235 5800
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 9876 5732 10057 5760
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 4709 5695 4767 5701
rect 4580 5664 4660 5692
rect 4580 5652 4586 5664
rect 1394 5584 1400 5636
rect 1452 5624 1458 5636
rect 4632 5633 4660 5664
rect 4709 5661 4721 5695
rect 4755 5692 4767 5695
rect 7742 5692 7748 5704
rect 4755 5664 5396 5692
rect 7655 5664 7748 5692
rect 4755 5661 4767 5664
rect 4709 5655 4767 5661
rect 2777 5627 2835 5633
rect 2777 5624 2789 5627
rect 1452 5596 2789 5624
rect 1452 5584 1458 5596
rect 2777 5593 2789 5596
rect 2823 5593 2835 5627
rect 2777 5587 2835 5593
rect 4617 5627 4675 5633
rect 4617 5593 4629 5627
rect 4663 5624 4675 5627
rect 4890 5624 4896 5636
rect 4663 5596 4896 5624
rect 4663 5593 4675 5596
rect 4617 5587 4675 5593
rect 4890 5584 4896 5596
rect 4948 5584 4954 5636
rect 5368 5568 5396 5664
rect 7742 5652 7748 5664
rect 7800 5692 7806 5704
rect 9490 5692 9496 5704
rect 7800 5664 9496 5692
rect 7800 5652 7806 5664
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 8343 5627 8401 5633
rect 8343 5593 8355 5627
rect 8389 5624 8401 5627
rect 9398 5624 9404 5636
rect 8389 5596 9404 5624
rect 8389 5593 8401 5596
rect 8343 5587 8401 5593
rect 9398 5584 9404 5596
rect 9456 5584 9462 5636
rect 3786 5516 3792 5568
rect 3844 5556 3850 5568
rect 4338 5556 4344 5568
rect 3844 5528 4344 5556
rect 3844 5516 3850 5528
rect 4338 5516 4344 5528
rect 4396 5556 4402 5568
rect 4479 5559 4537 5565
rect 4479 5556 4491 5559
rect 4396 5528 4491 5556
rect 4396 5516 4402 5528
rect 4479 5525 4491 5528
rect 4525 5525 4537 5559
rect 5350 5556 5356 5568
rect 5311 5528 5356 5556
rect 4479 5519 4537 5525
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 5721 5559 5779 5565
rect 5721 5556 5733 5559
rect 5684 5528 5733 5556
rect 5684 5516 5690 5528
rect 5721 5525 5733 5528
rect 5767 5525 5779 5559
rect 6178 5556 6184 5568
rect 6139 5528 6184 5556
rect 5721 5519 5779 5525
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 7834 5516 7840 5568
rect 7892 5556 7898 5568
rect 9876 5565 9904 5732
rect 10045 5729 10057 5732
rect 10091 5729 10103 5763
rect 10045 5723 10103 5729
rect 10192 5763 10250 5769
rect 10192 5729 10204 5763
rect 10238 5760 10250 5763
rect 11422 5760 11428 5772
rect 10238 5732 11428 5760
rect 10238 5729 10250 5732
rect 10192 5723 10250 5729
rect 11422 5720 11428 5732
rect 11480 5720 11486 5772
rect 12250 5720 12256 5772
rect 12308 5760 12314 5772
rect 12621 5763 12679 5769
rect 12621 5760 12633 5763
rect 12308 5732 12633 5760
rect 12308 5720 12314 5732
rect 12621 5729 12633 5732
rect 12667 5729 12679 5763
rect 12621 5723 12679 5729
rect 9950 5652 9956 5704
rect 10008 5692 10014 5704
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 10008 5664 10425 5692
rect 10008 5652 10014 5664
rect 10413 5661 10425 5664
rect 10459 5692 10471 5695
rect 10502 5692 10508 5704
rect 10459 5664 10508 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5692 10839 5695
rect 14458 5692 14464 5704
rect 10827 5664 14464 5692
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 10321 5627 10379 5633
rect 10321 5624 10333 5627
rect 10100 5596 10333 5624
rect 10100 5584 10106 5596
rect 10321 5593 10333 5596
rect 10367 5593 10379 5627
rect 10321 5587 10379 5593
rect 9861 5559 9919 5565
rect 9861 5556 9873 5559
rect 7892 5528 9873 5556
rect 7892 5516 7898 5528
rect 9861 5525 9873 5528
rect 9907 5525 9919 5559
rect 9861 5519 9919 5525
rect 1104 5466 22816 5488
rect 1104 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 12982 5466
rect 13034 5414 13046 5466
rect 13098 5414 13110 5466
rect 13162 5414 13174 5466
rect 13226 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 22816 5466
rect 1104 5392 22816 5414
rect 2961 5355 3019 5361
rect 2961 5321 2973 5355
rect 3007 5352 3019 5355
rect 3786 5352 3792 5364
rect 3007 5324 3792 5352
rect 3007 5321 3019 5324
rect 2961 5315 3019 5321
rect 2976 5284 3004 5315
rect 3786 5312 3792 5324
rect 3844 5312 3850 5364
rect 4522 5352 4528 5364
rect 4483 5324 4528 5352
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 5997 5355 6055 5361
rect 5997 5352 6009 5355
rect 5500 5324 6009 5352
rect 5500 5312 5506 5324
rect 5997 5321 6009 5324
rect 6043 5321 6055 5355
rect 6454 5352 6460 5364
rect 6415 5324 6460 5352
rect 5997 5315 6055 5321
rect 6454 5312 6460 5324
rect 6512 5352 6518 5364
rect 9769 5355 9827 5361
rect 9769 5352 9781 5355
rect 6512 5324 9781 5352
rect 6512 5312 6518 5324
rect 9769 5321 9781 5324
rect 9815 5321 9827 5355
rect 9950 5352 9956 5364
rect 9911 5324 9956 5352
rect 9769 5315 9827 5321
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 10042 5312 10048 5364
rect 10100 5352 10106 5364
rect 10321 5355 10379 5361
rect 10321 5352 10333 5355
rect 10100 5324 10333 5352
rect 10100 5312 10106 5324
rect 10321 5321 10333 5324
rect 10367 5321 10379 5355
rect 10321 5315 10379 5321
rect 2240 5256 3004 5284
rect 5261 5287 5319 5293
rect 2240 5157 2268 5256
rect 5261 5253 5273 5287
rect 5307 5284 5319 5287
rect 5534 5284 5540 5296
rect 5307 5256 5540 5284
rect 5307 5253 5319 5256
rect 5261 5247 5319 5253
rect 5534 5244 5540 5256
rect 5592 5284 5598 5296
rect 9858 5284 9864 5296
rect 5592 5256 9864 5284
rect 5592 5244 5598 5256
rect 9858 5244 9864 5256
rect 9916 5244 9922 5296
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5216 2651 5219
rect 3602 5216 3608 5228
rect 2639 5188 3608 5216
rect 2639 5185 2651 5188
rect 2593 5179 2651 5185
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 5350 5216 5356 5228
rect 4212 5188 4257 5216
rect 4816 5188 5356 5216
rect 4212 5176 4218 5188
rect 2225 5151 2283 5157
rect 2225 5117 2237 5151
rect 2271 5117 2283 5151
rect 2225 5111 2283 5117
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5148 3387 5151
rect 3513 5151 3571 5157
rect 3513 5148 3525 5151
rect 3375 5120 3525 5148
rect 3375 5117 3387 5120
rect 3329 5111 3387 5117
rect 3513 5117 3525 5120
rect 3559 5117 3571 5151
rect 3513 5111 3571 5117
rect 1854 5040 1860 5092
rect 1912 5080 1918 5092
rect 1949 5083 2007 5089
rect 1949 5080 1961 5083
rect 1912 5052 1961 5080
rect 1912 5040 1918 5052
rect 1949 5049 1961 5052
rect 1995 5080 2007 5083
rect 2041 5083 2099 5089
rect 2041 5080 2053 5083
rect 1995 5052 2053 5080
rect 1995 5049 2007 5052
rect 1949 5043 2007 5049
rect 2041 5049 2053 5052
rect 2087 5080 2099 5083
rect 3344 5080 3372 5111
rect 2087 5052 3372 5080
rect 2087 5049 2099 5052
rect 2041 5043 2099 5049
rect 3786 4972 3792 5024
rect 3844 5012 3850 5024
rect 3970 5012 3976 5024
rect 3844 4984 3976 5012
rect 3844 4972 3850 4984
rect 3970 4972 3976 4984
rect 4028 5012 4034 5024
rect 4816 5021 4844 5188
rect 5350 5176 5356 5188
rect 5408 5216 5414 5228
rect 9493 5219 9551 5225
rect 9493 5216 9505 5219
rect 5408 5188 9505 5216
rect 5408 5176 5414 5188
rect 9493 5185 9505 5188
rect 9539 5216 9551 5219
rect 9968 5216 9996 5312
rect 10183 5287 10241 5293
rect 10183 5284 10195 5287
rect 9539 5188 9996 5216
rect 10060 5256 10195 5284
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 4982 5148 4988 5160
rect 4943 5120 4988 5148
rect 4982 5108 4988 5120
rect 5040 5108 5046 5160
rect 5132 5151 5190 5157
rect 5132 5117 5144 5151
rect 5178 5148 5190 5151
rect 6454 5148 6460 5160
rect 5178 5120 6460 5148
rect 5178 5117 5190 5120
rect 5132 5111 5190 5117
rect 6454 5108 6460 5120
rect 6512 5108 6518 5160
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 6860 5151 6918 5157
rect 6860 5148 6872 5151
rect 6788 5120 6872 5148
rect 6788 5108 6794 5120
rect 6860 5117 6872 5120
rect 6906 5148 6918 5151
rect 7285 5151 7343 5157
rect 7285 5148 7297 5151
rect 6906 5120 7297 5148
rect 6906 5117 6918 5120
rect 6860 5111 6918 5117
rect 7285 5117 7297 5120
rect 7331 5117 7343 5151
rect 7285 5111 7343 5117
rect 7745 5151 7803 5157
rect 7745 5117 7757 5151
rect 7791 5148 7803 5151
rect 8570 5148 8576 5160
rect 7791 5120 8576 5148
rect 7791 5117 7803 5120
rect 7745 5111 7803 5117
rect 8570 5108 8576 5120
rect 8628 5108 8634 5160
rect 9766 5148 9772 5160
rect 9679 5120 9772 5148
rect 9766 5108 9772 5120
rect 9824 5148 9830 5160
rect 10060 5148 10088 5256
rect 10183 5253 10195 5256
rect 10229 5253 10241 5287
rect 10336 5284 10364 5315
rect 10410 5312 10416 5364
rect 10468 5352 10474 5364
rect 10689 5355 10747 5361
rect 10689 5352 10701 5355
rect 10468 5324 10701 5352
rect 10468 5312 10474 5324
rect 10689 5321 10701 5324
rect 10735 5352 10747 5355
rect 12066 5352 12072 5364
rect 10735 5324 12072 5352
rect 10735 5321 10747 5324
rect 10689 5315 10747 5321
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 12250 5352 12256 5364
rect 12211 5324 12256 5352
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 10778 5284 10784 5296
rect 10336 5256 10784 5284
rect 10183 5247 10241 5253
rect 10778 5244 10784 5256
rect 10836 5284 10842 5296
rect 11057 5287 11115 5293
rect 11057 5284 11069 5287
rect 10836 5256 11069 5284
rect 10836 5244 10842 5256
rect 11057 5253 11069 5256
rect 11103 5253 11115 5287
rect 11422 5284 11428 5296
rect 11383 5256 11428 5284
rect 11057 5247 11115 5253
rect 11422 5244 11428 5256
rect 11480 5244 11486 5296
rect 10413 5219 10471 5225
rect 10413 5185 10425 5219
rect 10459 5216 10471 5219
rect 10502 5216 10508 5228
rect 10459 5188 10508 5216
rect 10459 5185 10471 5188
rect 10413 5179 10471 5185
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 15562 5216 15568 5228
rect 15523 5188 15568 5216
rect 15562 5176 15568 5188
rect 15620 5176 15626 5228
rect 9824 5120 10088 5148
rect 9824 5108 9830 5120
rect 12158 5108 12164 5160
rect 12216 5148 12222 5160
rect 12472 5151 12530 5157
rect 12472 5148 12484 5151
rect 12216 5120 12484 5148
rect 12216 5108 12222 5120
rect 12472 5117 12484 5120
rect 12518 5148 12530 5151
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12518 5120 12909 5148
rect 12518 5117 12530 5120
rect 12472 5111 12530 5117
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 13538 5148 13544 5160
rect 13451 5120 13544 5148
rect 12897 5111 12955 5117
rect 13538 5108 13544 5120
rect 13596 5148 13602 5160
rect 13633 5151 13691 5157
rect 13633 5148 13645 5151
rect 13596 5120 13645 5148
rect 13596 5108 13602 5120
rect 13633 5117 13645 5120
rect 13679 5117 13691 5151
rect 14182 5148 14188 5160
rect 14095 5120 14188 5148
rect 13633 5111 13691 5117
rect 14182 5108 14188 5120
rect 14240 5148 14246 5160
rect 14458 5148 14464 5160
rect 14240 5120 14464 5148
rect 14240 5108 14246 5120
rect 14458 5108 14464 5120
rect 14516 5108 14522 5160
rect 6963 5083 7021 5089
rect 6963 5049 6975 5083
rect 7009 5080 7021 5083
rect 8662 5080 8668 5092
rect 7009 5052 8668 5080
rect 7009 5049 7021 5052
rect 6963 5043 7021 5049
rect 8662 5040 8668 5052
rect 8720 5040 8726 5092
rect 8941 5083 8999 5089
rect 8941 5049 8953 5083
rect 8987 5080 8999 5083
rect 9306 5080 9312 5092
rect 8987 5052 9312 5080
rect 8987 5049 8999 5052
rect 8941 5043 8999 5049
rect 9306 5040 9312 5052
rect 9364 5040 9370 5092
rect 9490 5040 9496 5092
rect 9548 5080 9554 5092
rect 10045 5083 10103 5089
rect 10045 5080 10057 5083
rect 9548 5052 10057 5080
rect 9548 5040 9554 5052
rect 10045 5049 10057 5052
rect 10091 5080 10103 5083
rect 11793 5083 11851 5089
rect 11793 5080 11805 5083
rect 10091 5052 11805 5080
rect 10091 5049 10103 5052
rect 10045 5043 10103 5049
rect 11793 5049 11805 5052
rect 11839 5049 11851 5083
rect 11793 5043 11851 5049
rect 11974 5040 11980 5092
rect 12032 5080 12038 5092
rect 12575 5083 12633 5089
rect 12575 5080 12587 5083
rect 12032 5052 12587 5080
rect 12032 5040 12038 5052
rect 12575 5049 12587 5052
rect 12621 5049 12633 5083
rect 14366 5080 14372 5092
rect 14327 5052 14372 5080
rect 12575 5043 12633 5049
rect 14366 5040 14372 5052
rect 14424 5040 14430 5092
rect 15886 5083 15944 5089
rect 15886 5049 15898 5083
rect 15932 5049 15944 5083
rect 15886 5043 15944 5049
rect 4801 5015 4859 5021
rect 4801 5012 4813 5015
rect 4028 4984 4813 5012
rect 4028 4972 4034 4984
rect 4801 4981 4813 4984
rect 4847 4981 4859 5015
rect 5626 5012 5632 5024
rect 5587 4984 5632 5012
rect 4801 4975 4859 4981
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 8113 5015 8171 5021
rect 8113 4981 8125 5015
rect 8159 5012 8171 5015
rect 8202 5012 8208 5024
rect 8159 4984 8208 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 8202 4972 8208 4984
rect 8260 5012 8266 5024
rect 8846 5012 8852 5024
rect 8260 4984 8852 5012
rect 8260 4972 8266 4984
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 15378 5012 15384 5024
rect 15339 4984 15384 5012
rect 15378 4972 15384 4984
rect 15436 5012 15442 5024
rect 15901 5012 15929 5043
rect 16482 5012 16488 5024
rect 15436 4984 15929 5012
rect 16443 4984 16488 5012
rect 15436 4972 15442 4984
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 1104 4922 22816 4944
rect 1104 4870 8982 4922
rect 9034 4870 9046 4922
rect 9098 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 17174 4922
rect 17226 4870 22816 4922
rect 1104 4848 22816 4870
rect 1946 4808 1952 4820
rect 1907 4780 1952 4808
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 4338 4808 4344 4820
rect 4299 4780 4344 4808
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 5534 4808 5540 4820
rect 5495 4780 5540 4808
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 5994 4808 6000 4820
rect 5955 4780 6000 4808
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7101 4811 7159 4817
rect 7101 4808 7113 4811
rect 7064 4780 7113 4808
rect 7064 4768 7070 4780
rect 7101 4777 7113 4780
rect 7147 4777 7159 4811
rect 7101 4771 7159 4777
rect 2317 4743 2375 4749
rect 2317 4709 2329 4743
rect 2363 4740 2375 4743
rect 4614 4740 4620 4752
rect 2363 4712 4620 4740
rect 2363 4709 2375 4712
rect 2317 4703 2375 4709
rect 1464 4675 1522 4681
rect 1464 4641 1476 4675
rect 1510 4672 1522 4675
rect 1578 4672 1584 4684
rect 1510 4644 1584 4672
rect 1510 4641 1522 4644
rect 1464 4635 1522 4641
rect 1578 4632 1584 4644
rect 1636 4632 1642 4684
rect 2682 4672 2688 4684
rect 2643 4644 2688 4672
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 2976 4681 3004 4712
rect 4614 4700 4620 4712
rect 4672 4740 4678 4752
rect 4672 4712 5120 4740
rect 4672 4700 4678 4712
rect 2961 4675 3019 4681
rect 2961 4641 2973 4675
rect 3007 4641 3019 4675
rect 2961 4635 3019 4641
rect 4062 4632 4068 4684
rect 4120 4672 4126 4684
rect 4522 4672 4528 4684
rect 4120 4644 4528 4672
rect 4120 4632 4126 4644
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 5092 4681 5120 4712
rect 6178 4700 6184 4752
rect 6236 4740 6242 4752
rect 6273 4743 6331 4749
rect 6273 4740 6285 4743
rect 6236 4712 6285 4740
rect 6236 4700 6242 4712
rect 6273 4709 6285 4712
rect 6319 4709 6331 4743
rect 7116 4740 7144 4771
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 13219 4811 13277 4817
rect 13219 4808 13231 4811
rect 8812 4780 13231 4808
rect 8812 4768 8818 4780
rect 13219 4777 13231 4780
rect 13265 4777 13277 4811
rect 13219 4771 13277 4777
rect 13725 4811 13783 4817
rect 13725 4777 13737 4811
rect 13771 4808 13783 4811
rect 14182 4808 14188 4820
rect 13771 4780 14188 4808
rect 13771 4777 13783 4780
rect 13725 4771 13783 4777
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 14277 4811 14335 4817
rect 14277 4777 14289 4811
rect 14323 4808 14335 4811
rect 14366 4808 14372 4820
rect 14323 4780 14372 4808
rect 14323 4777 14335 4780
rect 14277 4771 14335 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 7742 4740 7748 4752
rect 7116 4712 7748 4740
rect 6273 4703 6331 4709
rect 7742 4700 7748 4712
rect 7800 4740 7806 4752
rect 9493 4743 9551 4749
rect 7800 4712 8248 4740
rect 7800 4700 7806 4712
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 5626 4672 5632 4684
rect 5123 4644 5632 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4672 7711 4675
rect 7834 4672 7840 4684
rect 7699 4644 7840 4672
rect 7699 4641 7711 4644
rect 7653 4635 7711 4641
rect 3142 4604 3148 4616
rect 3103 4576 3148 4604
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 3970 4564 3976 4616
rect 4028 4604 4034 4616
rect 4982 4604 4988 4616
rect 4028 4576 4988 4604
rect 4028 4564 4034 4576
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4604 5319 4607
rect 5350 4604 5356 4616
rect 5307 4576 5356 4604
rect 5307 4573 5319 4576
rect 5261 4567 5319 4573
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4604 6239 4607
rect 6454 4604 6460 4616
rect 6227 4576 6460 4604
rect 6227 4573 6239 4576
rect 6181 4567 6239 4573
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 1535 4539 1593 4545
rect 1535 4505 1547 4539
rect 1581 4536 1593 4539
rect 4706 4536 4712 4548
rect 1581 4508 4712 4536
rect 1581 4505 1593 4508
rect 1535 4499 1593 4505
rect 4706 4496 4712 4508
rect 4764 4496 4770 4548
rect 6733 4539 6791 4545
rect 6733 4505 6745 4539
rect 6779 4536 6791 4539
rect 7650 4536 7656 4548
rect 6779 4508 7656 4536
rect 6779 4505 6791 4508
rect 6733 4499 6791 4505
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 7469 4471 7527 4477
rect 7469 4468 7481 4471
rect 6880 4440 7481 4468
rect 6880 4428 6886 4440
rect 7469 4437 7481 4440
rect 7515 4468 7527 4471
rect 7760 4468 7788 4644
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 8220 4681 8248 4712
rect 9493 4709 9505 4743
rect 9539 4740 9551 4743
rect 9766 4740 9772 4752
rect 9539 4712 9772 4740
rect 9539 4709 9551 4712
rect 9493 4703 9551 4709
rect 9766 4700 9772 4712
rect 9824 4700 9830 4752
rect 10778 4740 10784 4752
rect 10739 4712 10784 4740
rect 10778 4700 10784 4712
rect 10836 4700 10842 4752
rect 11695 4743 11753 4749
rect 11695 4709 11707 4743
rect 11741 4740 11753 4743
rect 11790 4740 11796 4752
rect 11741 4712 11796 4740
rect 11741 4709 11753 4712
rect 11695 4703 11753 4709
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 16482 4700 16488 4752
rect 16540 4740 16546 4752
rect 17218 4740 17224 4752
rect 16540 4712 17224 4740
rect 16540 4700 16546 4712
rect 17218 4700 17224 4712
rect 17276 4740 17282 4752
rect 17313 4743 17371 4749
rect 17313 4740 17325 4743
rect 17276 4712 17325 4740
rect 17276 4700 17282 4712
rect 17313 4709 17325 4712
rect 17359 4709 17371 4743
rect 17313 4703 17371 4709
rect 8205 4675 8263 4681
rect 8205 4641 8217 4675
rect 8251 4641 8263 4675
rect 8205 4635 8263 4641
rect 8386 4632 8392 4684
rect 8444 4672 8450 4684
rect 8481 4675 8539 4681
rect 8481 4672 8493 4675
rect 8444 4644 8493 4672
rect 8444 4632 8450 4644
rect 8481 4641 8493 4644
rect 8527 4641 8539 4675
rect 10042 4672 10048 4684
rect 10003 4644 10048 4672
rect 8481 4635 8539 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 10321 4675 10379 4681
rect 10321 4641 10333 4675
rect 10367 4672 10379 4675
rect 10410 4672 10416 4684
rect 10367 4644 10416 4672
rect 10367 4641 10379 4644
rect 10321 4635 10379 4641
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 11054 4632 11060 4684
rect 11112 4672 11118 4684
rect 12526 4672 12532 4684
rect 11112 4644 12532 4672
rect 11112 4632 11118 4644
rect 12526 4632 12532 4644
rect 12584 4632 12590 4684
rect 13148 4675 13206 4681
rect 13148 4641 13160 4675
rect 13194 4672 13206 4675
rect 13446 4672 13452 4684
rect 13194 4644 13452 4672
rect 13194 4641 13206 4644
rect 13148 4635 13206 4641
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 15933 4675 15991 4681
rect 15933 4641 15945 4675
rect 15979 4672 15991 4675
rect 16114 4672 16120 4684
rect 15979 4644 16120 4672
rect 15979 4641 15991 4644
rect 15933 4635 15991 4641
rect 16114 4632 16120 4644
rect 16172 4632 16178 4684
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4604 10563 4607
rect 11146 4604 11152 4616
rect 10551 4576 11152 4604
rect 10551 4573 10563 4576
rect 10505 4567 10563 4573
rect 11146 4564 11152 4576
rect 11204 4604 11210 4616
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 11204 4576 11345 4604
rect 11204 4564 11210 4576
rect 11333 4573 11345 4576
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 17221 4607 17279 4613
rect 17221 4573 17233 4607
rect 17267 4604 17279 4607
rect 17494 4604 17500 4616
rect 17267 4576 17500 4604
rect 17267 4573 17279 4576
rect 17221 4567 17279 4573
rect 17494 4564 17500 4576
rect 17552 4564 17558 4616
rect 17865 4607 17923 4613
rect 17865 4573 17877 4607
rect 17911 4604 17923 4607
rect 18414 4604 18420 4616
rect 17911 4576 18420 4604
rect 17911 4573 17923 4576
rect 17865 4567 17923 4573
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 7515 4440 7788 4468
rect 7515 4437 7527 4440
rect 7469 4431 7527 4437
rect 8754 4428 8760 4480
rect 8812 4468 8818 4480
rect 12250 4468 12256 4480
rect 8812 4440 8857 4468
rect 12211 4440 12256 4468
rect 8812 4428 8818 4440
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 15562 4468 15568 4480
rect 15523 4440 15568 4468
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 18046 4428 18052 4480
rect 18104 4468 18110 4480
rect 18141 4471 18199 4477
rect 18141 4468 18153 4471
rect 18104 4440 18153 4468
rect 18104 4428 18110 4440
rect 18141 4437 18153 4440
rect 18187 4437 18199 4471
rect 18141 4431 18199 4437
rect 1104 4378 22816 4400
rect 1104 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 12982 4378
rect 13034 4326 13046 4378
rect 13098 4326 13110 4378
rect 13162 4326 13174 4378
rect 13226 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 22816 4378
rect 1104 4304 22816 4326
rect 1578 4264 1584 4276
rect 1539 4236 1584 4264
rect 1578 4224 1584 4236
rect 1636 4224 1642 4276
rect 2682 4224 2688 4276
rect 2740 4264 2746 4276
rect 3237 4267 3295 4273
rect 3237 4264 3249 4267
rect 2740 4236 3249 4264
rect 2740 4224 2746 4236
rect 3237 4233 3249 4236
rect 3283 4264 3295 4267
rect 3694 4264 3700 4276
rect 3283 4236 3700 4264
rect 3283 4233 3295 4236
rect 3237 4227 3295 4233
rect 3694 4224 3700 4236
rect 3752 4224 3758 4276
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 4893 4267 4951 4273
rect 4893 4264 4905 4267
rect 4580 4236 4905 4264
rect 4580 4224 4586 4236
rect 4893 4233 4905 4236
rect 4939 4233 4951 4267
rect 4893 4227 4951 4233
rect 5353 4267 5411 4273
rect 5353 4233 5365 4267
rect 5399 4264 5411 4267
rect 6178 4264 6184 4276
rect 5399 4236 6184 4264
rect 5399 4233 5411 4236
rect 5353 4227 5411 4233
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3694 4128 3700 4140
rect 3200 4100 3700 4128
rect 3200 4088 3206 4100
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 4908 4128 4936 4227
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 8205 4267 8263 4273
rect 8205 4233 8217 4267
rect 8251 4264 8263 4267
rect 10042 4264 10048 4276
rect 8251 4236 10048 4264
rect 8251 4233 8263 4236
rect 8205 4227 8263 4233
rect 10042 4224 10048 4236
rect 10100 4224 10106 4276
rect 10410 4224 10416 4276
rect 10468 4264 10474 4276
rect 10689 4267 10747 4273
rect 10689 4264 10701 4267
rect 10468 4236 10701 4264
rect 10468 4224 10474 4236
rect 10689 4233 10701 4236
rect 10735 4233 10747 4267
rect 11146 4264 11152 4276
rect 11107 4236 11152 4264
rect 10689 4227 10747 4233
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 11790 4264 11796 4276
rect 11751 4236 11796 4264
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 13814 4224 13820 4276
rect 13872 4264 13878 4276
rect 14642 4264 14648 4276
rect 13872 4236 14648 4264
rect 13872 4224 13878 4236
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 17218 4264 17224 4276
rect 17179 4236 17224 4264
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 8110 4156 8116 4208
rect 8168 4196 8174 4208
rect 11808 4196 11836 4224
rect 14001 4199 14059 4205
rect 14001 4196 14013 4199
rect 8168 4168 14013 4196
rect 8168 4156 8174 4168
rect 14001 4165 14013 4168
rect 14047 4165 14059 4199
rect 14001 4159 14059 4165
rect 15105 4199 15163 4205
rect 15105 4165 15117 4199
rect 15151 4196 15163 4199
rect 15473 4199 15531 4205
rect 15473 4196 15485 4199
rect 15151 4168 15485 4196
rect 15151 4165 15163 4168
rect 15105 4159 15163 4165
rect 15473 4165 15485 4168
rect 15519 4196 15531 4199
rect 15841 4199 15899 4205
rect 15841 4196 15853 4199
rect 15519 4168 15853 4196
rect 15519 4165 15531 4168
rect 15473 4159 15531 4165
rect 15841 4165 15853 4168
rect 15887 4196 15899 4199
rect 16114 4196 16120 4208
rect 15887 4168 16120 4196
rect 15887 4165 15899 4168
rect 15841 4159 15899 4165
rect 6641 4131 6699 4137
rect 4908 4100 6040 4128
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4029 2559 4063
rect 2501 4023 2559 4029
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4060 2927 4063
rect 3878 4060 3884 4072
rect 2915 4032 3884 4060
rect 2915 4029 2927 4032
rect 2869 4023 2927 4029
rect 2314 3992 2320 4004
rect 2275 3964 2320 3992
rect 2314 3952 2320 3964
rect 2372 3952 2378 4004
rect 2130 3924 2136 3936
rect 2091 3896 2136 3924
rect 2130 3884 2136 3896
rect 2188 3924 2194 3936
rect 2516 3924 2544 4023
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 4798 4020 4804 4072
rect 4856 4060 4862 4072
rect 5480 4063 5538 4069
rect 5480 4060 5492 4063
rect 4856 4032 5492 4060
rect 4856 4020 4862 4032
rect 5480 4029 5492 4032
rect 5526 4060 5538 4063
rect 5905 4063 5963 4069
rect 5905 4060 5917 4063
rect 5526 4032 5917 4060
rect 5526 4029 5538 4032
rect 5480 4023 5538 4029
rect 5905 4029 5917 4032
rect 5951 4029 5963 4063
rect 5905 4023 5963 4029
rect 4018 3995 4076 4001
rect 4018 3992 4030 3995
rect 3528 3964 4030 3992
rect 2188 3896 2544 3924
rect 2188 3884 2194 3896
rect 2590 3884 2596 3936
rect 2648 3924 2654 3936
rect 3528 3933 3556 3964
rect 4018 3961 4030 3964
rect 4064 3992 4076 3995
rect 4522 3992 4528 4004
rect 4064 3964 4528 3992
rect 4064 3961 4076 3964
rect 4018 3955 4076 3961
rect 4522 3952 4528 3964
rect 4580 3952 4586 4004
rect 6012 3992 6040 4100
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 7742 4128 7748 4140
rect 6687 4100 7144 4128
rect 7703 4100 7748 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 6822 4020 6828 4072
rect 6880 4060 6886 4072
rect 7009 4063 7067 4069
rect 7009 4060 7021 4063
rect 6880 4032 7021 4060
rect 6880 4020 6886 4032
rect 7009 4029 7021 4032
rect 7055 4029 7067 4063
rect 7116 4060 7144 4100
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 8754 4088 8760 4140
rect 8812 4128 8818 4140
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 8812 4100 9137 4128
rect 8812 4088 8818 4100
rect 9125 4097 9137 4100
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10413 4131 10471 4137
rect 10413 4128 10425 4131
rect 10100 4100 10425 4128
rect 10100 4088 10106 4100
rect 10413 4097 10425 4100
rect 10459 4097 10471 4131
rect 12526 4128 12532 4140
rect 12487 4100 12532 4128
rect 10413 4091 10471 4097
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 12802 4128 12808 4140
rect 12763 4100 12808 4128
rect 12802 4088 12808 4100
rect 12860 4088 12866 4140
rect 7466 4060 7472 4072
rect 7116 4032 7472 4060
rect 7009 4023 7067 4029
rect 7466 4020 7472 4032
rect 7524 4060 7530 4072
rect 7837 4063 7895 4069
rect 7837 4060 7849 4063
rect 7524 4032 7849 4060
rect 7524 4020 7530 4032
rect 7837 4029 7849 4032
rect 7883 4060 7895 4063
rect 8205 4063 8263 4069
rect 8205 4060 8217 4063
rect 7883 4032 8217 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 8205 4029 8217 4032
rect 8251 4029 8263 4063
rect 8205 4023 8263 4029
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 11368 4063 11426 4069
rect 11368 4060 11380 4063
rect 11204 4032 11380 4060
rect 11204 4020 11210 4032
rect 11368 4029 11380 4032
rect 11414 4029 11426 4063
rect 11368 4023 11426 4029
rect 8386 3992 8392 4004
rect 6012 3964 8392 3992
rect 8386 3952 8392 3964
rect 8444 3952 8450 4004
rect 9446 3995 9504 4001
rect 9446 3961 9458 3995
rect 9492 3961 9504 3995
rect 9446 3955 9504 3961
rect 12253 3995 12311 4001
rect 12253 3961 12265 3995
rect 12299 3992 12311 3995
rect 12621 3995 12679 4001
rect 12621 3992 12633 3995
rect 12299 3964 12633 3992
rect 12299 3961 12311 3964
rect 12253 3955 12311 3961
rect 12621 3961 12633 3964
rect 12667 3992 12679 3995
rect 12894 3992 12900 4004
rect 12667 3964 12900 3992
rect 12667 3961 12679 3964
rect 12621 3955 12679 3961
rect 3513 3927 3571 3933
rect 3513 3924 3525 3927
rect 2648 3896 3525 3924
rect 2648 3884 2654 3896
rect 3513 3893 3525 3896
rect 3559 3893 3571 3927
rect 3513 3887 3571 3893
rect 4154 3884 4160 3936
rect 4212 3924 4218 3936
rect 4617 3927 4675 3933
rect 4617 3924 4629 3927
rect 4212 3896 4629 3924
rect 4212 3884 4218 3896
rect 4617 3893 4629 3896
rect 4663 3893 4675 3927
rect 4617 3887 4675 3893
rect 4798 3884 4804 3936
rect 4856 3924 4862 3936
rect 5583 3927 5641 3933
rect 5583 3924 5595 3927
rect 4856 3896 5595 3924
rect 4856 3884 4862 3896
rect 5583 3893 5595 3896
rect 5629 3893 5641 3927
rect 7282 3924 7288 3936
rect 7243 3896 7288 3924
rect 5583 3887 5641 3893
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8941 3927 8999 3933
rect 8941 3924 8953 3927
rect 8168 3896 8953 3924
rect 8168 3884 8174 3896
rect 8941 3893 8953 3896
rect 8987 3924 8999 3927
rect 9461 3924 9489 3955
rect 12894 3952 12900 3964
rect 12952 3952 12958 4004
rect 14016 3992 14044 4159
rect 16114 4156 16120 4168
rect 16172 4156 16178 4208
rect 14185 4131 14243 4137
rect 14185 4097 14197 4131
rect 14231 4128 14243 4131
rect 14366 4128 14372 4140
rect 14231 4100 14372 4128
rect 14231 4097 14243 4100
rect 14185 4091 14243 4097
rect 14366 4088 14372 4100
rect 14424 4088 14430 4140
rect 16298 4128 16304 4140
rect 16259 4100 16304 4128
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 18414 4128 18420 4140
rect 18375 4100 18420 4128
rect 18414 4088 18420 4100
rect 18472 4088 18478 4140
rect 14506 3995 14564 4001
rect 14506 3992 14518 3995
rect 14016 3964 14518 3992
rect 14506 3961 14518 3964
rect 14552 3992 14564 3995
rect 15378 3992 15384 4004
rect 14552 3964 15384 3992
rect 14552 3961 14564 3964
rect 14506 3955 14564 3961
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 16025 3995 16083 4001
rect 16025 3961 16037 3995
rect 16071 3961 16083 3995
rect 16025 3955 16083 3961
rect 10042 3924 10048 3936
rect 8987 3896 9489 3924
rect 10003 3896 10048 3924
rect 8987 3893 8999 3896
rect 8941 3887 8999 3893
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 11471 3927 11529 3933
rect 11471 3893 11483 3927
rect 11517 3924 11529 3927
rect 12526 3924 12532 3936
rect 11517 3896 12532 3924
rect 11517 3893 11529 3896
rect 11471 3887 11529 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 13446 3924 13452 3936
rect 13407 3896 13452 3924
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 16040 3924 16068 3955
rect 16114 3952 16120 4004
rect 16172 3992 16178 4004
rect 18141 3995 18199 4001
rect 16172 3964 16217 3992
rect 16172 3952 16178 3964
rect 18141 3961 18153 3995
rect 18187 3961 18199 3995
rect 18141 3955 18199 3961
rect 16390 3924 16396 3936
rect 16040 3896 16396 3924
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 17770 3924 17776 3936
rect 17731 3896 17776 3924
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 18046 3884 18052 3936
rect 18104 3924 18110 3936
rect 18156 3924 18184 3955
rect 18230 3952 18236 4004
rect 18288 3992 18294 4004
rect 18288 3964 18333 3992
rect 18288 3952 18294 3964
rect 18104 3896 18184 3924
rect 18104 3884 18110 3896
rect 1104 3834 22816 3856
rect 1104 3782 8982 3834
rect 9034 3782 9046 3834
rect 9098 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 17174 3834
rect 17226 3782 22816 3834
rect 1104 3760 22816 3782
rect 3694 3720 3700 3732
rect 3655 3692 3700 3720
rect 3694 3680 3700 3692
rect 3752 3680 3758 3732
rect 4614 3720 4620 3732
rect 4575 3692 4620 3720
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 5994 3680 6000 3732
rect 6052 3720 6058 3732
rect 6181 3723 6239 3729
rect 6181 3720 6193 3723
rect 6052 3692 6193 3720
rect 6052 3680 6058 3692
rect 6181 3689 6193 3692
rect 6227 3689 6239 3723
rect 6181 3683 6239 3689
rect 7469 3723 7527 3729
rect 7469 3689 7481 3723
rect 7515 3720 7527 3723
rect 7742 3720 7748 3732
rect 7515 3692 7748 3720
rect 7515 3689 7527 3692
rect 7469 3683 7527 3689
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 8478 3720 8484 3732
rect 8439 3692 8484 3720
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 8754 3680 8760 3732
rect 8812 3720 8818 3732
rect 9125 3723 9183 3729
rect 9125 3720 9137 3723
rect 8812 3692 9137 3720
rect 8812 3680 8818 3692
rect 9125 3689 9137 3692
rect 9171 3689 9183 3723
rect 12250 3720 12256 3732
rect 9125 3683 9183 3689
rect 12084 3692 12256 3720
rect 12084 3664 12112 3692
rect 12250 3680 12256 3692
rect 12308 3720 12314 3732
rect 12308 3692 13584 3720
rect 12308 3680 12314 3692
rect 4522 3612 4528 3664
rect 4580 3652 4586 3664
rect 5442 3652 5448 3664
rect 4580 3624 5448 3652
rect 4580 3612 4586 3624
rect 5442 3612 5448 3624
rect 5500 3652 5506 3664
rect 5582 3655 5640 3661
rect 5582 3652 5594 3655
rect 5500 3624 5594 3652
rect 5500 3612 5506 3624
rect 5582 3621 5594 3624
rect 5628 3652 5640 3655
rect 7882 3655 7940 3661
rect 7882 3652 7894 3655
rect 5628 3624 7894 3652
rect 5628 3621 5640 3624
rect 5582 3615 5640 3621
rect 7882 3621 7894 3624
rect 7928 3652 7940 3655
rect 8110 3652 8116 3664
rect 7928 3624 8116 3652
rect 7928 3621 7940 3624
rect 7882 3615 7940 3621
rect 8110 3612 8116 3624
rect 8168 3612 8174 3664
rect 9490 3612 9496 3664
rect 9548 3652 9554 3664
rect 10042 3652 10048 3664
rect 9548 3624 10048 3652
rect 9548 3612 9554 3624
rect 10042 3612 10048 3624
rect 10100 3652 10106 3664
rect 10137 3655 10195 3661
rect 10137 3652 10149 3655
rect 10100 3624 10149 3652
rect 10100 3612 10106 3624
rect 10137 3621 10149 3624
rect 10183 3652 10195 3655
rect 10686 3652 10692 3664
rect 10183 3624 10692 3652
rect 10183 3621 10195 3624
rect 10137 3615 10195 3621
rect 10686 3612 10692 3624
rect 10744 3612 10750 3664
rect 12066 3652 12072 3664
rect 11979 3624 12072 3652
rect 12066 3612 12072 3624
rect 12124 3612 12130 3664
rect 12621 3655 12679 3661
rect 12621 3621 12633 3655
rect 12667 3652 12679 3655
rect 12802 3652 12808 3664
rect 12667 3624 12808 3652
rect 12667 3621 12679 3624
rect 12621 3615 12679 3621
rect 12802 3612 12808 3624
rect 12860 3612 12866 3664
rect 12894 3612 12900 3664
rect 12952 3652 12958 3664
rect 13449 3655 13507 3661
rect 13449 3652 13461 3655
rect 12952 3624 13461 3652
rect 12952 3612 12958 3624
rect 13449 3621 13461 3624
rect 13495 3621 13507 3655
rect 13449 3615 13507 3621
rect 13556 3596 13584 3692
rect 17494 3680 17500 3732
rect 17552 3720 17558 3732
rect 17865 3723 17923 3729
rect 17865 3720 17877 3723
rect 17552 3692 17877 3720
rect 17552 3680 17558 3692
rect 17865 3689 17877 3692
rect 17911 3689 17923 3723
rect 17865 3683 17923 3689
rect 15473 3655 15531 3661
rect 15473 3621 15485 3655
rect 15519 3652 15531 3655
rect 15562 3652 15568 3664
rect 15519 3624 15568 3652
rect 15519 3621 15531 3624
rect 15473 3615 15531 3621
rect 15562 3612 15568 3624
rect 15620 3652 15626 3664
rect 15746 3652 15752 3664
rect 15620 3624 15752 3652
rect 15620 3612 15626 3624
rect 15746 3612 15752 3624
rect 15804 3612 15810 3664
rect 16022 3652 16028 3664
rect 15935 3624 16028 3652
rect 16022 3612 16028 3624
rect 16080 3652 16086 3664
rect 16298 3652 16304 3664
rect 16080 3624 16304 3652
rect 16080 3612 16086 3624
rect 16298 3612 16304 3624
rect 16356 3612 16362 3664
rect 17589 3655 17647 3661
rect 17589 3621 17601 3655
rect 17635 3652 17647 3655
rect 17770 3652 17776 3664
rect 17635 3624 17776 3652
rect 17635 3621 17647 3624
rect 17589 3615 17647 3621
rect 17770 3612 17776 3624
rect 17828 3652 17834 3664
rect 18230 3652 18236 3664
rect 17828 3624 18236 3652
rect 17828 3612 17834 3624
rect 18230 3612 18236 3624
rect 18288 3612 18294 3664
rect 2222 3584 2228 3596
rect 2183 3556 2228 3584
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 2314 3544 2320 3596
rect 2372 3584 2378 3596
rect 2777 3587 2835 3593
rect 2777 3584 2789 3587
rect 2372 3556 2789 3584
rect 2372 3544 2378 3556
rect 2777 3553 2789 3556
rect 2823 3584 2835 3587
rect 3053 3587 3111 3593
rect 3053 3584 3065 3587
rect 2823 3556 3065 3584
rect 2823 3553 2835 3556
rect 2777 3547 2835 3553
rect 3053 3553 3065 3556
rect 3099 3553 3111 3587
rect 3053 3547 3111 3553
rect 4132 3587 4190 3593
rect 4132 3553 4144 3587
rect 4178 3584 4190 3587
rect 4614 3584 4620 3596
rect 4178 3556 4620 3584
rect 4178 3553 4190 3556
rect 4132 3547 4190 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 5261 3587 5319 3593
rect 5261 3553 5273 3587
rect 5307 3584 5319 3587
rect 5350 3584 5356 3596
rect 5307 3556 5356 3584
rect 5307 3553 5319 3556
rect 5261 3547 5319 3553
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 7561 3587 7619 3593
rect 7561 3584 7573 3587
rect 7340 3556 7573 3584
rect 7340 3544 7346 3556
rect 7561 3553 7573 3556
rect 7607 3553 7619 3587
rect 7561 3547 7619 3553
rect 8662 3544 8668 3596
rect 8720 3584 8726 3596
rect 8757 3587 8815 3593
rect 8757 3584 8769 3587
rect 8720 3556 8769 3584
rect 8720 3544 8726 3556
rect 8757 3553 8769 3556
rect 8803 3553 8815 3587
rect 13538 3584 13544 3596
rect 13499 3556 13544 3584
rect 8757 3547 8815 3553
rect 13538 3544 13544 3556
rect 13596 3544 13602 3596
rect 17310 3584 17316 3596
rect 17271 3556 17316 3584
rect 17310 3544 17316 3556
rect 17368 3544 17374 3596
rect 3970 3476 3976 3528
rect 4028 3516 4034 3528
rect 6822 3516 6828 3528
rect 4028 3488 6828 3516
rect 4028 3476 4034 3488
rect 6822 3476 6828 3488
rect 6880 3516 6886 3528
rect 7009 3519 7067 3525
rect 7009 3516 7021 3519
rect 6880 3488 7021 3516
rect 6880 3476 6886 3488
rect 7009 3485 7021 3488
rect 7055 3485 7067 3519
rect 10042 3516 10048 3528
rect 10003 3488 10048 3516
rect 7009 3479 7067 3485
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 11974 3516 11980 3528
rect 11935 3488 11980 3516
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3516 15439 3519
rect 16114 3516 16120 3528
rect 15427 3488 16120 3516
rect 15427 3485 15439 3488
rect 15381 3479 15439 3485
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 16390 3516 16396 3528
rect 16303 3488 16396 3516
rect 16390 3476 16396 3488
rect 16448 3516 16454 3528
rect 18414 3516 18420 3528
rect 16448 3488 18420 3516
rect 16448 3476 16454 3488
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 10597 3451 10655 3457
rect 10597 3417 10609 3451
rect 10643 3417 10655 3451
rect 10597 3411 10655 3417
rect 1949 3383 2007 3389
rect 1949 3349 1961 3383
rect 1995 3380 2007 3383
rect 2498 3380 2504 3392
rect 1995 3352 2504 3380
rect 1995 3349 2007 3352
rect 1949 3343 2007 3349
rect 2498 3340 2504 3352
rect 2556 3340 2562 3392
rect 4203 3383 4261 3389
rect 4203 3349 4215 3383
rect 4249 3380 4261 3383
rect 4338 3380 4344 3392
rect 4249 3352 4344 3380
rect 4249 3349 4261 3352
rect 4203 3343 4261 3349
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 6454 3380 6460 3392
rect 6415 3352 6460 3380
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 10612 3380 10640 3411
rect 11146 3380 11152 3392
rect 10612 3352 11152 3380
rect 11146 3340 11152 3352
rect 11204 3380 11210 3392
rect 11333 3383 11391 3389
rect 11333 3380 11345 3383
rect 11204 3352 11345 3380
rect 11204 3340 11210 3352
rect 11333 3349 11345 3352
rect 11379 3349 11391 3383
rect 11333 3343 11391 3349
rect 1104 3290 22816 3312
rect 1104 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 12982 3290
rect 13034 3238 13046 3290
rect 13098 3238 13110 3290
rect 13162 3238 13174 3290
rect 13226 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 22816 3290
rect 1104 3216 22816 3238
rect 1394 3136 1400 3188
rect 1452 3176 1458 3188
rect 1535 3179 1593 3185
rect 1535 3176 1547 3179
rect 1452 3148 1547 3176
rect 1452 3136 1458 3148
rect 1535 3145 1547 3148
rect 1581 3145 1593 3179
rect 4154 3176 4160 3188
rect 1535 3139 1593 3145
rect 3436 3148 4160 3176
rect 1210 2932 1216 2984
rect 1268 2972 1274 2984
rect 1432 2975 1490 2981
rect 1432 2972 1444 2975
rect 1268 2944 1444 2972
rect 1268 2932 1274 2944
rect 1432 2941 1444 2944
rect 1478 2972 1490 2975
rect 1857 2975 1915 2981
rect 1857 2972 1869 2975
rect 1478 2944 1869 2972
rect 1478 2941 1490 2944
rect 1432 2935 1490 2941
rect 1857 2941 1869 2944
rect 1903 2941 1915 2975
rect 2498 2972 2504 2984
rect 2459 2944 2504 2972
rect 1857 2935 1915 2941
rect 2498 2932 2504 2944
rect 2556 2972 2562 2984
rect 3436 2981 3464 3148
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 5353 3179 5411 3185
rect 5353 3145 5365 3179
rect 5399 3176 5411 3179
rect 5442 3176 5448 3188
rect 5399 3148 5448 3176
rect 5399 3145 5411 3148
rect 5353 3139 5411 3145
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 5905 3179 5963 3185
rect 5905 3176 5917 3179
rect 5868 3148 5917 3176
rect 5868 3136 5874 3148
rect 5905 3145 5917 3148
rect 5951 3145 5963 3179
rect 5905 3139 5963 3145
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 7282 3176 7288 3188
rect 7239 3148 7288 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 8110 3176 8116 3188
rect 8071 3148 8116 3176
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9585 3179 9643 3185
rect 9585 3176 9597 3179
rect 9364 3148 9597 3176
rect 9364 3136 9370 3148
rect 9585 3145 9597 3148
rect 9631 3176 9643 3179
rect 9677 3179 9735 3185
rect 9677 3176 9689 3179
rect 9631 3148 9689 3176
rect 9631 3145 9643 3148
rect 9585 3139 9643 3145
rect 9677 3145 9689 3148
rect 9723 3145 9735 3179
rect 9677 3139 9735 3145
rect 11885 3179 11943 3185
rect 11885 3145 11897 3179
rect 11931 3176 11943 3179
rect 12066 3176 12072 3188
rect 11931 3148 12072 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 13538 3176 13544 3188
rect 13499 3148 13544 3176
rect 13538 3136 13544 3148
rect 13596 3136 13602 3188
rect 15746 3176 15752 3188
rect 15707 3148 15752 3176
rect 15746 3136 15752 3148
rect 15804 3136 15810 3188
rect 16114 3176 16120 3188
rect 16075 3148 16120 3176
rect 16114 3136 16120 3148
rect 16172 3176 16178 3188
rect 16945 3179 17003 3185
rect 16172 3148 16344 3176
rect 16172 3136 16178 3148
rect 4246 3068 4252 3120
rect 4304 3108 4310 3120
rect 7423 3111 7481 3117
rect 7423 3108 7435 3111
rect 4304 3080 7435 3108
rect 4304 3068 4310 3080
rect 7423 3077 7435 3080
rect 7469 3077 7481 3111
rect 7423 3071 7481 3077
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 10873 3111 10931 3117
rect 10873 3108 10885 3111
rect 9456 3080 10885 3108
rect 9456 3068 9462 3080
rect 10873 3077 10885 3080
rect 10919 3077 10931 3111
rect 10873 3071 10931 3077
rect 15197 3111 15255 3117
rect 15197 3077 15209 3111
rect 15243 3108 15255 3111
rect 16022 3108 16028 3120
rect 15243 3080 16028 3108
rect 15243 3077 15255 3080
rect 15197 3071 15255 3077
rect 4798 3040 4804 3052
rect 3896 3012 4804 3040
rect 3421 2975 3479 2981
rect 3421 2972 3433 2975
rect 2556 2944 3433 2972
rect 2556 2932 2562 2944
rect 3421 2941 3433 2944
rect 3467 2941 3479 2975
rect 3421 2935 3479 2941
rect 3142 2904 3148 2916
rect 3103 2876 3148 2904
rect 3142 2864 3148 2876
rect 3200 2864 3206 2916
rect 3510 2864 3516 2916
rect 3568 2904 3574 2916
rect 3896 2904 3924 3012
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 8389 3043 8447 3049
rect 8389 3009 8401 3043
rect 8435 3040 8447 3043
rect 8662 3040 8668 3052
rect 8435 3012 8668 3040
rect 8435 3009 8447 3012
rect 8389 3003 8447 3009
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 10042 3040 10048 3052
rect 9079 3012 10048 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 10042 3000 10048 3012
rect 10100 3040 10106 3052
rect 10229 3043 10287 3049
rect 10229 3040 10241 3043
rect 10100 3012 10241 3040
rect 10100 3000 10106 3012
rect 10229 3009 10241 3012
rect 10275 3040 10287 3043
rect 11241 3043 11299 3049
rect 11241 3040 11253 3043
rect 10275 3012 11253 3040
rect 10275 3009 10287 3012
rect 10229 3003 10287 3009
rect 11241 3009 11253 3012
rect 11287 3009 11299 3043
rect 11241 3003 11299 3009
rect 5696 2975 5754 2981
rect 5696 2941 5708 2975
rect 5742 2972 5754 2975
rect 7352 2975 7410 2981
rect 5742 2944 6224 2972
rect 5742 2941 5754 2944
rect 5696 2935 5754 2941
rect 4065 2907 4123 2913
rect 4065 2904 4077 2907
rect 3568 2876 4077 2904
rect 3568 2864 3574 2876
rect 4065 2873 4077 2876
rect 4111 2873 4123 2907
rect 4065 2867 4123 2873
rect 4154 2864 4160 2916
rect 4212 2904 4218 2916
rect 4706 2904 4712 2916
rect 4212 2876 4257 2904
rect 4667 2876 4712 2904
rect 4212 2864 4218 2876
rect 4706 2864 4712 2876
rect 4764 2864 4770 2916
rect 6196 2848 6224 2944
rect 7352 2941 7364 2975
rect 7398 2972 7410 2975
rect 9309 2975 9367 2981
rect 7398 2944 7880 2972
rect 7398 2941 7410 2944
rect 7352 2935 7410 2941
rect 7852 2848 7880 2944
rect 9309 2941 9321 2975
rect 9355 2972 9367 2975
rect 9490 2972 9496 2984
rect 9355 2944 9496 2972
rect 9355 2941 9367 2944
rect 9309 2935 9367 2941
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 10686 2932 10692 2984
rect 10744 2972 10750 2984
rect 15339 2981 15367 3080
rect 16022 3068 16028 3080
rect 16080 3068 16086 3120
rect 16316 3049 16344 3148
rect 16945 3145 16957 3179
rect 16991 3176 17003 3179
rect 17310 3176 17316 3188
rect 16991 3148 17316 3176
rect 16991 3145 17003 3148
rect 16945 3139 17003 3145
rect 17310 3136 17316 3148
rect 17368 3136 17374 3188
rect 18046 3136 18052 3188
rect 18104 3176 18110 3188
rect 18187 3179 18245 3185
rect 18187 3176 18199 3179
rect 18104 3148 18199 3176
rect 18104 3136 18110 3148
rect 18187 3145 18199 3148
rect 18233 3145 18245 3179
rect 18187 3139 18245 3145
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3009 16359 3043
rect 16301 3003 16359 3009
rect 12253 2975 12311 2981
rect 12253 2972 12265 2975
rect 10744 2944 12265 2972
rect 10744 2932 10750 2944
rect 12253 2941 12265 2944
rect 12299 2972 12311 2975
rect 12529 2975 12587 2981
rect 12529 2972 12541 2975
rect 12299 2944 12541 2972
rect 12299 2941 12311 2944
rect 12253 2935 12311 2941
rect 12529 2941 12541 2944
rect 12575 2941 12587 2975
rect 12529 2935 12587 2941
rect 14185 2975 14243 2981
rect 14185 2941 14197 2975
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 15324 2975 15382 2981
rect 15324 2941 15336 2975
rect 15370 2941 15382 2975
rect 15324 2935 15382 2941
rect 18116 2975 18174 2981
rect 18116 2941 18128 2975
rect 18162 2972 18174 2975
rect 18162 2944 18644 2972
rect 18162 2941 18174 2944
rect 18116 2935 18174 2941
rect 8478 2864 8484 2916
rect 8536 2904 8542 2916
rect 8536 2876 8581 2904
rect 8536 2864 8542 2876
rect 9398 2864 9404 2916
rect 9456 2904 9462 2916
rect 9953 2907 10011 2913
rect 9953 2904 9965 2907
rect 9456 2876 9965 2904
rect 9456 2864 9462 2876
rect 9953 2873 9965 2876
rect 9999 2873 10011 2907
rect 9953 2867 10011 2873
rect 10045 2907 10103 2913
rect 10045 2873 10057 2907
rect 10091 2873 10103 2907
rect 10045 2867 10103 2873
rect 2222 2836 2228 2848
rect 2183 2808 2228 2836
rect 2222 2796 2228 2808
rect 2280 2796 2286 2848
rect 3881 2839 3939 2845
rect 3881 2805 3893 2839
rect 3927 2836 3939 2839
rect 4614 2836 4620 2848
rect 3927 2808 4620 2836
rect 3927 2805 3939 2808
rect 3881 2799 3939 2805
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 6178 2836 6184 2848
rect 6139 2808 6184 2836
rect 6178 2796 6184 2808
rect 6236 2796 6242 2848
rect 7834 2836 7840 2848
rect 7795 2808 7840 2836
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 9585 2839 9643 2845
rect 9585 2805 9597 2839
rect 9631 2836 9643 2839
rect 10060 2836 10088 2867
rect 10778 2864 10784 2916
rect 10836 2904 10842 2916
rect 12437 2907 12495 2913
rect 12437 2904 12449 2907
rect 10836 2876 12449 2904
rect 10836 2864 10842 2876
rect 12437 2873 12449 2876
rect 12483 2873 12495 2907
rect 14200 2904 14228 2935
rect 14829 2907 14887 2913
rect 14829 2904 14841 2907
rect 14200 2876 14841 2904
rect 12437 2867 12495 2873
rect 14829 2873 14841 2876
rect 14875 2904 14887 2907
rect 15427 2907 15485 2913
rect 15427 2904 15439 2907
rect 14875 2876 15439 2904
rect 14875 2873 14887 2876
rect 14829 2867 14887 2873
rect 15427 2873 15439 2876
rect 15473 2873 15485 2907
rect 15427 2867 15485 2873
rect 18616 2848 18644 2944
rect 14366 2836 14372 2848
rect 9631 2808 10088 2836
rect 14327 2808 14372 2836
rect 9631 2805 9643 2808
rect 9585 2799 9643 2805
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 18598 2836 18604 2848
rect 18559 2808 18604 2836
rect 18598 2796 18604 2808
rect 18656 2796 18662 2848
rect 1104 2746 22816 2768
rect 1104 2694 8982 2746
rect 9034 2694 9046 2746
rect 9098 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 17174 2746
rect 17226 2694 22816 2746
rect 1104 2672 22816 2694
rect 3510 2632 3516 2644
rect 3471 2604 3516 2632
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 5350 2632 5356 2644
rect 5311 2604 5356 2632
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2632 5871 2635
rect 6454 2632 6460 2644
rect 5859 2604 6460 2632
rect 5859 2601 5871 2604
rect 5813 2595 5871 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 8389 2635 8447 2641
rect 6595 2604 7144 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 3142 2524 3148 2576
rect 3200 2564 3206 2576
rect 3789 2567 3847 2573
rect 3789 2564 3801 2567
rect 3200 2536 3801 2564
rect 3200 2524 3206 2536
rect 3789 2533 3801 2536
rect 3835 2564 3847 2567
rect 4433 2567 4491 2573
rect 4433 2564 4445 2567
rect 3835 2536 4445 2564
rect 3835 2533 3847 2536
rect 3789 2527 3847 2533
rect 4433 2533 4445 2536
rect 4479 2533 4491 2567
rect 4433 2527 4491 2533
rect 4706 2524 4712 2576
rect 4764 2564 4770 2576
rect 7116 2573 7144 2604
rect 8389 2601 8401 2635
rect 8435 2632 8447 2635
rect 8478 2632 8484 2644
rect 8435 2604 8484 2632
rect 8435 2601 8447 2604
rect 8389 2595 8447 2601
rect 8478 2592 8484 2604
rect 8536 2592 8542 2644
rect 11974 2632 11980 2644
rect 11935 2604 11980 2632
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 4985 2567 5043 2573
rect 4985 2564 4997 2567
rect 4764 2536 4997 2564
rect 4764 2524 4770 2536
rect 4985 2533 4997 2536
rect 5031 2564 5043 2567
rect 6273 2567 6331 2573
rect 6273 2564 6285 2567
rect 5031 2536 6285 2564
rect 5031 2533 5043 2536
rect 4985 2527 5043 2533
rect 6273 2533 6285 2536
rect 6319 2564 6331 2567
rect 7009 2567 7067 2573
rect 7009 2564 7021 2567
rect 6319 2536 7021 2564
rect 6319 2533 6331 2536
rect 6273 2527 6331 2533
rect 7009 2533 7021 2536
rect 7055 2533 7067 2567
rect 7009 2527 7067 2533
rect 7101 2567 7159 2573
rect 7101 2533 7113 2567
rect 7147 2533 7159 2567
rect 7101 2527 7159 2533
rect 10321 2567 10379 2573
rect 10321 2533 10333 2567
rect 10367 2564 10379 2567
rect 10597 2567 10655 2573
rect 10597 2564 10609 2567
rect 10367 2536 10609 2564
rect 10367 2533 10379 2536
rect 10321 2527 10379 2533
rect 10597 2533 10609 2536
rect 10643 2564 10655 2567
rect 10778 2564 10784 2576
rect 10643 2536 10784 2564
rect 10643 2533 10655 2536
rect 10597 2527 10655 2533
rect 10778 2524 10784 2536
rect 10836 2524 10842 2576
rect 11146 2564 11152 2576
rect 11107 2536 11152 2564
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 13998 2524 14004 2576
rect 14056 2564 14062 2576
rect 16025 2567 16083 2573
rect 16025 2564 16037 2567
rect 14056 2536 16037 2564
rect 14056 2524 14062 2536
rect 2222 2496 2228 2508
rect 1780 2468 2228 2496
rect 1026 2252 1032 2304
rect 1084 2292 1090 2304
rect 1780 2301 1808 2468
rect 2222 2456 2228 2468
rect 2280 2496 2286 2508
rect 2317 2499 2375 2505
rect 2317 2496 2329 2499
rect 2280 2468 2329 2496
rect 2280 2456 2286 2468
rect 2317 2465 2329 2468
rect 2363 2465 2375 2499
rect 2869 2499 2927 2505
rect 2869 2496 2881 2499
rect 2317 2459 2375 2465
rect 2608 2468 2881 2496
rect 1765 2295 1823 2301
rect 1765 2292 1777 2295
rect 1084 2264 1777 2292
rect 1084 2252 1090 2264
rect 1765 2261 1777 2264
rect 1811 2261 1823 2295
rect 2130 2292 2136 2304
rect 2091 2264 2136 2292
rect 1765 2255 1823 2261
rect 2130 2252 2136 2264
rect 2188 2292 2194 2304
rect 2608 2292 2636 2468
rect 2869 2465 2881 2468
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 6549 2499 6607 2505
rect 6549 2496 6561 2499
rect 6052 2468 6561 2496
rect 6052 2456 6058 2468
rect 6549 2465 6561 2468
rect 6595 2496 6607 2499
rect 6641 2499 6699 2505
rect 6641 2496 6653 2499
rect 6595 2468 6653 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 6641 2465 6653 2468
rect 6687 2465 6699 2499
rect 6641 2459 6699 2465
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12584 2468 12633 2496
rect 12584 2456 12590 2468
rect 12621 2465 12633 2468
rect 12667 2496 12679 2499
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12667 2468 13185 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 13630 2456 13636 2508
rect 13688 2496 13694 2508
rect 15488 2505 15516 2536
rect 16025 2533 16037 2536
rect 16071 2533 16083 2567
rect 16025 2527 16083 2533
rect 13725 2499 13783 2505
rect 13725 2496 13737 2499
rect 13688 2468 13737 2496
rect 13688 2456 13694 2468
rect 13725 2465 13737 2468
rect 13771 2496 13783 2499
rect 14277 2499 14335 2505
rect 14277 2496 14289 2499
rect 13771 2468 14289 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 14277 2465 14289 2468
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2465 15531 2499
rect 15473 2459 15531 2465
rect 16942 2456 16948 2508
rect 17000 2496 17006 2508
rect 17256 2499 17314 2505
rect 17256 2496 17268 2499
rect 17000 2468 17268 2496
rect 17000 2456 17006 2468
rect 17256 2465 17268 2468
rect 17302 2465 17314 2499
rect 17256 2459 17314 2465
rect 17359 2499 17417 2505
rect 17359 2465 17371 2499
rect 17405 2496 17417 2499
rect 18601 2499 18659 2505
rect 18601 2496 18613 2499
rect 17405 2468 18613 2496
rect 17405 2465 17417 2468
rect 17359 2459 17417 2465
rect 18601 2465 18613 2468
rect 18647 2496 18659 2499
rect 19153 2499 19211 2505
rect 19153 2496 19165 2499
rect 18647 2468 19165 2496
rect 18647 2465 18659 2468
rect 18601 2459 18659 2465
rect 19153 2465 19165 2468
rect 19199 2465 19211 2499
rect 19978 2496 19984 2508
rect 19939 2468 19984 2496
rect 19153 2459 19211 2465
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2428 2743 2431
rect 3970 2428 3976 2440
rect 2731 2400 3976 2428
rect 2731 2397 2743 2400
rect 2685 2391 2743 2397
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 4338 2428 4344 2440
rect 4299 2400 4344 2428
rect 4338 2388 4344 2400
rect 4396 2428 4402 2440
rect 5629 2431 5687 2437
rect 5629 2428 5641 2431
rect 4396 2400 5641 2428
rect 4396 2388 4402 2400
rect 5629 2397 5641 2400
rect 5675 2397 5687 2431
rect 7650 2428 7656 2440
rect 7611 2400 7656 2428
rect 5629 2391 5687 2397
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2428 8723 2431
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 8711 2400 9505 2428
rect 8711 2397 8723 2400
rect 8665 2391 8723 2397
rect 9493 2397 9505 2400
rect 9539 2428 9551 2431
rect 10505 2431 10563 2437
rect 10505 2428 10517 2431
rect 9539 2400 10517 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 10505 2397 10517 2400
rect 10551 2397 10563 2431
rect 17271 2428 17299 2459
rect 19978 2456 19984 2468
rect 20036 2496 20042 2508
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20036 2468 20545 2496
rect 20036 2456 20042 2468
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 17271 2400 17693 2428
rect 10505 2391 10563 2397
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 13262 2320 13268 2372
rect 13320 2360 13326 2372
rect 13909 2363 13967 2369
rect 13909 2360 13921 2363
rect 13320 2332 13921 2360
rect 13320 2320 13326 2332
rect 13909 2329 13921 2332
rect 13955 2329 13967 2363
rect 13909 2323 13967 2329
rect 12802 2292 12808 2304
rect 2188 2264 2636 2292
rect 12763 2264 12808 2292
rect 2188 2252 2194 2264
rect 12802 2252 12808 2264
rect 12860 2252 12866 2304
rect 15657 2295 15715 2301
rect 15657 2261 15669 2295
rect 15703 2292 15715 2295
rect 15930 2292 15936 2304
rect 15703 2264 15936 2292
rect 15703 2261 15715 2264
rect 15657 2255 15715 2261
rect 15930 2252 15936 2264
rect 15988 2252 15994 2304
rect 18785 2295 18843 2301
rect 18785 2261 18797 2295
rect 18831 2292 18843 2295
rect 20070 2292 20076 2304
rect 18831 2264 20076 2292
rect 18831 2261 18843 2264
rect 18785 2255 18843 2261
rect 20070 2252 20076 2264
rect 20128 2252 20134 2304
rect 20165 2295 20223 2301
rect 20165 2261 20177 2295
rect 20211 2292 20223 2295
rect 21542 2292 21548 2304
rect 20211 2264 21548 2292
rect 20211 2261 20223 2264
rect 20165 2255 20223 2261
rect 21542 2252 21548 2264
rect 21600 2252 21606 2304
rect 1104 2202 22816 2224
rect 1104 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 12982 2202
rect 13034 2150 13046 2202
rect 13098 2150 13110 2202
rect 13162 2150 13174 2202
rect 13226 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 22816 2202
rect 1104 2128 22816 2150
rect 8018 2048 8024 2100
rect 8076 2088 8082 2100
rect 13446 2088 13452 2100
rect 8076 2060 13452 2088
rect 8076 2048 8082 2060
rect 13446 2048 13452 2060
rect 13504 2048 13510 2100
rect 7834 1912 7840 1964
rect 7892 1952 7898 1964
rect 10226 1952 10232 1964
rect 7892 1924 10232 1952
rect 7892 1912 7898 1924
rect 10226 1912 10232 1924
rect 10284 1912 10290 1964
<< via1 >>
rect 20 23536 72 23588
rect 848 23536 900 23588
rect 4982 21734 5034 21786
rect 5046 21734 5098 21786
rect 5110 21734 5162 21786
rect 5174 21734 5226 21786
rect 12982 21734 13034 21786
rect 13046 21734 13098 21786
rect 13110 21734 13162 21786
rect 13174 21734 13226 21786
rect 20982 21734 21034 21786
rect 21046 21734 21098 21786
rect 21110 21734 21162 21786
rect 21174 21734 21226 21786
rect 8982 21190 9034 21242
rect 9046 21190 9098 21242
rect 9110 21190 9162 21242
rect 9174 21190 9226 21242
rect 16982 21190 17034 21242
rect 17046 21190 17098 21242
rect 17110 21190 17162 21242
rect 17174 21190 17226 21242
rect 112 20952 164 21004
rect 9956 20995 10008 21004
rect 9956 20961 10000 20995
rect 10000 20961 10008 20995
rect 9956 20952 10008 20961
rect 10232 20748 10284 20800
rect 4982 20646 5034 20698
rect 5046 20646 5098 20698
rect 5110 20646 5162 20698
rect 5174 20646 5226 20698
rect 12982 20646 13034 20698
rect 13046 20646 13098 20698
rect 13110 20646 13162 20698
rect 13174 20646 13226 20698
rect 20982 20646 21034 20698
rect 21046 20646 21098 20698
rect 21110 20646 21162 20698
rect 21174 20646 21226 20698
rect 4528 20587 4580 20596
rect 4528 20553 4537 20587
rect 4537 20553 4571 20587
rect 4571 20553 4580 20587
rect 4528 20544 4580 20553
rect 6092 20587 6144 20596
rect 6092 20553 6101 20587
rect 6101 20553 6135 20587
rect 6135 20553 6144 20587
rect 6092 20544 6144 20553
rect 7380 20587 7432 20596
rect 7380 20553 7389 20587
rect 7389 20553 7423 20587
rect 7423 20553 7432 20587
rect 7380 20544 7432 20553
rect 9312 20544 9364 20596
rect 9956 20587 10008 20596
rect 9956 20553 9965 20587
rect 9965 20553 9999 20587
rect 9999 20553 10008 20587
rect 9956 20544 10008 20553
rect 10968 20587 11020 20596
rect 10968 20553 10977 20587
rect 10977 20553 11011 20587
rect 11011 20553 11020 20587
rect 10968 20544 11020 20553
rect 1216 20340 1268 20392
rect 4528 20340 4580 20392
rect 6092 20340 6144 20392
rect 7380 20340 7432 20392
rect 10968 20340 11020 20392
rect 14280 20544 14332 20596
rect 15844 20544 15896 20596
rect 14556 20383 14608 20392
rect 14556 20349 14565 20383
rect 14565 20349 14599 20383
rect 14599 20349 14608 20383
rect 14556 20340 14608 20349
rect 17684 20544 17736 20596
rect 21272 20544 21324 20596
rect 21456 20587 21508 20596
rect 21456 20553 21465 20587
rect 21465 20553 21499 20587
rect 21499 20553 21508 20587
rect 21456 20544 21508 20553
rect 21456 20340 21508 20392
rect 1952 20204 2004 20256
rect 3792 20204 3844 20256
rect 6276 20204 6328 20256
rect 6644 20204 6696 20256
rect 9404 20247 9456 20256
rect 9404 20213 9413 20247
rect 9413 20213 9447 20247
rect 9447 20213 9456 20247
rect 9404 20204 9456 20213
rect 12532 20204 12584 20256
rect 13360 20204 13412 20256
rect 14924 20204 14976 20256
rect 17500 20204 17552 20256
rect 20628 20204 20680 20256
rect 8982 20102 9034 20154
rect 9046 20102 9098 20154
rect 9110 20102 9162 20154
rect 9174 20102 9226 20154
rect 16982 20102 17034 20154
rect 17046 20102 17098 20154
rect 17110 20102 17162 20154
rect 17174 20102 17226 20154
rect 1584 20043 1636 20052
rect 1584 20009 1593 20043
rect 1593 20009 1627 20043
rect 1627 20009 1636 20043
rect 1584 20000 1636 20009
rect 9404 20000 9456 20052
rect 10232 19932 10284 19984
rect 11336 19932 11388 19984
rect 12624 19975 12676 19984
rect 12624 19941 12633 19975
rect 12633 19941 12667 19975
rect 12667 19941 12676 19975
rect 12624 19932 12676 19941
rect 1308 19864 1360 19916
rect 2780 19864 2832 19916
rect 5632 19864 5684 19916
rect 10048 19864 10100 19916
rect 18696 19864 18748 19916
rect 12532 19839 12584 19848
rect 12532 19805 12541 19839
rect 12541 19805 12575 19839
rect 12575 19805 12584 19839
rect 12532 19796 12584 19805
rect 12716 19796 12768 19848
rect 3424 19660 3476 19712
rect 6460 19703 6512 19712
rect 6460 19669 6469 19703
rect 6469 19669 6503 19703
rect 6503 19669 6512 19703
rect 6460 19660 6512 19669
rect 10048 19660 10100 19712
rect 17868 19660 17920 19712
rect 4982 19558 5034 19610
rect 5046 19558 5098 19610
rect 5110 19558 5162 19610
rect 5174 19558 5226 19610
rect 12982 19558 13034 19610
rect 13046 19558 13098 19610
rect 13110 19558 13162 19610
rect 13174 19558 13226 19610
rect 20982 19558 21034 19610
rect 21046 19558 21098 19610
rect 21110 19558 21162 19610
rect 21174 19558 21226 19610
rect 2780 19456 2832 19508
rect 6460 19456 6512 19508
rect 10232 19499 10284 19508
rect 10232 19465 10241 19499
rect 10241 19465 10275 19499
rect 10275 19465 10284 19499
rect 10232 19456 10284 19465
rect 12532 19456 12584 19508
rect 12808 19456 12860 19508
rect 1584 19431 1636 19440
rect 1584 19397 1593 19431
rect 1593 19397 1627 19431
rect 1627 19397 1636 19431
rect 1584 19388 1636 19397
rect 12624 19320 12676 19372
rect 9496 19295 9548 19304
rect 9496 19261 9505 19295
rect 9505 19261 9539 19295
rect 9539 19261 9548 19295
rect 9496 19252 9548 19261
rect 11336 19295 11388 19304
rect 11336 19261 11345 19295
rect 11345 19261 11379 19295
rect 11379 19261 11388 19295
rect 11336 19252 11388 19261
rect 12808 19252 12860 19304
rect 19432 19456 19484 19508
rect 7564 19227 7616 19236
rect 1308 19116 1360 19168
rect 2044 19116 2096 19168
rect 5632 19159 5684 19168
rect 5632 19125 5641 19159
rect 5641 19125 5675 19159
rect 5675 19125 5684 19159
rect 5632 19116 5684 19125
rect 6460 19116 6512 19168
rect 7564 19193 7573 19227
rect 7573 19193 7607 19227
rect 7607 19193 7616 19227
rect 7564 19184 7616 19193
rect 9772 19227 9824 19236
rect 9772 19193 9781 19227
rect 9781 19193 9815 19227
rect 9815 19193 9824 19227
rect 9772 19184 9824 19193
rect 18696 19227 18748 19236
rect 18696 19193 18705 19227
rect 18705 19193 18739 19227
rect 18739 19193 18748 19227
rect 18696 19184 18748 19193
rect 22836 19184 22888 19236
rect 12440 19116 12492 19168
rect 12808 19116 12860 19168
rect 8982 19014 9034 19066
rect 9046 19014 9098 19066
rect 9110 19014 9162 19066
rect 9174 19014 9226 19066
rect 16982 19014 17034 19066
rect 17046 19014 17098 19066
rect 17110 19014 17162 19066
rect 17174 19014 17226 19066
rect 112 18912 164 18964
rect 2044 18955 2096 18964
rect 2044 18921 2053 18955
rect 2053 18921 2087 18955
rect 2087 18921 2096 18955
rect 2044 18912 2096 18921
rect 12440 18955 12492 18964
rect 12440 18921 12449 18955
rect 12449 18921 12483 18955
rect 12483 18921 12492 18955
rect 12440 18912 12492 18921
rect 6736 18887 6788 18896
rect 6736 18853 6745 18887
rect 6745 18853 6779 18887
rect 6779 18853 6788 18887
rect 6736 18844 6788 18853
rect 9772 18844 9824 18896
rect 12900 18887 12952 18896
rect 12900 18853 12909 18887
rect 12909 18853 12943 18887
rect 12943 18853 12952 18887
rect 12900 18844 12952 18853
rect 2596 18776 2648 18828
rect 4344 18819 4396 18828
rect 4344 18785 4353 18819
rect 4353 18785 4387 18819
rect 4387 18785 4396 18819
rect 4344 18776 4396 18785
rect 21272 18776 21324 18828
rect 3516 18708 3568 18760
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 6920 18751 6972 18760
rect 6920 18717 6929 18751
rect 6929 18717 6963 18751
rect 6963 18717 6972 18751
rect 6920 18708 6972 18717
rect 9128 18708 9180 18760
rect 10048 18751 10100 18760
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 11888 18708 11940 18760
rect 12808 18751 12860 18760
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 13268 18751 13320 18760
rect 13268 18717 13277 18751
rect 13277 18717 13311 18751
rect 13311 18717 13320 18751
rect 13268 18708 13320 18717
rect 4804 18640 4856 18692
rect 8760 18572 8812 18624
rect 9404 18615 9456 18624
rect 9404 18581 9413 18615
rect 9413 18581 9447 18615
rect 9447 18581 9456 18615
rect 9404 18572 9456 18581
rect 11336 18572 11388 18624
rect 16396 18572 16448 18624
rect 4982 18470 5034 18522
rect 5046 18470 5098 18522
rect 5110 18470 5162 18522
rect 5174 18470 5226 18522
rect 12982 18470 13034 18522
rect 13046 18470 13098 18522
rect 13110 18470 13162 18522
rect 13174 18470 13226 18522
rect 20982 18470 21034 18522
rect 21046 18470 21098 18522
rect 21110 18470 21162 18522
rect 21174 18470 21226 18522
rect 4344 18411 4396 18420
rect 4344 18377 4353 18411
rect 4353 18377 4387 18411
rect 4387 18377 4396 18411
rect 4344 18368 4396 18377
rect 4804 18368 4856 18420
rect 6736 18368 6788 18420
rect 9128 18411 9180 18420
rect 9128 18377 9137 18411
rect 9137 18377 9171 18411
rect 9171 18377 9180 18411
rect 9128 18368 9180 18377
rect 9772 18368 9824 18420
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 21272 18368 21324 18420
rect 2504 18300 2556 18352
rect 2044 18232 2096 18284
rect 3424 18275 3476 18284
rect 3424 18241 3433 18275
rect 3433 18241 3467 18275
rect 3467 18241 3476 18275
rect 3424 18232 3476 18241
rect 12440 18300 12492 18352
rect 6644 18232 6696 18284
rect 6920 18275 6972 18284
rect 6920 18241 6929 18275
rect 6929 18241 6963 18275
rect 6963 18241 6972 18275
rect 6920 18232 6972 18241
rect 7564 18275 7616 18284
rect 7564 18241 7573 18275
rect 7573 18241 7607 18275
rect 7607 18241 7616 18275
rect 7564 18232 7616 18241
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 10048 18275 10100 18284
rect 10048 18241 10057 18275
rect 10057 18241 10091 18275
rect 10091 18241 10100 18275
rect 10048 18232 10100 18241
rect 13268 18232 13320 18284
rect 1676 18028 1728 18080
rect 2504 18096 2556 18148
rect 3516 18139 3568 18148
rect 3516 18105 3525 18139
rect 3525 18105 3559 18139
rect 3559 18105 3568 18139
rect 4068 18139 4120 18148
rect 3516 18096 3568 18105
rect 4068 18105 4077 18139
rect 4077 18105 4111 18139
rect 4111 18105 4120 18139
rect 4068 18096 4120 18105
rect 5632 18096 5684 18148
rect 7012 18139 7064 18148
rect 7012 18105 7021 18139
rect 7021 18105 7055 18139
rect 7055 18105 7064 18139
rect 7012 18096 7064 18105
rect 9496 18139 9548 18148
rect 9496 18105 9505 18139
rect 9505 18105 9539 18139
rect 9539 18105 9548 18139
rect 9496 18096 9548 18105
rect 2136 18028 2188 18080
rect 2596 18028 2648 18080
rect 12256 18071 12308 18080
rect 12256 18037 12265 18071
rect 12265 18037 12299 18071
rect 12299 18037 12308 18071
rect 12256 18028 12308 18037
rect 12900 18028 12952 18080
rect 8982 17926 9034 17978
rect 9046 17926 9098 17978
rect 9110 17926 9162 17978
rect 9174 17926 9226 17978
rect 16982 17926 17034 17978
rect 17046 17926 17098 17978
rect 17110 17926 17162 17978
rect 17174 17926 17226 17978
rect 3424 17867 3476 17876
rect 3424 17833 3433 17867
rect 3433 17833 3467 17867
rect 3467 17833 3476 17867
rect 3424 17824 3476 17833
rect 6920 17824 6972 17876
rect 2320 17799 2372 17808
rect 2320 17765 2329 17799
rect 2329 17765 2363 17799
rect 2363 17765 2372 17799
rect 2320 17756 2372 17765
rect 4344 17756 4396 17808
rect 6460 17799 6512 17808
rect 6460 17765 6469 17799
rect 6469 17765 6503 17799
rect 6503 17765 6512 17799
rect 6460 17756 6512 17765
rect 8760 17867 8812 17876
rect 8760 17833 8769 17867
rect 8769 17833 8803 17867
rect 8803 17833 8812 17867
rect 8760 17824 8812 17833
rect 9772 17756 9824 17808
rect 12256 17799 12308 17808
rect 12256 17765 12265 17799
rect 12265 17765 12299 17799
rect 12299 17765 12308 17799
rect 12256 17756 12308 17765
rect 12900 17731 12952 17740
rect 12900 17697 12909 17731
rect 12909 17697 12943 17731
rect 12943 17697 12952 17731
rect 12900 17688 12952 17697
rect 2504 17663 2556 17672
rect 2504 17629 2513 17663
rect 2513 17629 2547 17663
rect 2547 17629 2556 17663
rect 2504 17620 2556 17629
rect 4252 17620 4304 17672
rect 4068 17552 4120 17604
rect 5908 17620 5960 17672
rect 9864 17620 9916 17672
rect 9404 17552 9456 17604
rect 13728 17620 13780 17672
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 9496 17484 9548 17536
rect 11244 17484 11296 17536
rect 4982 17382 5034 17434
rect 5046 17382 5098 17434
rect 5110 17382 5162 17434
rect 5174 17382 5226 17434
rect 12982 17382 13034 17434
rect 13046 17382 13098 17434
rect 13110 17382 13162 17434
rect 13174 17382 13226 17434
rect 20982 17382 21034 17434
rect 21046 17382 21098 17434
rect 21110 17382 21162 17434
rect 21174 17382 21226 17434
rect 4344 17280 4396 17332
rect 12808 17280 12860 17332
rect 8760 17212 8812 17264
rect 9404 17255 9456 17264
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 4160 17144 4212 17196
rect 6460 17144 6512 17196
rect 9404 17221 9413 17255
rect 9413 17221 9447 17255
rect 9447 17221 9456 17255
rect 9404 17212 9456 17221
rect 9864 17144 9916 17196
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 13268 17144 13320 17196
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 2320 17076 2372 17128
rect 6736 17076 6788 17128
rect 2044 16940 2096 16992
rect 4252 16940 4304 16992
rect 5908 16983 5960 16992
rect 5908 16949 5917 16983
rect 5917 16949 5951 16983
rect 5951 16949 5960 16983
rect 5908 16940 5960 16949
rect 9312 17008 9364 17060
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 10140 16940 10192 16992
rect 10692 17008 10744 17060
rect 11520 17051 11572 17060
rect 11520 17017 11529 17051
rect 11529 17017 11563 17051
rect 11563 17017 11572 17051
rect 11520 17008 11572 17017
rect 13636 17051 13688 17060
rect 12992 16940 13044 16992
rect 13636 17017 13645 17051
rect 13645 17017 13679 17051
rect 13679 17017 13688 17051
rect 13636 17008 13688 17017
rect 13268 16940 13320 16992
rect 14464 17051 14516 17060
rect 14464 17017 14473 17051
rect 14473 17017 14507 17051
rect 14507 17017 14516 17051
rect 14464 17008 14516 17017
rect 8982 16838 9034 16890
rect 9046 16838 9098 16890
rect 9110 16838 9162 16890
rect 9174 16838 9226 16890
rect 16982 16838 17034 16890
rect 17046 16838 17098 16890
rect 17110 16838 17162 16890
rect 17174 16838 17226 16890
rect 1768 16779 1820 16788
rect 1768 16745 1777 16779
rect 1777 16745 1811 16779
rect 1811 16745 1820 16779
rect 1768 16736 1820 16745
rect 2872 16736 2924 16788
rect 6368 16779 6420 16788
rect 6368 16745 6377 16779
rect 6377 16745 6411 16779
rect 6411 16745 6420 16779
rect 6368 16736 6420 16745
rect 6736 16736 6788 16788
rect 2044 16668 2096 16720
rect 4068 16668 4120 16720
rect 3884 16600 3936 16652
rect 4712 16600 4764 16652
rect 5448 16600 5500 16652
rect 8116 16600 8168 16652
rect 10140 16736 10192 16788
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 12808 16736 12860 16788
rect 12992 16779 13044 16788
rect 12992 16745 13001 16779
rect 13001 16745 13035 16779
rect 13035 16745 13044 16779
rect 12992 16736 13044 16745
rect 9312 16668 9364 16720
rect 13452 16711 13504 16720
rect 13452 16677 13461 16711
rect 13461 16677 13495 16711
rect 13495 16677 13504 16711
rect 13452 16668 13504 16677
rect 14464 16668 14516 16720
rect 8668 16600 8720 16652
rect 9496 16600 9548 16652
rect 9772 16643 9824 16652
rect 9772 16609 9781 16643
rect 9781 16609 9815 16643
rect 9815 16609 9824 16643
rect 9772 16600 9824 16609
rect 15384 16600 15436 16652
rect 2872 16532 2924 16584
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 11520 16575 11572 16584
rect 11520 16541 11529 16575
rect 11529 16541 11563 16575
rect 11563 16541 11572 16575
rect 11520 16532 11572 16541
rect 13636 16575 13688 16584
rect 13636 16541 13645 16575
rect 13645 16541 13679 16575
rect 13679 16541 13688 16575
rect 13636 16532 13688 16541
rect 13728 16464 13780 16516
rect 4160 16396 4212 16448
rect 5816 16439 5868 16448
rect 5816 16405 5825 16439
rect 5825 16405 5859 16439
rect 5859 16405 5868 16439
rect 5816 16396 5868 16405
rect 10692 16396 10744 16448
rect 14464 16396 14516 16448
rect 4982 16294 5034 16346
rect 5046 16294 5098 16346
rect 5110 16294 5162 16346
rect 5174 16294 5226 16346
rect 12982 16294 13034 16346
rect 13046 16294 13098 16346
rect 13110 16294 13162 16346
rect 13174 16294 13226 16346
rect 20982 16294 21034 16346
rect 21046 16294 21098 16346
rect 21110 16294 21162 16346
rect 21174 16294 21226 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 2872 16192 2924 16244
rect 8116 16235 8168 16244
rect 8116 16201 8125 16235
rect 8125 16201 8159 16235
rect 8159 16201 8168 16235
rect 8116 16192 8168 16201
rect 11244 16235 11296 16244
rect 11244 16201 11253 16235
rect 11253 16201 11287 16235
rect 11287 16201 11296 16235
rect 11244 16192 11296 16201
rect 13452 16192 13504 16244
rect 13728 16192 13780 16244
rect 15384 16235 15436 16244
rect 15384 16201 15393 16235
rect 15393 16201 15427 16235
rect 15427 16201 15436 16235
rect 15384 16192 15436 16201
rect 13268 16124 13320 16176
rect 5816 16099 5868 16108
rect 5816 16065 5825 16099
rect 5825 16065 5859 16099
rect 5859 16065 5868 16099
rect 5816 16056 5868 16065
rect 6644 16056 6696 16108
rect 8576 16099 8628 16108
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 3608 16031 3660 16040
rect 3608 15997 3617 16031
rect 3617 15997 3651 16031
rect 3651 15997 3660 16031
rect 3608 15988 3660 15997
rect 4344 15988 4396 16040
rect 5448 16031 5500 16040
rect 5448 15997 5457 16031
rect 5457 15997 5491 16031
rect 5491 15997 5500 16031
rect 5448 15988 5500 15997
rect 7288 16031 7340 16040
rect 2964 15963 3016 15972
rect 2964 15929 2973 15963
rect 2973 15929 3007 15963
rect 3007 15929 3016 15963
rect 2964 15920 3016 15929
rect 5264 15920 5316 15972
rect 7288 15997 7297 16031
rect 7297 15997 7331 16031
rect 7331 15997 7340 16031
rect 7288 15988 7340 15997
rect 8576 16065 8585 16099
rect 8585 16065 8619 16099
rect 8619 16065 8628 16099
rect 8576 16056 8628 16065
rect 8668 15988 8720 16040
rect 10324 16031 10376 16040
rect 10324 15997 10333 16031
rect 10333 15997 10367 16031
rect 10367 15997 10376 16031
rect 10324 15988 10376 15997
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 13636 15988 13688 16040
rect 10232 15920 10284 15972
rect 11888 15920 11940 15972
rect 12072 15920 12124 15972
rect 2044 15895 2096 15904
rect 2044 15861 2053 15895
rect 2053 15861 2087 15895
rect 2087 15861 2096 15895
rect 2044 15852 2096 15861
rect 3884 15852 3936 15904
rect 4712 15852 4764 15904
rect 6368 15852 6420 15904
rect 6460 15895 6512 15904
rect 6460 15861 6469 15895
rect 6469 15861 6503 15895
rect 6503 15861 6512 15895
rect 6460 15852 6512 15861
rect 6920 15895 6972 15904
rect 6920 15861 6929 15895
rect 6929 15861 6963 15895
rect 6963 15861 6972 15895
rect 6920 15852 6972 15861
rect 9496 15895 9548 15904
rect 9496 15861 9505 15895
rect 9505 15861 9539 15895
rect 9539 15861 9548 15895
rect 9496 15852 9548 15861
rect 13636 15852 13688 15904
rect 8982 15750 9034 15802
rect 9046 15750 9098 15802
rect 9110 15750 9162 15802
rect 9174 15750 9226 15802
rect 16982 15750 17034 15802
rect 17046 15750 17098 15802
rect 17110 15750 17162 15802
rect 17174 15750 17226 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 4160 15691 4212 15700
rect 4160 15657 4169 15691
rect 4169 15657 4203 15691
rect 4203 15657 4212 15691
rect 5264 15691 5316 15700
rect 4160 15648 4212 15657
rect 5264 15657 5273 15691
rect 5273 15657 5307 15691
rect 5307 15657 5316 15691
rect 5264 15648 5316 15657
rect 7012 15648 7064 15700
rect 8576 15648 8628 15700
rect 9496 15648 9548 15700
rect 11520 15648 11572 15700
rect 13360 15648 13412 15700
rect 14280 15648 14332 15700
rect 2964 15580 3016 15632
rect 6368 15580 6420 15632
rect 10324 15623 10376 15632
rect 10324 15589 10333 15623
rect 10333 15589 10367 15623
rect 10367 15589 10376 15623
rect 10324 15580 10376 15589
rect 12440 15580 12492 15632
rect 13728 15580 13780 15632
rect 4344 15555 4396 15564
rect 4344 15521 4353 15555
rect 4353 15521 4387 15555
rect 4387 15521 4396 15555
rect 4344 15512 4396 15521
rect 4712 15512 4764 15564
rect 5448 15512 5500 15564
rect 6920 15512 6972 15564
rect 8024 15555 8076 15564
rect 8024 15521 8033 15555
rect 8033 15521 8067 15555
rect 8067 15521 8076 15555
rect 8024 15512 8076 15521
rect 8668 15512 8720 15564
rect 10876 15555 10928 15564
rect 10876 15521 10885 15555
rect 10885 15521 10919 15555
rect 10919 15521 10928 15555
rect 10876 15512 10928 15521
rect 2688 15444 2740 15496
rect 3240 15444 3292 15496
rect 4620 15444 4672 15496
rect 6736 15376 6788 15428
rect 7288 15376 7340 15428
rect 14464 15444 14516 15496
rect 13452 15376 13504 15428
rect 1400 15308 1452 15360
rect 3516 15308 3568 15360
rect 10692 15351 10744 15360
rect 10692 15317 10701 15351
rect 10701 15317 10735 15351
rect 10735 15317 10744 15351
rect 10692 15308 10744 15317
rect 12348 15308 12400 15360
rect 4982 15206 5034 15258
rect 5046 15206 5098 15258
rect 5110 15206 5162 15258
rect 5174 15206 5226 15258
rect 12982 15206 13034 15258
rect 13046 15206 13098 15258
rect 13110 15206 13162 15258
rect 13174 15206 13226 15258
rect 20982 15206 21034 15258
rect 21046 15206 21098 15258
rect 21110 15206 21162 15258
rect 21174 15206 21226 15258
rect 2964 15104 3016 15156
rect 3700 15104 3752 15156
rect 4344 15104 4396 15156
rect 4712 15104 4764 15156
rect 5448 15147 5500 15156
rect 5448 15113 5457 15147
rect 5457 15113 5491 15147
rect 5491 15113 5500 15147
rect 5448 15104 5500 15113
rect 10232 15147 10284 15156
rect 10232 15113 10241 15147
rect 10241 15113 10275 15147
rect 10275 15113 10284 15147
rect 10232 15104 10284 15113
rect 11336 15147 11388 15156
rect 11336 15113 11345 15147
rect 11345 15113 11379 15147
rect 11379 15113 11388 15147
rect 11336 15104 11388 15113
rect 12072 15104 12124 15156
rect 13728 15147 13780 15156
rect 13728 15113 13737 15147
rect 13737 15113 13771 15147
rect 13771 15113 13780 15147
rect 13728 15104 13780 15113
rect 4620 15079 4672 15088
rect 4620 15045 4629 15079
rect 4629 15045 4663 15079
rect 4663 15045 4672 15079
rect 4620 15036 4672 15045
rect 13452 15036 13504 15088
rect 1952 14968 2004 15020
rect 2320 15011 2372 15020
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4068 14968 4120 14977
rect 4252 14968 4304 15020
rect 14280 15011 14332 15020
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 6000 14943 6052 14952
rect 6000 14909 6009 14943
rect 6009 14909 6043 14943
rect 6043 14909 6052 14943
rect 6000 14900 6052 14909
rect 10324 14900 10376 14952
rect 12348 14900 12400 14952
rect 18512 14900 18564 14952
rect 2596 14832 2648 14884
rect 3608 14832 3660 14884
rect 10232 14832 10284 14884
rect 10876 14832 10928 14884
rect 12072 14832 12124 14884
rect 4988 14807 5040 14816
rect 4988 14773 4997 14807
rect 4997 14773 5031 14807
rect 5031 14773 5040 14807
rect 4988 14764 5040 14773
rect 6368 14807 6420 14816
rect 6368 14773 6377 14807
rect 6377 14773 6411 14807
rect 6411 14773 6420 14807
rect 6368 14764 6420 14773
rect 6460 14764 6512 14816
rect 8024 14807 8076 14816
rect 8024 14773 8033 14807
rect 8033 14773 8067 14807
rect 8067 14773 8076 14807
rect 8024 14764 8076 14773
rect 8668 14764 8720 14816
rect 14096 14807 14148 14816
rect 14096 14773 14105 14807
rect 14105 14773 14139 14807
rect 14139 14773 14148 14807
rect 14096 14764 14148 14773
rect 19708 14764 19760 14816
rect 8982 14662 9034 14714
rect 9046 14662 9098 14714
rect 9110 14662 9162 14714
rect 9174 14662 9226 14714
rect 16982 14662 17034 14714
rect 17046 14662 17098 14714
rect 17110 14662 17162 14714
rect 17174 14662 17226 14714
rect 2688 14603 2740 14612
rect 2688 14569 2697 14603
rect 2697 14569 2731 14603
rect 2731 14569 2740 14603
rect 2688 14560 2740 14569
rect 1860 14535 1912 14544
rect 1860 14501 1869 14535
rect 1869 14501 1903 14535
rect 1903 14501 1912 14535
rect 1860 14492 1912 14501
rect 4252 14560 4304 14612
rect 4344 14560 4396 14612
rect 4988 14603 5040 14612
rect 4988 14569 4997 14603
rect 4997 14569 5031 14603
rect 5031 14569 5040 14603
rect 4988 14560 5040 14569
rect 10324 14603 10376 14612
rect 10324 14569 10333 14603
rect 10333 14569 10367 14603
rect 10367 14569 10376 14603
rect 10324 14560 10376 14569
rect 14464 14603 14516 14612
rect 14464 14569 14473 14603
rect 14473 14569 14507 14603
rect 14507 14569 14516 14603
rect 14464 14560 14516 14569
rect 19892 14603 19944 14612
rect 19892 14569 19901 14603
rect 19901 14569 19935 14603
rect 19935 14569 19944 14603
rect 19892 14560 19944 14569
rect 4068 14492 4120 14544
rect 6368 14492 6420 14544
rect 12348 14535 12400 14544
rect 12348 14501 12357 14535
rect 12357 14501 12391 14535
rect 12391 14501 12400 14535
rect 12348 14492 12400 14501
rect 14096 14535 14148 14544
rect 14096 14501 14105 14535
rect 14105 14501 14139 14535
rect 14139 14501 14148 14535
rect 14096 14492 14148 14501
rect 16764 14535 16816 14544
rect 16764 14501 16773 14535
rect 16773 14501 16807 14535
rect 16807 14501 16816 14535
rect 16764 14492 16816 14501
rect 10140 14467 10192 14476
rect 10140 14433 10149 14467
rect 10149 14433 10183 14467
rect 10183 14433 10192 14467
rect 10140 14424 10192 14433
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 5908 14399 5960 14408
rect 5908 14365 5917 14399
rect 5917 14365 5951 14399
rect 5951 14365 5960 14399
rect 5908 14356 5960 14365
rect 8116 14356 8168 14408
rect 10232 14356 10284 14408
rect 11888 14467 11940 14476
rect 11888 14433 11897 14467
rect 11897 14433 11931 14467
rect 11931 14433 11940 14467
rect 11888 14424 11940 14433
rect 12164 14467 12216 14476
rect 12164 14433 12173 14467
rect 12173 14433 12207 14467
rect 12207 14433 12216 14467
rect 12164 14424 12216 14433
rect 13728 14467 13780 14476
rect 13728 14433 13737 14467
rect 13737 14433 13771 14467
rect 13771 14433 13780 14467
rect 13728 14424 13780 14433
rect 18788 14467 18840 14476
rect 18788 14433 18797 14467
rect 18797 14433 18831 14467
rect 18831 14433 18840 14467
rect 18788 14424 18840 14433
rect 19708 14467 19760 14476
rect 19708 14433 19717 14467
rect 19717 14433 19751 14467
rect 19751 14433 19760 14467
rect 19708 14424 19760 14433
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 17316 14399 17368 14408
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 2320 14331 2372 14340
rect 2320 14297 2329 14331
rect 2329 14297 2363 14331
rect 2363 14297 2372 14331
rect 2320 14288 2372 14297
rect 2596 14288 2648 14340
rect 10784 14288 10836 14340
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 12808 14263 12860 14272
rect 12808 14229 12817 14263
rect 12817 14229 12851 14263
rect 12851 14229 12860 14263
rect 12808 14220 12860 14229
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 18420 14263 18472 14272
rect 18420 14229 18429 14263
rect 18429 14229 18463 14263
rect 18463 14229 18472 14263
rect 18420 14220 18472 14229
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 12982 14118 13034 14170
rect 13046 14118 13098 14170
rect 13110 14118 13162 14170
rect 13174 14118 13226 14170
rect 20982 14118 21034 14170
rect 21046 14118 21098 14170
rect 21110 14118 21162 14170
rect 21174 14118 21226 14170
rect 1860 14059 1912 14068
rect 1860 14025 1869 14059
rect 1869 14025 1903 14059
rect 1903 14025 1912 14059
rect 1860 14016 1912 14025
rect 2596 14059 2648 14068
rect 2596 14025 2605 14059
rect 2605 14025 2639 14059
rect 2639 14025 2648 14059
rect 2596 14016 2648 14025
rect 3700 14059 3752 14068
rect 3700 14025 3709 14059
rect 3709 14025 3743 14059
rect 3743 14025 3752 14059
rect 3700 14016 3752 14025
rect 5908 14016 5960 14068
rect 11060 14059 11112 14068
rect 11060 14025 11069 14059
rect 11069 14025 11103 14059
rect 11103 14025 11112 14059
rect 11060 14016 11112 14025
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 13728 14059 13780 14068
rect 13728 14025 13737 14059
rect 13737 14025 13771 14059
rect 13771 14025 13780 14059
rect 13728 14016 13780 14025
rect 16764 14059 16816 14068
rect 16764 14025 16773 14059
rect 16773 14025 16807 14059
rect 16807 14025 16816 14059
rect 16764 14016 16816 14025
rect 18052 14016 18104 14068
rect 18788 14016 18840 14068
rect 19708 14016 19760 14068
rect 2688 13948 2740 14000
rect 10140 13948 10192 14000
rect 16672 13948 16724 14000
rect 2320 13880 2372 13932
rect 9312 13923 9364 13932
rect 9312 13889 9321 13923
rect 9321 13889 9355 13923
rect 9355 13889 9364 13923
rect 9312 13880 9364 13889
rect 11152 13923 11204 13932
rect 11152 13889 11161 13923
rect 11161 13889 11195 13923
rect 11195 13889 11204 13923
rect 11152 13880 11204 13889
rect 11888 13923 11940 13932
rect 11888 13889 11897 13923
rect 11897 13889 11931 13923
rect 11931 13889 11940 13923
rect 11888 13880 11940 13889
rect 15200 13880 15252 13932
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 2596 13812 2648 13864
rect 3700 13812 3752 13864
rect 4528 13812 4580 13864
rect 5724 13812 5776 13864
rect 7472 13855 7524 13864
rect 7472 13821 7481 13855
rect 7481 13821 7515 13855
rect 7515 13821 7524 13855
rect 7472 13812 7524 13821
rect 10784 13855 10836 13864
rect 10784 13821 10793 13855
rect 10793 13821 10827 13855
rect 10827 13821 10836 13855
rect 10784 13812 10836 13821
rect 11520 13812 11572 13864
rect 12808 13855 12860 13864
rect 12808 13821 12817 13855
rect 12817 13821 12851 13855
rect 12851 13821 12860 13855
rect 12808 13812 12860 13821
rect 2044 13744 2096 13796
rect 3976 13744 4028 13796
rect 4068 13719 4120 13728
rect 4068 13685 4077 13719
rect 4077 13685 4111 13719
rect 4111 13685 4120 13719
rect 4068 13676 4120 13685
rect 4160 13676 4212 13728
rect 4344 13676 4396 13728
rect 6368 13676 6420 13728
rect 7932 13676 7984 13728
rect 9956 13787 10008 13796
rect 9956 13753 9965 13787
rect 9965 13753 9999 13787
rect 9999 13753 10008 13787
rect 9956 13744 10008 13753
rect 10232 13676 10284 13728
rect 10600 13676 10652 13728
rect 14740 13744 14792 13796
rect 13268 13676 13320 13728
rect 15936 13676 15988 13728
rect 17408 13676 17460 13728
rect 18420 13744 18472 13796
rect 18512 13744 18564 13796
rect 18788 13787 18840 13796
rect 18788 13753 18797 13787
rect 18797 13753 18831 13787
rect 18831 13753 18840 13787
rect 18788 13744 18840 13753
rect 8982 13574 9034 13626
rect 9046 13574 9098 13626
rect 9110 13574 9162 13626
rect 9174 13574 9226 13626
rect 16982 13574 17034 13626
rect 17046 13574 17098 13626
rect 17110 13574 17162 13626
rect 17174 13574 17226 13626
rect 1860 13472 1912 13524
rect 3240 13515 3292 13524
rect 3240 13481 3249 13515
rect 3249 13481 3283 13515
rect 3283 13481 3292 13515
rect 3240 13472 3292 13481
rect 3424 13472 3476 13524
rect 5908 13472 5960 13524
rect 7472 13515 7524 13524
rect 7472 13481 7481 13515
rect 7481 13481 7515 13515
rect 7515 13481 7524 13515
rect 7472 13472 7524 13481
rect 9312 13515 9364 13524
rect 9312 13481 9321 13515
rect 9321 13481 9355 13515
rect 9355 13481 9364 13515
rect 9312 13472 9364 13481
rect 10140 13472 10192 13524
rect 10784 13472 10836 13524
rect 11520 13515 11572 13524
rect 11520 13481 11529 13515
rect 11529 13481 11563 13515
rect 11563 13481 11572 13515
rect 11520 13472 11572 13481
rect 12808 13472 12860 13524
rect 13452 13472 13504 13524
rect 16764 13472 16816 13524
rect 2688 13404 2740 13456
rect 3700 13404 3752 13456
rect 10876 13404 10928 13456
rect 12072 13404 12124 13456
rect 15936 13404 15988 13456
rect 17408 13404 17460 13456
rect 18052 13404 18104 13456
rect 18788 13404 18840 13456
rect 4620 13379 4672 13388
rect 2320 13268 2372 13320
rect 3332 13268 3384 13320
rect 3884 13268 3936 13320
rect 4620 13345 4629 13379
rect 4629 13345 4663 13379
rect 4663 13345 4672 13379
rect 4620 13336 4672 13345
rect 6092 13379 6144 13388
rect 6092 13345 6101 13379
rect 6101 13345 6135 13379
rect 6135 13345 6144 13379
rect 6092 13336 6144 13345
rect 6460 13268 6512 13320
rect 3884 13175 3936 13184
rect 3884 13141 3893 13175
rect 3893 13141 3927 13175
rect 3927 13141 3936 13175
rect 3884 13132 3936 13141
rect 7932 13336 7984 13388
rect 10508 13379 10560 13388
rect 10508 13345 10517 13379
rect 10517 13345 10551 13379
rect 10551 13345 10560 13379
rect 10508 13336 10560 13345
rect 10784 13336 10836 13388
rect 12164 13336 12216 13388
rect 12624 13268 12676 13320
rect 13820 13311 13872 13320
rect 13820 13277 13829 13311
rect 13829 13277 13863 13311
rect 13863 13277 13872 13311
rect 15476 13311 15528 13320
rect 13820 13268 13872 13277
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 17316 13268 17368 13320
rect 18696 13268 18748 13320
rect 7288 13132 7340 13184
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 10416 13132 10468 13184
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 12982 13030 13034 13082
rect 13046 13030 13098 13082
rect 13110 13030 13162 13082
rect 13174 13030 13226 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 3332 12971 3384 12980
rect 3332 12937 3341 12971
rect 3341 12937 3375 12971
rect 3375 12937 3384 12971
rect 3332 12928 3384 12937
rect 3884 12928 3936 12980
rect 4620 12971 4672 12980
rect 4620 12937 4629 12971
rect 4629 12937 4663 12971
rect 4663 12937 4672 12971
rect 4620 12928 4672 12937
rect 8116 12971 8168 12980
rect 8116 12937 8125 12971
rect 8125 12937 8159 12971
rect 8159 12937 8168 12971
rect 8116 12928 8168 12937
rect 8484 12971 8536 12980
rect 8484 12937 8493 12971
rect 8493 12937 8527 12971
rect 8527 12937 8536 12971
rect 8484 12928 8536 12937
rect 8576 12928 8628 12980
rect 10784 12971 10836 12980
rect 4344 12860 4396 12912
rect 6276 12860 6328 12912
rect 4528 12835 4580 12844
rect 4528 12801 4537 12835
rect 4537 12801 4571 12835
rect 4571 12801 4580 12835
rect 4528 12792 4580 12801
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 12072 12971 12124 12980
rect 12072 12937 12081 12971
rect 12081 12937 12115 12971
rect 12115 12937 12124 12971
rect 12072 12928 12124 12937
rect 12624 12971 12676 12980
rect 12624 12937 12633 12971
rect 12633 12937 12667 12971
rect 12667 12937 12676 12971
rect 12624 12928 12676 12937
rect 12808 12928 12860 12980
rect 3424 12724 3476 12776
rect 2044 12656 2096 12708
rect 2412 12656 2464 12708
rect 4160 12699 4212 12708
rect 4160 12665 4169 12699
rect 4169 12665 4203 12699
rect 4203 12665 4212 12699
rect 4160 12656 4212 12665
rect 2780 12631 2832 12640
rect 2780 12597 2789 12631
rect 2789 12597 2823 12631
rect 2823 12597 2832 12631
rect 2780 12588 2832 12597
rect 6184 12724 6236 12776
rect 5356 12588 5408 12640
rect 5724 12631 5776 12640
rect 5724 12597 5733 12631
rect 5733 12597 5767 12631
rect 5767 12597 5776 12631
rect 5724 12588 5776 12597
rect 6092 12588 6144 12640
rect 6460 12588 6512 12640
rect 7288 12767 7340 12776
rect 7288 12733 7297 12767
rect 7297 12733 7331 12767
rect 7331 12733 7340 12767
rect 7288 12724 7340 12733
rect 9956 12724 10008 12776
rect 10232 12724 10284 12776
rect 10140 12699 10192 12708
rect 8484 12588 8536 12640
rect 10140 12665 10149 12699
rect 10149 12665 10183 12699
rect 10183 12665 10192 12699
rect 10140 12656 10192 12665
rect 10416 12724 10468 12776
rect 16764 12928 16816 12980
rect 17408 12971 17460 12980
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 18696 12903 18748 12912
rect 18696 12869 18705 12903
rect 18705 12869 18739 12903
rect 18739 12869 18748 12903
rect 18696 12860 18748 12869
rect 13452 12792 13504 12844
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 15384 12835 15436 12844
rect 15384 12801 15393 12835
rect 15393 12801 15427 12835
rect 15427 12801 15436 12835
rect 15384 12792 15436 12801
rect 18144 12835 18196 12844
rect 18144 12801 18153 12835
rect 18153 12801 18187 12835
rect 18187 12801 18196 12835
rect 18144 12792 18196 12801
rect 9588 12631 9640 12640
rect 9588 12597 9597 12631
rect 9597 12597 9631 12631
rect 9631 12597 9640 12631
rect 9588 12588 9640 12597
rect 10324 12588 10376 12640
rect 10508 12588 10560 12640
rect 13452 12588 13504 12640
rect 14832 12724 14884 12776
rect 16764 12767 16816 12776
rect 16764 12733 16773 12767
rect 16773 12733 16807 12767
rect 16807 12733 16816 12767
rect 16764 12724 16816 12733
rect 15936 12588 15988 12640
rect 8982 12486 9034 12538
rect 9046 12486 9098 12538
rect 9110 12486 9162 12538
rect 9174 12486 9226 12538
rect 16982 12486 17034 12538
rect 17046 12486 17098 12538
rect 17110 12486 17162 12538
rect 17174 12486 17226 12538
rect 3424 12384 3476 12436
rect 3884 12427 3936 12436
rect 3884 12393 3893 12427
rect 3893 12393 3927 12427
rect 3927 12393 3936 12427
rect 3884 12384 3936 12393
rect 7932 12427 7984 12436
rect 7932 12393 7941 12427
rect 7941 12393 7975 12427
rect 7975 12393 7984 12427
rect 7932 12384 7984 12393
rect 8668 12427 8720 12436
rect 8668 12393 8677 12427
rect 8677 12393 8711 12427
rect 8711 12393 8720 12427
rect 8668 12384 8720 12393
rect 10692 12427 10744 12436
rect 10692 12393 10701 12427
rect 10701 12393 10735 12427
rect 10735 12393 10744 12427
rect 10692 12384 10744 12393
rect 10784 12384 10836 12436
rect 12440 12384 12492 12436
rect 14740 12427 14792 12436
rect 2044 12316 2096 12368
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 4620 12291 4672 12300
rect 2780 12248 2832 12257
rect 4620 12257 4629 12291
rect 4629 12257 4663 12291
rect 4663 12257 4672 12291
rect 4620 12248 4672 12257
rect 6184 12248 6236 12300
rect 9588 12316 9640 12368
rect 13268 12316 13320 12368
rect 14740 12393 14749 12427
rect 14749 12393 14783 12427
rect 14783 12393 14792 12427
rect 14740 12384 14792 12393
rect 15476 12384 15528 12436
rect 18144 12384 18196 12436
rect 21088 12427 21140 12436
rect 21088 12393 21097 12427
rect 21097 12393 21131 12427
rect 21131 12393 21140 12427
rect 21088 12384 21140 12393
rect 13728 12316 13780 12368
rect 6552 12248 6604 12300
rect 1952 12180 2004 12232
rect 5724 12180 5776 12232
rect 6644 12180 6696 12232
rect 9496 12248 9548 12300
rect 10232 12248 10284 12300
rect 15200 12248 15252 12300
rect 19432 12316 19484 12368
rect 16672 12248 16724 12300
rect 17684 12248 17736 12300
rect 20812 12248 20864 12300
rect 8116 12180 8168 12232
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 10416 12223 10468 12232
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 10416 12180 10468 12189
rect 13360 12180 13412 12232
rect 13820 12180 13872 12232
rect 18696 12223 18748 12232
rect 18696 12189 18705 12223
rect 18705 12189 18739 12223
rect 18739 12189 18748 12223
rect 18696 12180 18748 12189
rect 18972 12223 19024 12232
rect 18972 12189 18981 12223
rect 18981 12189 19015 12223
rect 19015 12189 19024 12223
rect 18972 12180 19024 12189
rect 2320 12155 2372 12164
rect 2320 12121 2329 12155
rect 2329 12121 2363 12155
rect 2363 12121 2372 12155
rect 2320 12112 2372 12121
rect 5356 12112 5408 12164
rect 7288 12112 7340 12164
rect 11520 12112 11572 12164
rect 5632 12044 5684 12096
rect 5724 12044 5776 12096
rect 6552 12044 6604 12096
rect 7104 12044 7156 12096
rect 7380 12087 7432 12096
rect 7380 12053 7389 12087
rect 7389 12053 7423 12087
rect 7423 12053 7432 12087
rect 7380 12044 7432 12053
rect 8300 12087 8352 12096
rect 8300 12053 8309 12087
rect 8309 12053 8343 12087
rect 8343 12053 8352 12087
rect 8300 12044 8352 12053
rect 9128 12087 9180 12096
rect 9128 12053 9137 12087
rect 9137 12053 9171 12087
rect 9171 12053 9180 12087
rect 9128 12044 9180 12053
rect 9404 12044 9456 12096
rect 10232 12044 10284 12096
rect 10324 12087 10376 12096
rect 10324 12053 10333 12087
rect 10333 12053 10367 12087
rect 10367 12053 10376 12087
rect 20720 12112 20772 12164
rect 14004 12087 14056 12096
rect 10324 12044 10376 12053
rect 14004 12053 14013 12087
rect 14013 12053 14047 12087
rect 14047 12053 14056 12087
rect 14004 12044 14056 12053
rect 18420 12044 18472 12096
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 12982 11942 13034 11994
rect 13046 11942 13098 11994
rect 13110 11942 13162 11994
rect 13174 11942 13226 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 2044 11883 2096 11892
rect 2044 11849 2053 11883
rect 2053 11849 2087 11883
rect 2087 11849 2096 11883
rect 2044 11840 2096 11849
rect 4620 11883 4672 11892
rect 4620 11849 4629 11883
rect 4629 11849 4663 11883
rect 4663 11849 4672 11883
rect 4620 11840 4672 11849
rect 10048 11840 10100 11892
rect 10600 11883 10652 11892
rect 10600 11849 10609 11883
rect 10609 11849 10643 11883
rect 10643 11849 10652 11883
rect 10600 11840 10652 11849
rect 11152 11883 11204 11892
rect 11152 11849 11161 11883
rect 11161 11849 11195 11883
rect 11195 11849 11204 11883
rect 11152 11840 11204 11849
rect 11520 11883 11572 11892
rect 11520 11849 11529 11883
rect 11529 11849 11563 11883
rect 11563 11849 11572 11883
rect 11520 11840 11572 11849
rect 13360 11883 13412 11892
rect 13360 11849 13369 11883
rect 13369 11849 13403 11883
rect 13403 11849 13412 11883
rect 13360 11840 13412 11849
rect 15200 11840 15252 11892
rect 16672 11883 16724 11892
rect 16672 11849 16681 11883
rect 16681 11849 16715 11883
rect 16715 11849 16724 11883
rect 16672 11840 16724 11849
rect 112 11772 164 11824
rect 2688 11772 2740 11824
rect 4528 11772 4580 11824
rect 6644 11772 6696 11824
rect 3976 11747 4028 11756
rect 3976 11713 3985 11747
rect 3985 11713 4019 11747
rect 4019 11713 4028 11747
rect 3976 11704 4028 11713
rect 2688 11611 2740 11620
rect 2688 11577 2697 11611
rect 2697 11577 2731 11611
rect 2731 11577 2740 11611
rect 2688 11568 2740 11577
rect 3148 11568 3200 11620
rect 5632 11679 5684 11688
rect 2872 11500 2924 11552
rect 3516 11500 3568 11552
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 10232 11772 10284 11824
rect 8392 11704 8444 11756
rect 10140 11704 10192 11756
rect 12072 11772 12124 11824
rect 10784 11704 10836 11756
rect 13268 11772 13320 11824
rect 18420 11772 18472 11824
rect 20812 11772 20864 11824
rect 18972 11747 19024 11756
rect 18972 11713 18981 11747
rect 18981 11713 19015 11747
rect 19015 11713 19024 11747
rect 18972 11704 19024 11713
rect 10416 11636 10468 11688
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12440 11636 12492 11645
rect 5908 11611 5960 11620
rect 5908 11577 5917 11611
rect 5917 11577 5951 11611
rect 5951 11577 5960 11611
rect 5908 11568 5960 11577
rect 6092 11500 6144 11552
rect 7012 11611 7064 11620
rect 7012 11577 7021 11611
rect 7021 11577 7055 11611
rect 7055 11577 7064 11611
rect 7012 11568 7064 11577
rect 7380 11568 7432 11620
rect 9128 11568 9180 11620
rect 9496 11568 9548 11620
rect 8300 11500 8352 11552
rect 9680 11500 9732 11552
rect 10324 11500 10376 11552
rect 13452 11500 13504 11552
rect 14004 11636 14056 11688
rect 15936 11568 15988 11620
rect 18328 11611 18380 11620
rect 18328 11577 18337 11611
rect 18337 11577 18371 11611
rect 18371 11577 18380 11611
rect 18328 11568 18380 11577
rect 18420 11611 18472 11620
rect 18420 11577 18429 11611
rect 18429 11577 18463 11611
rect 18463 11577 18472 11611
rect 18420 11568 18472 11577
rect 18696 11568 18748 11620
rect 17684 11543 17736 11552
rect 17684 11509 17693 11543
rect 17693 11509 17727 11543
rect 17727 11509 17736 11543
rect 17684 11500 17736 11509
rect 19432 11500 19484 11552
rect 8982 11398 9034 11450
rect 9046 11398 9098 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 16982 11398 17034 11450
rect 17046 11398 17098 11450
rect 17110 11398 17162 11450
rect 17174 11398 17226 11450
rect 2688 11296 2740 11348
rect 4712 11296 4764 11348
rect 7012 11296 7064 11348
rect 8392 11296 8444 11348
rect 14004 11296 14056 11348
rect 15936 11339 15988 11348
rect 15936 11305 15945 11339
rect 15945 11305 15979 11339
rect 15979 11305 15988 11339
rect 15936 11296 15988 11305
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 19432 11339 19484 11348
rect 19432 11305 19441 11339
rect 19441 11305 19475 11339
rect 19475 11305 19484 11339
rect 19432 11296 19484 11305
rect 1952 11271 2004 11280
rect 1952 11237 1961 11271
rect 1961 11237 1995 11271
rect 1995 11237 2004 11271
rect 1952 11228 2004 11237
rect 2596 11271 2648 11280
rect 2596 11237 2605 11271
rect 2605 11237 2639 11271
rect 2639 11237 2648 11271
rect 2596 11228 2648 11237
rect 6000 11228 6052 11280
rect 8116 11228 8168 11280
rect 9404 11228 9456 11280
rect 1467 11203 1519 11212
rect 1467 11169 1476 11203
rect 1476 11169 1510 11203
rect 1510 11169 1519 11203
rect 1467 11160 1519 11169
rect 4160 11160 4212 11212
rect 4436 11160 4488 11212
rect 5724 11203 5776 11212
rect 5724 11169 5733 11203
rect 5733 11169 5767 11203
rect 5767 11169 5776 11203
rect 5724 11160 5776 11169
rect 2136 11092 2188 11144
rect 2780 11092 2832 11144
rect 2964 11135 3016 11144
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 5448 11092 5500 11144
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 7380 11092 7432 11144
rect 2320 11024 2372 11076
rect 9496 11160 9548 11212
rect 10048 11228 10100 11280
rect 11060 11228 11112 11280
rect 11520 11228 11572 11280
rect 12072 11228 12124 11280
rect 12256 11228 12308 11280
rect 13544 11228 13596 11280
rect 17408 11228 17460 11280
rect 18328 11271 18380 11280
rect 18328 11237 18337 11271
rect 18337 11237 18371 11271
rect 18371 11237 18380 11271
rect 18328 11228 18380 11237
rect 18420 11160 18472 11212
rect 19156 11160 19208 11212
rect 20720 11160 20772 11212
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 11336 11135 11388 11144
rect 11336 11101 11345 11135
rect 11345 11101 11379 11135
rect 11379 11101 11388 11135
rect 11336 11092 11388 11101
rect 12716 11092 12768 11144
rect 13268 11092 13320 11144
rect 13360 11092 13412 11144
rect 15568 11135 15620 11144
rect 15568 11101 15577 11135
rect 15577 11101 15611 11135
rect 15611 11101 15620 11135
rect 15568 11092 15620 11101
rect 17868 11092 17920 11144
rect 2228 10999 2280 11008
rect 2228 10965 2237 10999
rect 2237 10965 2271 10999
rect 2271 10965 2280 10999
rect 2228 10956 2280 10965
rect 4528 10999 4580 11008
rect 4528 10965 4552 10999
rect 4552 10965 4580 10999
rect 4528 10956 4580 10965
rect 4712 10956 4764 11008
rect 5448 10999 5500 11008
rect 5448 10965 5457 10999
rect 5457 10965 5491 10999
rect 5491 10965 5500 10999
rect 5448 10956 5500 10965
rect 7104 10999 7156 11008
rect 7104 10965 7113 10999
rect 7113 10965 7147 10999
rect 7147 10965 7156 10999
rect 7104 10956 7156 10965
rect 7196 10956 7248 11008
rect 8300 10956 8352 11008
rect 9496 10999 9548 11008
rect 9496 10965 9505 10999
rect 9505 10965 9539 10999
rect 9539 10965 9548 10999
rect 9496 10956 9548 10965
rect 9680 10956 9732 11008
rect 12256 10999 12308 11008
rect 12256 10965 12265 10999
rect 12265 10965 12299 10999
rect 12299 10965 12308 10999
rect 12256 10956 12308 10965
rect 12716 10999 12768 11008
rect 12716 10965 12725 10999
rect 12725 10965 12759 10999
rect 12759 10965 12768 10999
rect 12716 10956 12768 10965
rect 17408 10956 17460 11008
rect 23572 10956 23624 11008
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 12982 10854 13034 10906
rect 13046 10854 13098 10906
rect 13110 10854 13162 10906
rect 13174 10854 13226 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 1492 10752 1544 10804
rect 2412 10752 2464 10804
rect 3424 10752 3476 10804
rect 4344 10795 4396 10804
rect 4344 10761 4353 10795
rect 4353 10761 4387 10795
rect 4387 10761 4396 10795
rect 4344 10752 4396 10761
rect 4712 10752 4764 10804
rect 6000 10795 6052 10804
rect 6000 10761 6009 10795
rect 6009 10761 6043 10795
rect 6043 10761 6052 10795
rect 6000 10752 6052 10761
rect 7104 10752 7156 10804
rect 9404 10795 9456 10804
rect 112 10684 164 10736
rect 2596 10684 2648 10736
rect 2872 10684 2924 10736
rect 4436 10684 4488 10736
rect 5540 10684 5592 10736
rect 8576 10727 8628 10736
rect 8576 10693 8600 10727
rect 8600 10693 8628 10727
rect 8576 10684 8628 10693
rect 9404 10761 9413 10795
rect 9413 10761 9447 10795
rect 9447 10761 9456 10795
rect 9404 10752 9456 10761
rect 10140 10795 10192 10804
rect 10140 10761 10149 10795
rect 10149 10761 10183 10795
rect 10183 10761 10192 10795
rect 10140 10752 10192 10761
rect 11520 10795 11572 10804
rect 11520 10761 11529 10795
rect 11529 10761 11563 10795
rect 11563 10761 11572 10795
rect 11520 10752 11572 10761
rect 13544 10752 13596 10804
rect 15936 10752 15988 10804
rect 17408 10795 17460 10804
rect 17408 10761 17417 10795
rect 17417 10761 17451 10795
rect 17451 10761 17460 10795
rect 17408 10752 17460 10761
rect 19156 10795 19208 10804
rect 19156 10761 19165 10795
rect 19165 10761 19199 10795
rect 19199 10761 19208 10795
rect 19156 10752 19208 10761
rect 20720 10752 20772 10804
rect 10048 10684 10100 10736
rect 5448 10616 5500 10668
rect 6368 10616 6420 10668
rect 17868 10684 17920 10736
rect 11336 10616 11388 10668
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 13360 10659 13412 10668
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 14464 10616 14516 10668
rect 1676 10548 1728 10600
rect 2228 10548 2280 10600
rect 3056 10591 3108 10600
rect 3056 10557 3065 10591
rect 3065 10557 3099 10591
rect 3099 10557 3108 10591
rect 3056 10548 3108 10557
rect 3148 10548 3200 10600
rect 7012 10591 7064 10600
rect 7012 10557 7021 10591
rect 7021 10557 7055 10591
rect 7055 10557 7064 10591
rect 7012 10548 7064 10557
rect 10508 10591 10560 10600
rect 10508 10557 10517 10591
rect 10517 10557 10551 10591
rect 10551 10557 10560 10591
rect 10508 10548 10560 10557
rect 10600 10548 10652 10600
rect 15200 10616 15252 10668
rect 15568 10616 15620 10668
rect 18328 10616 18380 10668
rect 15108 10591 15160 10600
rect 15108 10557 15117 10591
rect 15117 10557 15151 10591
rect 15151 10557 15160 10591
rect 15108 10548 15160 10557
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 4988 10523 5040 10532
rect 4988 10489 4997 10523
rect 4997 10489 5031 10523
rect 5031 10489 5040 10523
rect 4988 10480 5040 10489
rect 5448 10480 5500 10532
rect 5724 10480 5776 10532
rect 8392 10523 8444 10532
rect 8392 10489 8401 10523
rect 8401 10489 8435 10523
rect 8435 10489 8444 10523
rect 8392 10480 8444 10489
rect 12532 10480 12584 10532
rect 18144 10523 18196 10532
rect 18144 10489 18153 10523
rect 18153 10489 18187 10523
rect 18187 10489 18196 10523
rect 18144 10480 18196 10489
rect 3424 10412 3476 10421
rect 4804 10412 4856 10464
rect 5632 10455 5684 10464
rect 5632 10421 5641 10455
rect 5641 10421 5675 10455
rect 5675 10421 5684 10455
rect 5632 10412 5684 10421
rect 6000 10412 6052 10464
rect 6184 10412 6236 10464
rect 8300 10412 8352 10464
rect 8484 10412 8536 10464
rect 9680 10412 9732 10464
rect 17776 10455 17828 10464
rect 17776 10421 17785 10455
rect 17785 10421 17819 10455
rect 17819 10421 17828 10455
rect 17776 10412 17828 10421
rect 8982 10310 9034 10362
rect 9046 10310 9098 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 16982 10310 17034 10362
rect 17046 10310 17098 10362
rect 17110 10310 17162 10362
rect 17174 10310 17226 10362
rect 1676 10251 1728 10260
rect 1676 10217 1685 10251
rect 1685 10217 1719 10251
rect 1719 10217 1728 10251
rect 1676 10208 1728 10217
rect 2136 10208 2188 10260
rect 3056 10208 3108 10260
rect 2596 10183 2648 10192
rect 2596 10149 2605 10183
rect 2605 10149 2639 10183
rect 2639 10149 2648 10183
rect 2596 10140 2648 10149
rect 2964 10140 3016 10192
rect 4160 10140 4212 10192
rect 4988 10208 5040 10260
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 7012 10251 7064 10260
rect 7012 10217 7021 10251
rect 7021 10217 7055 10251
rect 7055 10217 7064 10251
rect 7012 10208 7064 10217
rect 7380 10251 7432 10260
rect 7380 10217 7389 10251
rect 7389 10217 7423 10251
rect 7423 10217 7432 10251
rect 7380 10208 7432 10217
rect 8392 10208 8444 10260
rect 9496 10208 9548 10260
rect 10048 10208 10100 10260
rect 10600 10208 10652 10260
rect 12532 10251 12584 10260
rect 12532 10217 12541 10251
rect 12541 10217 12575 10251
rect 12575 10217 12584 10251
rect 12532 10208 12584 10217
rect 13268 10251 13320 10260
rect 13268 10217 13277 10251
rect 13277 10217 13311 10251
rect 13311 10217 13320 10251
rect 13268 10208 13320 10217
rect 14004 10208 14056 10260
rect 15108 10208 15160 10260
rect 4344 10072 4396 10124
rect 6552 10140 6604 10192
rect 6736 10183 6788 10192
rect 6736 10149 6745 10183
rect 6745 10149 6779 10183
rect 6779 10149 6788 10183
rect 6736 10140 6788 10149
rect 8576 10140 8628 10192
rect 17776 10183 17828 10192
rect 17776 10149 17785 10183
rect 17785 10149 17819 10183
rect 17819 10149 17828 10183
rect 17776 10140 17828 10149
rect 4804 10072 4856 10124
rect 5724 10072 5776 10124
rect 2136 10004 2188 10056
rect 3516 10004 3568 10056
rect 7196 10072 7248 10124
rect 8300 10115 8352 10124
rect 8300 10081 8309 10115
rect 8309 10081 8343 10115
rect 8343 10081 8352 10115
rect 8300 10072 8352 10081
rect 8484 10115 8536 10124
rect 8484 10081 8493 10115
rect 8493 10081 8527 10115
rect 8527 10081 8536 10115
rect 8484 10072 8536 10081
rect 9680 10072 9732 10124
rect 12256 10072 12308 10124
rect 13360 10072 13412 10124
rect 13820 10115 13872 10124
rect 13820 10081 13864 10115
rect 13864 10081 13872 10115
rect 17408 10115 17460 10124
rect 13820 10072 13872 10081
rect 17408 10081 17417 10115
rect 17417 10081 17451 10115
rect 17451 10081 17460 10115
rect 17408 10072 17460 10081
rect 6368 10047 6420 10056
rect 1400 9936 1452 9988
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 6552 10004 6604 10056
rect 8760 10047 8812 10056
rect 8760 10013 8769 10047
rect 8769 10013 8803 10047
rect 8803 10013 8812 10047
rect 8760 10004 8812 10013
rect 6460 9936 6512 9988
rect 4160 9868 4212 9920
rect 5540 9868 5592 9920
rect 6000 9868 6052 9920
rect 6276 9911 6328 9920
rect 6276 9877 6285 9911
rect 6285 9877 6319 9911
rect 6319 9877 6328 9911
rect 9680 9936 9732 9988
rect 6276 9868 6328 9877
rect 10508 9868 10560 9920
rect 11704 9868 11756 9920
rect 14096 9868 14148 9920
rect 18052 9911 18104 9920
rect 18052 9877 18061 9911
rect 18061 9877 18095 9911
rect 18095 9877 18104 9911
rect 18052 9868 18104 9877
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 12982 9766 13034 9818
rect 13046 9766 13098 9818
rect 13110 9766 13162 9818
rect 13174 9766 13226 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 2136 9707 2188 9716
rect 2136 9673 2145 9707
rect 2145 9673 2179 9707
rect 2179 9673 2188 9707
rect 2136 9664 2188 9673
rect 4068 9664 4120 9716
rect 4344 9664 4396 9716
rect 4804 9707 4856 9716
rect 4804 9673 4813 9707
rect 4813 9673 4847 9707
rect 4847 9673 4856 9707
rect 4804 9664 4856 9673
rect 6276 9664 6328 9716
rect 6368 9664 6420 9716
rect 8300 9664 8352 9716
rect 10508 9664 10560 9716
rect 12256 9664 12308 9716
rect 13820 9707 13872 9716
rect 13820 9673 13829 9707
rect 13829 9673 13863 9707
rect 13863 9673 13872 9707
rect 13820 9664 13872 9673
rect 18052 9664 18104 9716
rect 112 9596 164 9648
rect 2596 9528 2648 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 4988 9460 5040 9512
rect 5448 9460 5500 9512
rect 9956 9596 10008 9648
rect 11520 9596 11572 9648
rect 17408 9596 17460 9648
rect 10232 9528 10284 9580
rect 12716 9528 12768 9580
rect 7196 9503 7248 9512
rect 7196 9469 7205 9503
rect 7205 9469 7239 9503
rect 7239 9469 7248 9503
rect 7196 9460 7248 9469
rect 4160 9392 4212 9444
rect 4528 9392 4580 9444
rect 6460 9392 6512 9444
rect 9956 9460 10008 9512
rect 7840 9392 7892 9444
rect 8484 9392 8536 9444
rect 5356 9367 5408 9376
rect 5356 9333 5365 9367
rect 5365 9333 5399 9367
rect 5399 9333 5408 9367
rect 5356 9324 5408 9333
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 9772 9324 9824 9376
rect 10232 9435 10284 9444
rect 10232 9401 10241 9435
rect 10241 9401 10275 9435
rect 10275 9401 10284 9435
rect 10232 9392 10284 9401
rect 11152 9392 11204 9444
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 17408 9324 17460 9333
rect 8982 9222 9034 9274
rect 9046 9222 9098 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 16982 9222 17034 9274
rect 17046 9222 17098 9274
rect 17110 9222 17162 9274
rect 17174 9222 17226 9274
rect 2872 9120 2924 9172
rect 2964 9120 3016 9172
rect 3608 9120 3660 9172
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 6460 9163 6512 9172
rect 6460 9129 6469 9163
rect 6469 9129 6503 9163
rect 6503 9129 6512 9163
rect 6460 9120 6512 9129
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 9956 9120 10008 9172
rect 10232 9120 10284 9172
rect 3792 9052 3844 9104
rect 1952 9027 2004 9036
rect 1952 8993 1961 9027
rect 1961 8993 1995 9027
rect 1995 8993 2004 9027
rect 1952 8984 2004 8993
rect 2228 8984 2280 9036
rect 5356 9052 5408 9104
rect 5908 9052 5960 9104
rect 9772 9052 9824 9104
rect 6092 8984 6144 9036
rect 7840 9027 7892 9036
rect 5632 8916 5684 8968
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 8760 8984 8812 9036
rect 13728 9027 13780 9036
rect 13728 8993 13737 9027
rect 13737 8993 13771 9027
rect 13771 8993 13780 9027
rect 13728 8984 13780 8993
rect 14464 8984 14516 9036
rect 8116 8916 8168 8968
rect 13544 8916 13596 8968
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 5724 8780 5776 8832
rect 10876 8823 10928 8832
rect 10876 8789 10885 8823
rect 10885 8789 10919 8823
rect 10919 8789 10928 8823
rect 10876 8780 10928 8789
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 12982 8678 13034 8730
rect 13046 8678 13098 8730
rect 13110 8678 13162 8730
rect 13174 8678 13226 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 5356 8576 5408 8628
rect 7840 8576 7892 8628
rect 8760 8576 8812 8628
rect 9956 8619 10008 8628
rect 9956 8585 9965 8619
rect 9965 8585 9999 8619
rect 9999 8585 10008 8619
rect 9956 8576 10008 8585
rect 2228 8483 2280 8492
rect 2228 8449 2237 8483
rect 2237 8449 2271 8483
rect 2271 8449 2280 8483
rect 2228 8440 2280 8449
rect 4068 8440 4120 8492
rect 4712 8440 4764 8492
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 10876 8440 10928 8492
rect 3976 8415 4028 8424
rect 3976 8381 3985 8415
rect 3985 8381 4019 8415
rect 4019 8381 4028 8415
rect 3976 8372 4028 8381
rect 7748 8372 7800 8424
rect 1768 8304 1820 8356
rect 2596 8279 2648 8288
rect 2596 8245 2605 8279
rect 2605 8245 2639 8279
rect 2639 8245 2648 8279
rect 2596 8236 2648 8245
rect 2872 8279 2924 8288
rect 2872 8245 2881 8279
rect 2881 8245 2915 8279
rect 2915 8245 2924 8279
rect 2872 8236 2924 8245
rect 3792 8279 3844 8288
rect 3792 8245 3801 8279
rect 3801 8245 3835 8279
rect 3835 8245 3844 8279
rect 3792 8236 3844 8245
rect 5448 8304 5500 8356
rect 11152 8347 11204 8356
rect 7288 8279 7340 8288
rect 7288 8245 7297 8279
rect 7297 8245 7331 8279
rect 7331 8245 7340 8279
rect 7288 8236 7340 8245
rect 8116 8279 8168 8288
rect 8116 8245 8125 8279
rect 8125 8245 8159 8279
rect 8159 8245 8168 8279
rect 8116 8236 8168 8245
rect 10324 8279 10376 8288
rect 10324 8245 10333 8279
rect 10333 8245 10367 8279
rect 10367 8245 10376 8279
rect 11152 8313 11161 8347
rect 11161 8313 11195 8347
rect 11195 8313 11204 8347
rect 11152 8304 11204 8313
rect 13728 8279 13780 8288
rect 10324 8236 10376 8245
rect 13728 8245 13737 8279
rect 13737 8245 13771 8279
rect 13771 8245 13780 8279
rect 13728 8236 13780 8245
rect 8982 8134 9034 8186
rect 9046 8134 9098 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 16982 8134 17034 8186
rect 17046 8134 17098 8186
rect 17110 8134 17162 8186
rect 17174 8134 17226 8186
rect 1768 8032 1820 8084
rect 2872 8032 2924 8084
rect 3976 8032 4028 8084
rect 1952 8007 2004 8016
rect 1952 7973 1961 8007
rect 1961 7973 1995 8007
rect 1995 7973 2004 8007
rect 1952 7964 2004 7973
rect 2228 7964 2280 8016
rect 5632 8075 5684 8084
rect 5632 8041 5641 8075
rect 5641 8041 5675 8075
rect 5675 8041 5684 8075
rect 5632 8032 5684 8041
rect 10324 8075 10376 8084
rect 10324 8041 10333 8075
rect 10333 8041 10367 8075
rect 10367 8041 10376 8075
rect 10324 8032 10376 8041
rect 4344 8007 4396 8016
rect 4344 7973 4353 8007
rect 4353 7973 4387 8007
rect 4387 7973 4396 8007
rect 4344 7964 4396 7973
rect 7288 8007 7340 8016
rect 7288 7973 7297 8007
rect 7297 7973 7331 8007
rect 7331 7973 7340 8007
rect 7288 7964 7340 7973
rect 11152 7964 11204 8016
rect 3792 7896 3844 7948
rect 10232 7939 10284 7948
rect 10232 7905 10241 7939
rect 10241 7905 10275 7939
rect 10275 7905 10284 7939
rect 10232 7896 10284 7905
rect 12072 7939 12124 7948
rect 2136 7828 2188 7880
rect 6276 7828 6328 7880
rect 8208 7828 8260 7880
rect 11704 7828 11756 7880
rect 12072 7905 12081 7939
rect 12081 7905 12115 7939
rect 12115 7905 12124 7939
rect 12072 7896 12124 7905
rect 19248 7939 19300 7948
rect 19248 7905 19292 7939
rect 19292 7905 19300 7939
rect 19248 7896 19300 7905
rect 12348 7871 12400 7880
rect 1308 7760 1360 7812
rect 5724 7760 5776 7812
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 13544 7760 13596 7812
rect 3976 7692 4028 7744
rect 4528 7692 4580 7744
rect 4712 7692 4764 7744
rect 6828 7735 6880 7744
rect 6828 7701 6837 7735
rect 6837 7701 6871 7735
rect 6871 7701 6880 7735
rect 6828 7692 6880 7701
rect 8760 7692 8812 7744
rect 12716 7692 12768 7744
rect 19984 7692 20036 7744
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 12982 7590 13034 7642
rect 13046 7590 13098 7642
rect 13110 7590 13162 7642
rect 13174 7590 13226 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 112 7488 164 7540
rect 2136 7463 2188 7472
rect 2136 7429 2145 7463
rect 2145 7429 2179 7463
rect 2179 7429 2188 7463
rect 2136 7420 2188 7429
rect 3884 7420 3936 7472
rect 5724 7488 5776 7540
rect 6276 7531 6328 7540
rect 6276 7497 6285 7531
rect 6285 7497 6319 7531
rect 6319 7497 6328 7531
rect 6276 7488 6328 7497
rect 7748 7531 7800 7540
rect 7748 7497 7757 7531
rect 7757 7497 7791 7531
rect 7791 7497 7800 7531
rect 7748 7488 7800 7497
rect 8024 7488 8076 7540
rect 10232 7488 10284 7540
rect 11704 7531 11756 7540
rect 11704 7497 11713 7531
rect 11713 7497 11747 7531
rect 11747 7497 11756 7531
rect 11704 7488 11756 7497
rect 12072 7531 12124 7540
rect 12072 7497 12081 7531
rect 12081 7497 12115 7531
rect 12115 7497 12124 7531
rect 12072 7488 12124 7497
rect 14556 7488 14608 7540
rect 19248 7531 19300 7540
rect 19248 7497 19257 7531
rect 19257 7497 19291 7531
rect 19291 7497 19300 7531
rect 19248 7488 19300 7497
rect 21456 7531 21508 7540
rect 21456 7497 21465 7531
rect 21465 7497 21499 7531
rect 21499 7497 21508 7531
rect 21456 7488 21508 7497
rect 4804 7420 4856 7472
rect 6184 7420 6236 7472
rect 3976 7352 4028 7404
rect 4620 7352 4672 7404
rect 8760 7352 8812 7404
rect 13452 7395 13504 7404
rect 13452 7361 13461 7395
rect 13461 7361 13495 7395
rect 13495 7361 13504 7395
rect 13452 7352 13504 7361
rect 6000 7284 6052 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 9864 7284 9916 7336
rect 21456 7284 21508 7336
rect 1584 7259 1636 7268
rect 1584 7225 1593 7259
rect 1593 7225 1627 7259
rect 1627 7225 1636 7259
rect 1584 7216 1636 7225
rect 4160 7259 4212 7268
rect 4160 7225 4169 7259
rect 4169 7225 4203 7259
rect 4203 7225 4212 7259
rect 4160 7216 4212 7225
rect 4436 7216 4488 7268
rect 4620 7216 4672 7268
rect 2504 7191 2556 7200
rect 2504 7157 2513 7191
rect 2513 7157 2547 7191
rect 2547 7157 2556 7191
rect 2504 7148 2556 7157
rect 2872 7148 2924 7200
rect 3976 7148 4028 7200
rect 4528 7148 4580 7200
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 9312 7259 9364 7268
rect 5632 7191 5684 7200
rect 5172 7148 5224 7157
rect 5632 7157 5641 7191
rect 5641 7157 5675 7191
rect 5675 7157 5684 7191
rect 5632 7148 5684 7157
rect 9312 7225 9321 7259
rect 9321 7225 9355 7259
rect 9355 7225 9364 7259
rect 9312 7216 9364 7225
rect 11704 7216 11756 7268
rect 12716 7216 12768 7268
rect 12808 7191 12860 7200
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 12808 7148 12860 7157
rect 17316 7148 17368 7200
rect 8982 7046 9034 7098
rect 9046 7046 9098 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 17174 7046 17226 7098
rect 1584 6944 1636 6996
rect 2872 6987 2924 6996
rect 2872 6953 2881 6987
rect 2881 6953 2915 6987
rect 2915 6953 2924 6987
rect 2872 6944 2924 6953
rect 3792 6944 3844 6996
rect 2044 6876 2096 6928
rect 6092 6944 6144 6996
rect 6828 6987 6880 6996
rect 6828 6953 6837 6987
rect 6837 6953 6871 6987
rect 6871 6953 6880 6987
rect 6828 6944 6880 6953
rect 7288 6987 7340 6996
rect 7288 6953 7297 6987
rect 7297 6953 7331 6987
rect 7331 6953 7340 6987
rect 7288 6944 7340 6953
rect 2412 6808 2464 6860
rect 3792 6808 3844 6860
rect 6000 6876 6052 6928
rect 9312 6944 9364 6996
rect 11704 6987 11756 6996
rect 11704 6953 11713 6987
rect 11713 6953 11747 6987
rect 11747 6953 11756 6987
rect 11704 6944 11756 6953
rect 12348 6944 12400 6996
rect 4528 6851 4580 6860
rect 4528 6817 4537 6851
rect 4537 6817 4571 6851
rect 4571 6817 4580 6851
rect 4528 6808 4580 6817
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 6920 6851 6972 6860
rect 4160 6740 4212 6792
rect 6368 6740 6420 6792
rect 6920 6817 6929 6851
rect 6929 6817 6963 6851
rect 6963 6817 6972 6851
rect 6920 6808 6972 6817
rect 2044 6672 2096 6724
rect 4344 6672 4396 6724
rect 5172 6672 5224 6724
rect 8024 6919 8076 6928
rect 8024 6885 8033 6919
rect 8033 6885 8067 6919
rect 8067 6885 8076 6919
rect 9864 6919 9916 6928
rect 8024 6876 8076 6885
rect 9864 6885 9873 6919
rect 9873 6885 9907 6919
rect 9907 6885 9916 6919
rect 9864 6876 9916 6885
rect 12256 6876 12308 6928
rect 13452 6919 13504 6928
rect 13452 6885 13461 6919
rect 13461 6885 13495 6919
rect 13495 6885 13504 6919
rect 13452 6876 13504 6885
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 11244 6740 11296 6792
rect 9312 6672 9364 6724
rect 12716 6672 12768 6724
rect 1952 6604 2004 6656
rect 2504 6604 2556 6656
rect 3884 6647 3936 6656
rect 3884 6613 3893 6647
rect 3893 6613 3927 6647
rect 3927 6613 3936 6647
rect 3884 6604 3936 6613
rect 7012 6604 7064 6656
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 12982 6502 13034 6554
rect 13046 6502 13098 6554
rect 13110 6502 13162 6554
rect 13174 6502 13226 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 20 6400 72 6452
rect 3792 6443 3844 6452
rect 2136 6375 2188 6384
rect 2136 6341 2145 6375
rect 2145 6341 2179 6375
rect 2179 6341 2188 6375
rect 2136 6332 2188 6341
rect 3792 6409 3801 6443
rect 3801 6409 3835 6443
rect 3835 6409 3844 6443
rect 3792 6400 3844 6409
rect 5540 6400 5592 6452
rect 6184 6400 6236 6452
rect 6368 6443 6420 6452
rect 6368 6409 6377 6443
rect 6377 6409 6411 6443
rect 6411 6409 6420 6443
rect 6368 6400 6420 6409
rect 9864 6400 9916 6452
rect 3884 6332 3936 6384
rect 6460 6332 6512 6384
rect 3792 6264 3844 6316
rect 11060 6264 11112 6316
rect 11244 6307 11296 6316
rect 11244 6273 11253 6307
rect 11253 6273 11287 6307
rect 11287 6273 11296 6307
rect 11244 6264 11296 6273
rect 12348 6264 12400 6316
rect 12716 6264 12768 6316
rect 1400 6128 1452 6180
rect 1676 6171 1728 6180
rect 1676 6137 1685 6171
rect 1685 6137 1719 6171
rect 1719 6137 1728 6171
rect 5724 6196 5776 6248
rect 6184 6196 6236 6248
rect 7748 6239 7800 6248
rect 7748 6205 7757 6239
rect 7757 6205 7791 6239
rect 7791 6205 7800 6239
rect 7748 6196 7800 6205
rect 1676 6128 1728 6137
rect 5448 6128 5500 6180
rect 2044 6060 2096 6112
rect 2504 6103 2556 6112
rect 2504 6069 2513 6103
rect 2513 6069 2547 6103
rect 2547 6069 2556 6103
rect 2504 6060 2556 6069
rect 2872 6103 2924 6112
rect 2872 6069 2881 6103
rect 2881 6069 2915 6103
rect 2915 6069 2924 6103
rect 2872 6060 2924 6069
rect 3884 6060 3936 6112
rect 7012 6103 7064 6112
rect 7012 6069 7021 6103
rect 7021 6069 7055 6103
rect 7055 6069 7064 6103
rect 7012 6060 7064 6069
rect 7472 6103 7524 6112
rect 7472 6069 7481 6103
rect 7481 6069 7515 6103
rect 7515 6069 7524 6103
rect 7472 6060 7524 6069
rect 8116 6060 8168 6112
rect 9956 6171 10008 6180
rect 9956 6137 9959 6171
rect 9959 6137 9993 6171
rect 9993 6137 10008 6171
rect 9956 6128 10008 6137
rect 12256 6128 12308 6180
rect 13728 6196 13780 6248
rect 13820 6196 13872 6248
rect 14464 6196 14516 6248
rect 15108 6171 15160 6180
rect 15108 6137 15117 6171
rect 15117 6137 15151 6171
rect 15151 6137 15160 6171
rect 15108 6128 15160 6137
rect 11796 6060 11848 6112
rect 8982 5958 9034 6010
rect 9046 5958 9098 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 17174 5958 17226 6010
rect 2412 5899 2464 5908
rect 2412 5865 2421 5899
rect 2421 5865 2455 5899
rect 2455 5865 2464 5899
rect 2412 5856 2464 5865
rect 2596 5856 2648 5908
rect 4528 5856 4580 5908
rect 8024 5899 8076 5908
rect 8024 5865 8033 5899
rect 8033 5865 8067 5899
rect 8067 5865 8076 5899
rect 8024 5856 8076 5865
rect 9312 5856 9364 5908
rect 12808 5899 12860 5908
rect 12808 5865 12817 5899
rect 12817 5865 12851 5899
rect 12851 5865 12860 5899
rect 12808 5856 12860 5865
rect 14464 5899 14516 5908
rect 14464 5865 14473 5899
rect 14473 5865 14507 5899
rect 14507 5865 14516 5899
rect 14464 5856 14516 5865
rect 15108 5856 15160 5908
rect 15568 5899 15620 5908
rect 15568 5865 15577 5899
rect 15577 5865 15611 5899
rect 15611 5865 15620 5899
rect 15568 5856 15620 5865
rect 1676 5788 1728 5840
rect 2872 5788 2924 5840
rect 7012 5788 7064 5840
rect 9404 5788 9456 5840
rect 1952 5763 2004 5772
rect 1952 5729 1961 5763
rect 1961 5729 1995 5763
rect 1995 5729 2004 5763
rect 1952 5720 2004 5729
rect 4160 5720 4212 5772
rect 5448 5720 5500 5772
rect 6000 5763 6052 5772
rect 6000 5729 6009 5763
rect 6009 5729 6043 5763
rect 6043 5729 6052 5763
rect 6000 5720 6052 5729
rect 8208 5763 8260 5772
rect 8208 5729 8217 5763
rect 8217 5729 8251 5763
rect 8251 5729 8260 5763
rect 8208 5720 8260 5729
rect 4528 5652 4580 5704
rect 1400 5584 1452 5636
rect 7748 5695 7800 5704
rect 4896 5584 4948 5636
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 9496 5652 9548 5704
rect 9404 5584 9456 5636
rect 3792 5516 3844 5568
rect 4344 5516 4396 5568
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 5632 5516 5684 5568
rect 6184 5559 6236 5568
rect 6184 5525 6193 5559
rect 6193 5525 6227 5559
rect 6227 5525 6236 5559
rect 6184 5516 6236 5525
rect 7840 5516 7892 5568
rect 11428 5720 11480 5772
rect 12256 5720 12308 5772
rect 9956 5652 10008 5704
rect 10508 5652 10560 5704
rect 14464 5652 14516 5704
rect 10048 5584 10100 5636
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 12982 5414 13034 5466
rect 13046 5414 13098 5466
rect 13110 5414 13162 5466
rect 13174 5414 13226 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 3792 5312 3844 5364
rect 4528 5355 4580 5364
rect 4528 5321 4537 5355
rect 4537 5321 4571 5355
rect 4571 5321 4580 5355
rect 4528 5312 4580 5321
rect 5448 5312 5500 5364
rect 6460 5355 6512 5364
rect 6460 5321 6469 5355
rect 6469 5321 6503 5355
rect 6503 5321 6512 5355
rect 6460 5312 6512 5321
rect 9956 5355 10008 5364
rect 9956 5321 9965 5355
rect 9965 5321 9999 5355
rect 9999 5321 10008 5355
rect 9956 5312 10008 5321
rect 10048 5312 10100 5364
rect 5540 5244 5592 5296
rect 9864 5244 9916 5296
rect 3608 5176 3660 5228
rect 4160 5219 4212 5228
rect 4160 5185 4169 5219
rect 4169 5185 4203 5219
rect 4203 5185 4212 5219
rect 5356 5219 5408 5228
rect 4160 5176 4212 5185
rect 1860 5040 1912 5092
rect 3792 4972 3844 5024
rect 3976 4972 4028 5024
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 4988 5151 5040 5160
rect 4988 5117 4997 5151
rect 4997 5117 5031 5151
rect 5031 5117 5040 5151
rect 4988 5108 5040 5117
rect 6460 5108 6512 5160
rect 6736 5108 6788 5160
rect 8576 5151 8628 5160
rect 8576 5117 8585 5151
rect 8585 5117 8619 5151
rect 8619 5117 8628 5151
rect 8576 5108 8628 5117
rect 9772 5151 9824 5160
rect 9772 5117 9781 5151
rect 9781 5117 9815 5151
rect 9815 5117 9824 5151
rect 10416 5312 10468 5364
rect 12072 5312 12124 5364
rect 12256 5355 12308 5364
rect 12256 5321 12265 5355
rect 12265 5321 12299 5355
rect 12299 5321 12308 5355
rect 12256 5312 12308 5321
rect 10784 5244 10836 5296
rect 11428 5287 11480 5296
rect 11428 5253 11437 5287
rect 11437 5253 11471 5287
rect 11471 5253 11480 5287
rect 11428 5244 11480 5253
rect 10508 5176 10560 5228
rect 15568 5219 15620 5228
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 15568 5176 15620 5185
rect 9772 5108 9824 5117
rect 12164 5108 12216 5160
rect 13544 5151 13596 5160
rect 13544 5117 13553 5151
rect 13553 5117 13587 5151
rect 13587 5117 13596 5151
rect 13544 5108 13596 5117
rect 14188 5151 14240 5160
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 14464 5108 14516 5160
rect 8668 5040 8720 5092
rect 9312 5040 9364 5092
rect 9496 5040 9548 5092
rect 11980 5040 12032 5092
rect 14372 5083 14424 5092
rect 14372 5049 14381 5083
rect 14381 5049 14415 5083
rect 14415 5049 14424 5083
rect 14372 5040 14424 5049
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 5632 4972 5684 4981
rect 8208 4972 8260 5024
rect 8852 4972 8904 5024
rect 15384 5015 15436 5024
rect 15384 4981 15393 5015
rect 15393 4981 15427 5015
rect 15427 4981 15436 5015
rect 16488 5015 16540 5024
rect 15384 4972 15436 4981
rect 16488 4981 16497 5015
rect 16497 4981 16531 5015
rect 16531 4981 16540 5015
rect 16488 4972 16540 4981
rect 8982 4870 9034 4922
rect 9046 4870 9098 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 17174 4870 17226 4922
rect 1952 4811 2004 4820
rect 1952 4777 1961 4811
rect 1961 4777 1995 4811
rect 1995 4777 2004 4811
rect 1952 4768 2004 4777
rect 4344 4811 4396 4820
rect 4344 4777 4353 4811
rect 4353 4777 4387 4811
rect 4387 4777 4396 4811
rect 4344 4768 4396 4777
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 6000 4811 6052 4820
rect 6000 4777 6009 4811
rect 6009 4777 6043 4811
rect 6043 4777 6052 4811
rect 6000 4768 6052 4777
rect 7012 4768 7064 4820
rect 1584 4632 1636 4684
rect 2688 4675 2740 4684
rect 2688 4641 2697 4675
rect 2697 4641 2731 4675
rect 2731 4641 2740 4675
rect 2688 4632 2740 4641
rect 4620 4700 4672 4752
rect 4068 4632 4120 4684
rect 4528 4675 4580 4684
rect 4528 4641 4537 4675
rect 4537 4641 4571 4675
rect 4571 4641 4580 4675
rect 4528 4632 4580 4641
rect 6184 4700 6236 4752
rect 8760 4768 8812 4820
rect 14188 4768 14240 4820
rect 14372 4768 14424 4820
rect 7748 4700 7800 4752
rect 5632 4632 5684 4684
rect 3148 4607 3200 4616
rect 3148 4573 3157 4607
rect 3157 4573 3191 4607
rect 3191 4573 3200 4607
rect 3148 4564 3200 4573
rect 3976 4564 4028 4616
rect 4988 4564 5040 4616
rect 5356 4564 5408 4616
rect 6460 4564 6512 4616
rect 4712 4496 4764 4548
rect 7656 4496 7708 4548
rect 6828 4428 6880 4480
rect 7840 4632 7892 4684
rect 9772 4700 9824 4752
rect 10784 4743 10836 4752
rect 10784 4709 10793 4743
rect 10793 4709 10827 4743
rect 10827 4709 10836 4743
rect 10784 4700 10836 4709
rect 11796 4700 11848 4752
rect 16488 4700 16540 4752
rect 17224 4700 17276 4752
rect 8392 4632 8444 4684
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 10416 4632 10468 4684
rect 11060 4632 11112 4684
rect 12532 4675 12584 4684
rect 12532 4641 12541 4675
rect 12541 4641 12575 4675
rect 12575 4641 12584 4675
rect 12532 4632 12584 4641
rect 13452 4632 13504 4684
rect 16120 4632 16172 4684
rect 11152 4564 11204 4616
rect 17500 4564 17552 4616
rect 18420 4564 18472 4616
rect 8760 4471 8812 4480
rect 8760 4437 8769 4471
rect 8769 4437 8803 4471
rect 8803 4437 8812 4471
rect 12256 4471 12308 4480
rect 8760 4428 8812 4437
rect 12256 4437 12265 4471
rect 12265 4437 12299 4471
rect 12299 4437 12308 4471
rect 12256 4428 12308 4437
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 18052 4428 18104 4480
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 12982 4326 13034 4378
rect 13046 4326 13098 4378
rect 13110 4326 13162 4378
rect 13174 4326 13226 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 1584 4267 1636 4276
rect 1584 4233 1593 4267
rect 1593 4233 1627 4267
rect 1627 4233 1636 4267
rect 1584 4224 1636 4233
rect 2688 4224 2740 4276
rect 3700 4224 3752 4276
rect 4528 4224 4580 4276
rect 3148 4088 3200 4140
rect 3700 4131 3752 4140
rect 3700 4097 3709 4131
rect 3709 4097 3743 4131
rect 3743 4097 3752 4131
rect 3700 4088 3752 4097
rect 6184 4224 6236 4276
rect 10048 4224 10100 4276
rect 10416 4224 10468 4276
rect 11152 4267 11204 4276
rect 11152 4233 11161 4267
rect 11161 4233 11195 4267
rect 11195 4233 11204 4267
rect 11152 4224 11204 4233
rect 11796 4267 11848 4276
rect 11796 4233 11805 4267
rect 11805 4233 11839 4267
rect 11839 4233 11848 4267
rect 11796 4224 11848 4233
rect 13820 4224 13872 4276
rect 14648 4224 14700 4276
rect 17224 4267 17276 4276
rect 17224 4233 17233 4267
rect 17233 4233 17267 4267
rect 17267 4233 17276 4267
rect 17224 4224 17276 4233
rect 8116 4156 8168 4208
rect 2320 3995 2372 4004
rect 2320 3961 2329 3995
rect 2329 3961 2363 3995
rect 2363 3961 2372 3995
rect 2320 3952 2372 3961
rect 2136 3927 2188 3936
rect 2136 3893 2145 3927
rect 2145 3893 2179 3927
rect 2179 3893 2188 3927
rect 3884 4020 3936 4072
rect 4804 4020 4856 4072
rect 2136 3884 2188 3893
rect 2596 3884 2648 3936
rect 4528 3952 4580 4004
rect 7748 4131 7800 4140
rect 6828 4020 6880 4072
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 8760 4088 8812 4140
rect 10048 4088 10100 4140
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 12808 4131 12860 4140
rect 12808 4097 12817 4131
rect 12817 4097 12851 4131
rect 12851 4097 12860 4131
rect 12808 4088 12860 4097
rect 7472 4020 7524 4072
rect 11152 4020 11204 4072
rect 8392 3995 8444 4004
rect 8392 3961 8401 3995
rect 8401 3961 8435 3995
rect 8435 3961 8444 3995
rect 8392 3952 8444 3961
rect 4160 3884 4212 3936
rect 4804 3884 4856 3936
rect 7288 3927 7340 3936
rect 7288 3893 7297 3927
rect 7297 3893 7331 3927
rect 7331 3893 7340 3927
rect 7288 3884 7340 3893
rect 8116 3884 8168 3936
rect 12900 3952 12952 4004
rect 16120 4156 16172 4208
rect 14372 4088 14424 4140
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 18420 4131 18472 4140
rect 18420 4097 18429 4131
rect 18429 4097 18463 4131
rect 18463 4097 18472 4131
rect 18420 4088 18472 4097
rect 15384 3952 15436 4004
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 12532 3884 12584 3936
rect 13452 3927 13504 3936
rect 13452 3893 13461 3927
rect 13461 3893 13495 3927
rect 13495 3893 13504 3927
rect 13452 3884 13504 3893
rect 16120 3995 16172 4004
rect 16120 3961 16129 3995
rect 16129 3961 16163 3995
rect 16163 3961 16172 3995
rect 16120 3952 16172 3961
rect 16396 3884 16448 3936
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 18052 3884 18104 3936
rect 18236 3995 18288 4004
rect 18236 3961 18245 3995
rect 18245 3961 18279 3995
rect 18279 3961 18288 3995
rect 18236 3952 18288 3961
rect 8982 3782 9034 3834
rect 9046 3782 9098 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 17174 3782 17226 3834
rect 3700 3723 3752 3732
rect 3700 3689 3709 3723
rect 3709 3689 3743 3723
rect 3743 3689 3752 3723
rect 3700 3680 3752 3689
rect 4620 3723 4672 3732
rect 4620 3689 4629 3723
rect 4629 3689 4663 3723
rect 4663 3689 4672 3723
rect 4620 3680 4672 3689
rect 6000 3680 6052 3732
rect 7748 3680 7800 3732
rect 8484 3723 8536 3732
rect 8484 3689 8493 3723
rect 8493 3689 8527 3723
rect 8527 3689 8536 3723
rect 8484 3680 8536 3689
rect 8760 3680 8812 3732
rect 12256 3680 12308 3732
rect 4528 3612 4580 3664
rect 5448 3612 5500 3664
rect 8116 3612 8168 3664
rect 9496 3612 9548 3664
rect 10048 3612 10100 3664
rect 10692 3612 10744 3664
rect 12072 3655 12124 3664
rect 12072 3621 12081 3655
rect 12081 3621 12115 3655
rect 12115 3621 12124 3655
rect 12072 3612 12124 3621
rect 12808 3612 12860 3664
rect 12900 3612 12952 3664
rect 17500 3680 17552 3732
rect 15568 3612 15620 3664
rect 15752 3612 15804 3664
rect 16028 3655 16080 3664
rect 16028 3621 16037 3655
rect 16037 3621 16071 3655
rect 16071 3621 16080 3655
rect 16028 3612 16080 3621
rect 16304 3612 16356 3664
rect 17776 3612 17828 3664
rect 18236 3612 18288 3664
rect 2228 3587 2280 3596
rect 2228 3553 2237 3587
rect 2237 3553 2271 3587
rect 2271 3553 2280 3587
rect 2228 3544 2280 3553
rect 2320 3544 2372 3596
rect 4620 3544 4672 3596
rect 5356 3544 5408 3596
rect 7288 3544 7340 3596
rect 8668 3544 8720 3596
rect 13544 3587 13596 3596
rect 13544 3553 13553 3587
rect 13553 3553 13587 3587
rect 13587 3553 13596 3587
rect 13544 3544 13596 3553
rect 17316 3587 17368 3596
rect 17316 3553 17325 3587
rect 17325 3553 17359 3587
rect 17359 3553 17368 3587
rect 17316 3544 17368 3553
rect 3976 3476 4028 3528
rect 6828 3476 6880 3528
rect 10048 3519 10100 3528
rect 10048 3485 10057 3519
rect 10057 3485 10091 3519
rect 10091 3485 10100 3519
rect 10048 3476 10100 3485
rect 11980 3519 12032 3528
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 16120 3476 16172 3528
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 18420 3476 18472 3528
rect 2504 3340 2556 3392
rect 4344 3340 4396 3392
rect 6460 3383 6512 3392
rect 6460 3349 6469 3383
rect 6469 3349 6503 3383
rect 6503 3349 6512 3383
rect 6460 3340 6512 3349
rect 11152 3340 11204 3392
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 12982 3238 13034 3290
rect 13046 3238 13098 3290
rect 13110 3238 13162 3290
rect 13174 3238 13226 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 1400 3136 1452 3188
rect 1216 2932 1268 2984
rect 2504 2975 2556 2984
rect 2504 2941 2513 2975
rect 2513 2941 2547 2975
rect 2547 2941 2556 2975
rect 4160 3136 4212 3188
rect 5448 3136 5500 3188
rect 5816 3136 5868 3188
rect 7288 3136 7340 3188
rect 8116 3179 8168 3188
rect 8116 3145 8125 3179
rect 8125 3145 8159 3179
rect 8159 3145 8168 3179
rect 8116 3136 8168 3145
rect 9312 3136 9364 3188
rect 12072 3136 12124 3188
rect 13544 3179 13596 3188
rect 13544 3145 13553 3179
rect 13553 3145 13587 3179
rect 13587 3145 13596 3179
rect 13544 3136 13596 3145
rect 15752 3179 15804 3188
rect 15752 3145 15761 3179
rect 15761 3145 15795 3179
rect 15795 3145 15804 3179
rect 15752 3136 15804 3145
rect 16120 3179 16172 3188
rect 16120 3145 16129 3179
rect 16129 3145 16163 3179
rect 16163 3145 16172 3179
rect 16120 3136 16172 3145
rect 4252 3068 4304 3120
rect 9404 3068 9456 3120
rect 2504 2932 2556 2941
rect 3148 2907 3200 2916
rect 3148 2873 3157 2907
rect 3157 2873 3191 2907
rect 3191 2873 3200 2907
rect 3148 2864 3200 2873
rect 3516 2864 3568 2916
rect 4804 3000 4856 3052
rect 8668 3000 8720 3052
rect 10048 3000 10100 3052
rect 4160 2907 4212 2916
rect 4160 2873 4169 2907
rect 4169 2873 4203 2907
rect 4203 2873 4212 2907
rect 4712 2907 4764 2916
rect 4160 2864 4212 2873
rect 4712 2873 4721 2907
rect 4721 2873 4755 2907
rect 4755 2873 4764 2907
rect 4712 2864 4764 2873
rect 9496 2932 9548 2984
rect 10692 2932 10744 2984
rect 16028 3068 16080 3120
rect 17316 3136 17368 3188
rect 18052 3136 18104 3188
rect 8484 2907 8536 2916
rect 8484 2873 8493 2907
rect 8493 2873 8527 2907
rect 8527 2873 8536 2907
rect 8484 2864 8536 2873
rect 9404 2864 9456 2916
rect 2228 2839 2280 2848
rect 2228 2805 2237 2839
rect 2237 2805 2271 2839
rect 2271 2805 2280 2839
rect 2228 2796 2280 2805
rect 4620 2796 4672 2848
rect 6184 2839 6236 2848
rect 6184 2805 6193 2839
rect 6193 2805 6227 2839
rect 6227 2805 6236 2839
rect 6184 2796 6236 2805
rect 7840 2839 7892 2848
rect 7840 2805 7849 2839
rect 7849 2805 7883 2839
rect 7883 2805 7892 2839
rect 7840 2796 7892 2805
rect 10784 2864 10836 2916
rect 14372 2839 14424 2848
rect 14372 2805 14381 2839
rect 14381 2805 14415 2839
rect 14415 2805 14424 2839
rect 14372 2796 14424 2805
rect 18604 2839 18656 2848
rect 18604 2805 18613 2839
rect 18613 2805 18647 2839
rect 18647 2805 18656 2839
rect 18604 2796 18656 2805
rect 8982 2694 9034 2746
rect 9046 2694 9098 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 17174 2694 17226 2746
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 5356 2635 5408 2644
rect 5356 2601 5365 2635
rect 5365 2601 5399 2635
rect 5399 2601 5408 2635
rect 5356 2592 5408 2601
rect 6460 2592 6512 2644
rect 3148 2524 3200 2576
rect 4712 2524 4764 2576
rect 8484 2592 8536 2644
rect 11980 2635 12032 2644
rect 11980 2601 11989 2635
rect 11989 2601 12023 2635
rect 12023 2601 12032 2635
rect 11980 2592 12032 2601
rect 10784 2524 10836 2576
rect 11152 2567 11204 2576
rect 11152 2533 11161 2567
rect 11161 2533 11195 2567
rect 11195 2533 11204 2567
rect 11152 2524 11204 2533
rect 14004 2524 14056 2576
rect 1032 2252 1084 2304
rect 2228 2456 2280 2508
rect 2136 2295 2188 2304
rect 2136 2261 2145 2295
rect 2145 2261 2179 2295
rect 2179 2261 2188 2295
rect 6000 2456 6052 2508
rect 12532 2456 12584 2508
rect 13636 2456 13688 2508
rect 16948 2456 17000 2508
rect 19984 2499 20036 2508
rect 3976 2388 4028 2440
rect 4344 2431 4396 2440
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 7656 2431 7708 2440
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 19984 2465 19993 2499
rect 19993 2465 20027 2499
rect 20027 2465 20036 2499
rect 19984 2456 20036 2465
rect 13268 2320 13320 2372
rect 12808 2295 12860 2304
rect 2136 2252 2188 2261
rect 12808 2261 12817 2295
rect 12817 2261 12851 2295
rect 12851 2261 12860 2295
rect 12808 2252 12860 2261
rect 15936 2252 15988 2304
rect 20076 2252 20128 2304
rect 21548 2252 21600 2304
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 12982 2150 13034 2202
rect 13046 2150 13098 2202
rect 13110 2150 13162 2202
rect 13174 2150 13226 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 8024 2048 8076 2100
rect 13452 2048 13504 2100
rect 7840 1912 7892 1964
rect 10232 1912 10284 1964
<< metal2 >>
rect 20 23588 72 23594
rect 20 23530 72 23536
rect 846 23588 902 24000
rect 846 23536 848 23588
rect 900 23536 902 23588
rect 32 6458 60 23530
rect 846 23520 902 23536
rect 2502 23610 2558 24000
rect 4250 23610 4306 24000
rect 5906 23610 5962 24000
rect 7654 23610 7710 24000
rect 9402 23610 9458 24000
rect 11058 23610 11114 24000
rect 2502 23582 2820 23610
rect 2502 23520 2558 23582
rect 860 23499 888 23520
rect 110 23352 166 23361
rect 110 23287 166 23296
rect 124 21010 152 23287
rect 1214 21720 1270 21729
rect 1214 21655 1270 21664
rect 112 21004 164 21010
rect 112 20946 164 20952
rect 1228 20398 1256 21655
rect 1582 20496 1638 20505
rect 1582 20431 1638 20440
rect 1216 20392 1268 20398
rect 1216 20334 1268 20340
rect 1596 20058 1624 20431
rect 1952 20256 2004 20262
rect 1952 20198 2004 20204
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1308 19916 1360 19922
rect 1308 19858 1360 19864
rect 1320 19174 1348 19858
rect 1582 19544 1638 19553
rect 1582 19479 1638 19488
rect 1596 19446 1624 19479
rect 1584 19440 1636 19446
rect 1584 19382 1636 19388
rect 1308 19168 1360 19174
rect 1308 19110 1360 19116
rect 112 18964 164 18970
rect 112 18906 164 18912
rect 124 18873 152 18906
rect 110 18864 166 18873
rect 110 18799 166 18808
rect 110 11928 166 11937
rect 110 11863 166 11872
rect 124 11830 152 11863
rect 112 11824 164 11830
rect 112 11766 164 11772
rect 110 10840 166 10849
rect 110 10775 166 10784
rect 124 10742 152 10775
rect 112 10736 164 10742
rect 112 10678 164 10684
rect 110 9752 166 9761
rect 110 9687 166 9696
rect 124 9654 152 9687
rect 112 9648 164 9654
rect 112 9590 164 9596
rect 1320 7818 1348 19110
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1688 17542 1716 18022
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1688 17202 1716 17478
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1768 17128 1820 17134
rect 1582 17096 1638 17105
rect 1768 17070 1820 17076
rect 1582 17031 1638 17040
rect 1596 16250 1624 17031
rect 1780 16794 1808 17070
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1412 15366 1440 15982
rect 1964 15706 1992 20198
rect 2792 19922 2820 23582
rect 4250 23582 4568 23610
rect 4250 23520 4306 23582
rect 4540 20602 4568 23582
rect 5906 23582 6132 23610
rect 5906 23520 5962 23582
rect 4956 21788 5252 21808
rect 5012 21786 5036 21788
rect 5092 21786 5116 21788
rect 5172 21786 5196 21788
rect 5034 21734 5036 21786
rect 5098 21734 5110 21786
rect 5172 21734 5174 21786
rect 5012 21732 5036 21734
rect 5092 21732 5116 21734
rect 5172 21732 5196 21734
rect 4956 21712 5252 21732
rect 4956 20700 5252 20720
rect 5012 20698 5036 20700
rect 5092 20698 5116 20700
rect 5172 20698 5196 20700
rect 5034 20646 5036 20698
rect 5098 20646 5110 20698
rect 5172 20646 5174 20698
rect 5012 20644 5036 20646
rect 5092 20644 5116 20646
rect 5172 20644 5196 20646
rect 4956 20624 5252 20644
rect 6104 20602 6132 23582
rect 7392 23582 7710 23610
rect 7392 20602 7420 23582
rect 7654 23520 7710 23582
rect 9324 23582 9458 23610
rect 8956 21244 9252 21264
rect 9012 21242 9036 21244
rect 9092 21242 9116 21244
rect 9172 21242 9196 21244
rect 9034 21190 9036 21242
rect 9098 21190 9110 21242
rect 9172 21190 9174 21242
rect 9012 21188 9036 21190
rect 9092 21188 9116 21190
rect 9172 21188 9196 21190
rect 8956 21168 9252 21188
rect 9324 20602 9352 23582
rect 9402 23520 9458 23582
rect 10980 23582 11114 23610
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9968 20602 9996 20946
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 4528 20596 4580 20602
rect 4528 20538 4580 20544
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 4540 20398 4568 20538
rect 6104 20398 6132 20538
rect 7392 20398 7420 20538
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 3792 20256 3844 20262
rect 3792 20198 3844 20204
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2792 19514 2820 19858
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2044 19168 2096 19174
rect 2044 19110 2096 19116
rect 2056 18970 2084 19110
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 2056 18290 2084 18906
rect 2596 18828 2648 18834
rect 2596 18770 2648 18776
rect 2504 18352 2556 18358
rect 2504 18294 2556 18300
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2516 18154 2544 18294
rect 2504 18148 2556 18154
rect 2504 18090 2556 18096
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 2044 16992 2096 16998
rect 2044 16934 2096 16940
rect 2056 16726 2084 16934
rect 2044 16720 2096 16726
rect 2044 16662 2096 16668
rect 2056 15910 2084 16662
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1400 15360 1452 15366
rect 1400 15302 1452 15308
rect 1964 15026 1992 15642
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 1860 14544 1912 14550
rect 1860 14486 1912 14492
rect 1872 14074 1900 14486
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 1872 13530 1900 14010
rect 2056 13802 2084 15846
rect 2148 14793 2176 18022
rect 2320 17808 2372 17814
rect 2320 17750 2372 17756
rect 2332 17134 2360 17750
rect 2516 17678 2544 18090
rect 2608 18086 2636 18770
rect 3436 18290 3464 19654
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 3436 17882 3464 18226
rect 3528 18154 3556 18702
rect 3516 18148 3568 18154
rect 3516 18090 3568 18096
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2320 17128 2372 17134
rect 2320 17070 2372 17076
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2884 16590 2912 16730
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2884 16250 2912 16526
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2976 15638 3004 15914
rect 2964 15632 3016 15638
rect 2964 15574 3016 15580
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2134 14784 2190 14793
rect 2134 14719 2190 14728
rect 2332 14346 2360 14962
rect 2596 14884 2648 14890
rect 2596 14826 2648 14832
rect 2608 14346 2636 14826
rect 2700 14618 2728 15438
rect 2976 15162 3004 15574
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2320 14340 2372 14346
rect 2320 14282 2372 14288
rect 2596 14340 2648 14346
rect 2596 14282 2648 14288
rect 2332 13938 2360 14282
rect 2608 14074 2636 14282
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2608 13870 2636 14010
rect 2700 14006 2728 14554
rect 2688 14000 2740 14006
rect 2688 13942 2740 13948
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2044 13796 2096 13802
rect 2044 13738 2096 13744
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 2056 12714 2084 13738
rect 3252 13530 3280 15438
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3528 13814 3556 15302
rect 3620 14890 3648 15982
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3608 14884 3660 14890
rect 3608 14826 3660 14832
rect 3712 14074 3740 15098
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3712 13870 3740 14010
rect 3700 13864 3752 13870
rect 3528 13786 3648 13814
rect 3700 13806 3752 13812
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 2688 13456 2740 13462
rect 2740 13416 2820 13444
rect 2688 13398 2740 13404
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 1490 12608 1546 12617
rect 1490 12543 1546 12552
rect 1504 11234 1532 12543
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1964 11286 1992 12174
rect 2056 11898 2084 12310
rect 2332 12170 2360 13262
rect 2412 12708 2464 12714
rect 2412 12650 2464 12656
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 1479 11218 1532 11234
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 1467 11212 1532 11218
rect 1519 11160 1532 11212
rect 1467 11154 1532 11160
rect 1504 10810 1532 11154
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1688 10266 1716 10542
rect 2148 10266 2176 11086
rect 2332 11082 2360 12106
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 2228 11008 2280 11014
rect 2228 10950 2280 10956
rect 2240 10606 2268 10950
rect 2424 10810 2452 12650
rect 2792 12646 2820 13416
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3344 12986 3372 13262
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3436 12782 3464 13466
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2792 12306 2820 12582
rect 3436 12442 3464 12718
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2700 11626 2728 11766
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 2700 11354 2728 11562
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2596 11280 2648 11286
rect 2596 11222 2648 11228
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2608 10742 2636 11222
rect 2780 11144 2832 11150
rect 2884 11132 2912 11494
rect 2832 11104 2912 11132
rect 2964 11144 3016 11150
rect 2780 11086 2832 11092
rect 2964 11086 3016 11092
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 1400 9988 1452 9994
rect 1400 9930 1452 9936
rect 1412 9518 1440 9930
rect 2148 9722 2176 9998
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2608 9586 2636 10134
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2884 9518 2912 10678
rect 2976 10198 3004 11086
rect 3160 10606 3188 11562
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3068 10266 3096 10542
rect 3436 10470 3464 10746
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2884 9178 2912 9454
rect 2976 9178 3004 10134
rect 3528 10062 3556 11494
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3620 9178 3648 13786
rect 3712 13462 3740 13806
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3804 9110 3832 20198
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 4956 19612 5252 19632
rect 5012 19610 5036 19612
rect 5092 19610 5116 19612
rect 5172 19610 5196 19612
rect 5034 19558 5036 19610
rect 5098 19558 5110 19610
rect 5172 19558 5174 19610
rect 5012 19556 5036 19558
rect 5092 19556 5116 19558
rect 5172 19556 5196 19558
rect 4956 19536 5252 19556
rect 5644 19174 5672 19858
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 4344 18828 4396 18834
rect 4344 18770 4396 18776
rect 4356 18426 4384 18770
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 4816 18426 4844 18634
rect 4956 18524 5252 18544
rect 5012 18522 5036 18524
rect 5092 18522 5116 18524
rect 5172 18522 5196 18524
rect 5034 18470 5036 18522
rect 5098 18470 5110 18522
rect 5172 18470 5174 18522
rect 5012 18468 5036 18470
rect 5092 18468 5116 18470
rect 5172 18468 5196 18470
rect 4956 18448 5252 18468
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 4080 17610 4108 18090
rect 4356 17814 4384 18362
rect 5644 18154 5672 19110
rect 5632 18148 5684 18154
rect 5632 18090 5684 18096
rect 4344 17808 4396 17814
rect 4344 17750 4396 17756
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 4080 16726 4108 17546
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 3884 16652 3936 16658
rect 3884 16594 3936 16600
rect 3896 15910 3924 16594
rect 4172 16454 4200 17138
rect 4264 16998 4292 17614
rect 4356 17338 4384 17750
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 4956 17436 5252 17456
rect 5012 17434 5036 17436
rect 5092 17434 5116 17436
rect 5172 17434 5196 17436
rect 5034 17382 5036 17434
rect 5098 17382 5110 17434
rect 5172 17382 5174 17434
rect 5012 17380 5036 17382
rect 5092 17380 5116 17382
rect 5172 17380 5196 17382
rect 4956 17360 5252 17380
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 5920 16998 5948 17614
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 13326 3924 15846
rect 4172 15706 4200 16390
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4264 15586 4292 16934
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4172 15558 4292 15586
rect 4356 15570 4384 15982
rect 4724 15910 4752 16594
rect 4956 16348 5252 16368
rect 5012 16346 5036 16348
rect 5092 16346 5116 16348
rect 5172 16346 5196 16348
rect 5034 16294 5036 16346
rect 5098 16294 5110 16346
rect 5172 16294 5174 16346
rect 5012 16292 5036 16294
rect 5092 16292 5116 16294
rect 5172 16292 5196 16294
rect 4956 16272 5252 16292
rect 5460 16046 5488 16594
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 5828 16114 5856 16390
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5722 16008 5778 16017
rect 5264 15972 5316 15978
rect 5920 15994 5948 16934
rect 5722 15943 5778 15952
rect 5828 15966 5948 15994
rect 5264 15914 5316 15920
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4724 15570 4752 15846
rect 5276 15706 5304 15914
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 4344 15564 4396 15570
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 14929 4108 14962
rect 4066 14920 4122 14929
rect 4066 14855 4122 14864
rect 4080 14550 4108 14855
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3988 13546 4016 13738
rect 4080 13734 4108 14350
rect 4172 13814 4200 15558
rect 4344 15506 4396 15512
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 4356 15162 4384 15506
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4632 15094 4660 15438
rect 4724 15162 4752 15506
rect 4956 15260 5252 15280
rect 5012 15258 5036 15260
rect 5092 15258 5116 15260
rect 5172 15258 5196 15260
rect 5034 15206 5036 15258
rect 5098 15206 5110 15258
rect 5172 15206 5174 15258
rect 5012 15204 5036 15206
rect 5092 15204 5116 15206
rect 5172 15204 5196 15206
rect 4956 15184 5252 15204
rect 5460 15162 5488 15506
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4264 14618 4292 14962
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 4172 13786 4292 13814
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4160 13728 4212 13734
rect 4160 13670 4212 13676
rect 4172 13546 4200 13670
rect 3988 13518 4200 13546
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3896 12986 3924 13126
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3896 12442 3924 12922
rect 4160 12708 4212 12714
rect 4160 12650 4212 12656
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3988 11665 4016 11698
rect 3974 11656 4030 11665
rect 3974 11591 4030 11600
rect 4172 11218 4200 12650
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4172 10198 4200 11154
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8362 1808 8774
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1780 8090 1808 8298
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1964 8022 1992 8978
rect 2240 8498 2268 8978
rect 4080 8498 4108 9658
rect 4172 9450 4200 9862
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 2240 8022 2268 8434
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 1952 8016 2004 8022
rect 1952 7958 2004 7964
rect 2228 8016 2280 8022
rect 2228 7958 2280 7964
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 1308 7812 1360 7818
rect 1308 7754 1360 7760
rect 112 7540 164 7546
rect 112 7482 164 7488
rect 124 7449 152 7482
rect 2148 7478 2176 7822
rect 2136 7472 2188 7478
rect 110 7440 166 7449
rect 2136 7414 2188 7420
rect 110 7375 166 7384
rect 1584 7268 1636 7274
rect 1584 7210 1636 7216
rect 1596 7002 1624 7210
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 2044 6928 2096 6934
rect 2044 6870 2096 6876
rect 2056 6730 2084 6870
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 20 6452 72 6458
rect 20 6394 72 6400
rect 1400 6180 1452 6186
rect 1400 6122 1452 6128
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1412 5642 1440 6122
rect 1688 5846 1716 6122
rect 1676 5840 1728 5846
rect 1676 5782 1728 5788
rect 1964 5778 1992 6598
rect 2056 6118 2084 6666
rect 2148 6390 2176 7414
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 2424 5914 2452 6802
rect 2516 6662 2544 7142
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1400 5636 1452 5642
rect 1400 5578 1452 5584
rect 1214 3496 1270 3505
rect 1214 3431 1270 3440
rect 1228 2990 1256 3431
rect 1412 3194 1440 5578
rect 1860 5092 1912 5098
rect 1860 5034 1912 5040
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1596 4593 1624 4626
rect 1582 4584 1638 4593
rect 1582 4519 1638 4528
rect 1596 4282 1624 4519
rect 1584 4276 1636 4282
rect 1584 4218 1636 4224
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 1216 2984 1268 2990
rect 1216 2926 1268 2932
rect 1032 2304 1084 2310
rect 1032 2246 1084 2252
rect 662 82 718 480
rect 1044 82 1072 2246
rect 1872 2009 1900 5034
rect 1964 4826 1992 5714
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2516 4154 2544 6054
rect 2608 5914 2636 8230
rect 2884 8090 2912 8230
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 3804 7954 3832 8230
rect 3988 8090 4016 8366
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2884 7002 2912 7142
rect 3804 7002 3832 7890
rect 3988 7750 4016 8026
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 2872 6996 2924 7002
rect 2872 6938 2924 6944
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3804 6458 3832 6802
rect 3896 6662 3924 7414
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3988 7206 4016 7346
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3792 6452 3844 6458
rect 3712 6412 3792 6440
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2884 5846 2912 6054
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3620 5137 3648 5170
rect 3606 5128 3662 5137
rect 3606 5063 3662 5072
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2700 4282 2728 4626
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2424 4126 2544 4154
rect 3160 4146 3188 4558
rect 3712 4282 3740 6412
rect 3792 6394 3844 6400
rect 3896 6390 3924 6598
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3804 5574 3832 6258
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3804 5370 3832 5510
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3148 4140 3200 4146
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2148 2310 2176 3878
rect 2332 3602 2360 3946
rect 2424 3924 2452 4126
rect 3148 4082 3200 4088
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 2596 3936 2648 3942
rect 2424 3896 2596 3924
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2240 2854 2268 3538
rect 2228 2848 2280 2854
rect 2228 2790 2280 2796
rect 2240 2514 2268 2790
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 1858 2000 1914 2009
rect 1858 1935 1914 1944
rect 2148 1193 2176 2246
rect 2134 1184 2190 1193
rect 2134 1119 2190 1128
rect 662 54 1072 82
rect 2042 82 2098 480
rect 2424 82 2452 3896
rect 2596 3878 2648 3884
rect 3712 3738 3740 4082
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2516 2990 2544 3334
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 3148 2916 3200 2922
rect 3148 2858 3200 2864
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3160 2582 3188 2858
rect 3528 2650 3556 2858
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 2042 54 2452 82
rect 3422 82 3478 480
rect 3804 82 3832 4966
rect 3896 4078 3924 6054
rect 3988 5030 4016 7142
rect 4080 6780 4108 8434
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4172 7177 4200 7210
rect 4158 7168 4214 7177
rect 4158 7103 4214 7112
rect 4160 6792 4212 6798
rect 4080 6752 4160 6780
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 4080 4690 4108 6752
rect 4160 6734 4212 6740
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4172 5234 4200 5714
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3988 3534 4016 4558
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3988 2446 4016 3470
rect 4172 3194 4200 3878
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4172 2922 4200 3130
rect 4264 3126 4292 13786
rect 4356 13734 4384 14554
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4540 13376 4568 13806
rect 4620 13388 4672 13394
rect 4540 13348 4620 13376
rect 4620 13330 4672 13336
rect 4632 12986 4660 13330
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4356 10810 4384 12854
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4540 11830 4568 12786
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4632 11898 4660 12242
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4528 11824 4580 11830
rect 4528 11766 4580 11772
rect 4540 11370 4568 11766
rect 4540 11342 4660 11370
rect 4724 11354 4752 15098
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 5000 14618 5028 14758
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4956 14172 5252 14192
rect 5012 14170 5036 14172
rect 5092 14170 5116 14172
rect 5172 14170 5196 14172
rect 5034 14118 5036 14170
rect 5098 14118 5110 14170
rect 5172 14118 5174 14170
rect 5012 14116 5036 14118
rect 5092 14116 5116 14118
rect 5172 14116 5196 14118
rect 4956 14096 5252 14116
rect 5736 13870 5764 15943
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 4956 13084 5252 13104
rect 5012 13082 5036 13084
rect 5092 13082 5116 13084
rect 5172 13082 5196 13084
rect 5034 13030 5036 13082
rect 5098 13030 5110 13082
rect 5172 13030 5174 13082
rect 5012 13028 5036 13030
rect 5092 13028 5116 13030
rect 5172 13028 5196 13030
rect 4956 13008 5252 13028
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5368 12170 5396 12582
rect 5736 12238 5764 12582
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 4956 11996 5252 12016
rect 5012 11994 5036 11996
rect 5092 11994 5116 11996
rect 5172 11994 5196 11996
rect 5034 11942 5036 11994
rect 5098 11942 5110 11994
rect 5172 11942 5174 11994
rect 5012 11940 5036 11942
rect 5092 11940 5116 11942
rect 5172 11940 5196 11942
rect 4956 11920 5252 11940
rect 5644 11694 5672 12038
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4448 10742 4476 11154
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4436 10736 4488 10742
rect 4436 10678 4488 10684
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4356 9722 4384 10066
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 4356 6730 4384 7958
rect 4448 7274 4476 10678
rect 4540 9450 4568 10950
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4436 7268 4488 7274
rect 4436 7210 4488 7216
rect 4540 7206 4568 7686
rect 4632 7410 4660 11342
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5460 11014 5488 11086
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 4724 10810 4752 10950
rect 4956 10908 5252 10928
rect 5012 10906 5036 10908
rect 5092 10906 5116 10908
rect 5172 10906 5196 10908
rect 5034 10854 5036 10906
rect 5098 10854 5110 10906
rect 5172 10854 5174 10906
rect 5012 10852 5036 10854
rect 5092 10852 5116 10854
rect 5172 10852 5196 10854
rect 4956 10832 5252 10852
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 5460 10674 5488 10950
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4816 10130 4844 10406
rect 5000 10266 5028 10474
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4804 10124 4856 10130
rect 5460 10112 5488 10474
rect 5552 10266 5580 10678
rect 5644 10470 5672 11630
rect 5736 11218 5764 12038
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5736 10130 5764 10474
rect 5724 10124 5776 10130
rect 5460 10084 5580 10112
rect 4804 10066 4856 10072
rect 4816 9722 4844 10066
rect 5552 9926 5580 10084
rect 5724 10066 5776 10072
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 4956 9820 5252 9840
rect 5012 9818 5036 9820
rect 5092 9818 5116 9820
rect 5172 9818 5196 9820
rect 5034 9766 5036 9818
rect 5098 9766 5110 9818
rect 5172 9766 5174 9818
rect 5012 9764 5036 9766
rect 5092 9764 5116 9766
rect 5172 9764 5196 9766
rect 4956 9744 5252 9764
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5000 9178 5028 9454
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5368 9110 5396 9318
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 4956 8732 5252 8752
rect 5012 8730 5036 8732
rect 5092 8730 5116 8732
rect 5172 8730 5196 8732
rect 5034 8678 5036 8730
rect 5098 8678 5110 8730
rect 5172 8678 5174 8730
rect 5012 8676 5036 8678
rect 5092 8676 5116 8678
rect 5172 8676 5196 8678
rect 4956 8656 5252 8676
rect 5368 8634 5396 9046
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4724 7750 4752 8434
rect 5460 8362 5488 9454
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4540 6866 4568 7142
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4540 5914 4568 6802
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4356 4826 4384 5510
rect 4540 5370 4568 5646
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4632 5137 4660 7210
rect 4618 5128 4674 5137
rect 4618 5063 4674 5072
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4620 4752 4672 4758
rect 4620 4694 4672 4700
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4540 4282 4568 4626
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4540 3670 4568 3946
rect 4632 3738 4660 4694
rect 4724 4554 4752 7686
rect 4956 7644 5252 7664
rect 5012 7642 5036 7644
rect 5092 7642 5116 7644
rect 5172 7642 5196 7644
rect 5034 7590 5036 7642
rect 5098 7590 5110 7642
rect 5172 7590 5174 7642
rect 5012 7588 5036 7590
rect 5092 7588 5116 7590
rect 5172 7588 5196 7590
rect 4956 7568 5252 7588
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4816 5760 4844 7414
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5184 6730 5212 7142
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 4956 6556 5252 6576
rect 5012 6554 5036 6556
rect 5092 6554 5116 6556
rect 5172 6554 5196 6556
rect 5034 6502 5036 6554
rect 5098 6502 5110 6554
rect 5172 6502 5174 6554
rect 5012 6500 5036 6502
rect 5092 6500 5116 6502
rect 5172 6500 5196 6502
rect 4956 6480 5252 6500
rect 5552 6458 5580 9862
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5644 8090 5672 8910
rect 5736 8838 5764 10066
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5736 7970 5764 8774
rect 5644 7942 5764 7970
rect 5644 7206 5672 7942
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5736 7546 5764 7754
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5632 7200 5684 7206
rect 5630 7168 5632 7177
rect 5684 7168 5686 7177
rect 5630 7103 5686 7112
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5460 5778 5488 6122
rect 5448 5772 5500 5778
rect 4816 5732 4936 5760
rect 4802 5672 4858 5681
rect 4908 5642 4936 5732
rect 5448 5714 5500 5720
rect 4802 5607 4858 5616
rect 4896 5636 4948 5642
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4816 4078 4844 5607
rect 4896 5578 4948 5584
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 4956 5468 5252 5488
rect 5012 5466 5036 5468
rect 5092 5466 5116 5468
rect 5172 5466 5196 5468
rect 5034 5414 5036 5466
rect 5098 5414 5110 5466
rect 5172 5414 5174 5466
rect 5012 5412 5036 5414
rect 5092 5412 5116 5414
rect 5172 5412 5196 5414
rect 4956 5392 5252 5412
rect 4986 5264 5042 5273
rect 5368 5234 5396 5510
rect 5460 5370 5488 5714
rect 5644 5574 5672 7103
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5540 5296 5592 5302
rect 5644 5273 5672 5510
rect 5540 5238 5592 5244
rect 5630 5264 5686 5273
rect 4986 5199 5042 5208
rect 5356 5228 5408 5234
rect 5000 5166 5028 5199
rect 5356 5170 5408 5176
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5000 4622 5028 5102
rect 5552 4826 5580 5238
rect 5630 5199 5686 5208
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5644 4690 5672 4966
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 4956 4380 5252 4400
rect 5012 4378 5036 4380
rect 5092 4378 5116 4380
rect 5172 4378 5196 4380
rect 5034 4326 5036 4378
rect 5098 4326 5110 4378
rect 5172 4326 5174 4378
rect 5012 4324 5036 4326
rect 5092 4324 5116 4326
rect 5172 4324 5196 4326
rect 4956 4304 5252 4324
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 4160 2916 4212 2922
rect 4160 2858 4212 2864
rect 4356 2446 4384 3334
rect 4632 2854 4660 3538
rect 4816 3058 4844 3878
rect 5368 3602 5396 4558
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 4956 3292 5252 3312
rect 5012 3290 5036 3292
rect 5092 3290 5116 3292
rect 5172 3290 5196 3292
rect 5034 3238 5036 3290
rect 5098 3238 5110 3290
rect 5172 3238 5174 3290
rect 5012 3236 5036 3238
rect 5092 3236 5116 3238
rect 5172 3236 5196 3238
rect 4956 3216 5252 3236
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 3422 54 3832 82
rect 4632 82 4660 2790
rect 4724 2582 4752 2858
rect 5368 2650 5396 3538
rect 5460 3194 5488 3606
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5736 3097 5764 6190
rect 5828 3194 5856 15966
rect 6288 15065 6316 20198
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6472 19514 6500 19654
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6472 19174 6500 19450
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6656 18766 6684 20198
rect 8956 20156 9252 20176
rect 9012 20154 9036 20156
rect 9092 20154 9116 20156
rect 9172 20154 9196 20156
rect 9034 20102 9036 20154
rect 9098 20102 9110 20154
rect 9172 20102 9174 20154
rect 9012 20100 9036 20102
rect 9092 20100 9116 20102
rect 9172 20100 9196 20102
rect 8956 20080 9252 20100
rect 9416 20058 9444 20198
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 10244 19990 10272 20742
rect 10980 20602 11008 23582
rect 11058 23520 11114 23582
rect 12806 23520 12862 24000
rect 14554 23610 14610 24000
rect 16210 23610 16266 24000
rect 17958 23610 18014 24000
rect 19706 23610 19762 24000
rect 21362 23610 21418 24000
rect 23110 23610 23166 24000
rect 14292 23582 14610 23610
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 10980 20398 11008 20538
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 10232 19984 10284 19990
rect 10232 19926 10284 19932
rect 11336 19984 11388 19990
rect 11336 19926 11388 19932
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 10060 19718 10088 19858
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 6736 18896 6788 18902
rect 6736 18838 6788 18844
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6656 18290 6684 18702
rect 6748 18426 6776 18838
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6460 17808 6512 17814
rect 6460 17750 6512 17756
rect 6472 17202 6500 17750
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6748 17134 6776 18362
rect 6932 18290 6960 18702
rect 7576 18290 7604 19178
rect 8956 19068 9252 19088
rect 9012 19066 9036 19068
rect 9092 19066 9116 19068
rect 9172 19066 9196 19068
rect 9034 19014 9036 19066
rect 9098 19014 9110 19066
rect 9172 19014 9174 19066
rect 9012 19012 9036 19014
rect 9092 19012 9116 19014
rect 9172 19012 9196 19014
rect 8956 18992 9252 19012
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 6932 17882 6960 18226
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6748 16794 6776 17070
rect 6368 16788 6420 16794
rect 6368 16730 6420 16736
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6380 16096 6408 16730
rect 6644 16108 6696 16114
rect 6380 16068 6644 16096
rect 6380 15910 6408 16068
rect 6644 16050 6696 16056
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6380 15638 6408 15846
rect 6368 15632 6420 15638
rect 6368 15574 6420 15580
rect 5998 15056 6054 15065
rect 5998 14991 6054 15000
rect 6274 15056 6330 15065
rect 6274 14991 6330 15000
rect 6012 14958 6040 14991
rect 6000 14952 6052 14958
rect 6000 14894 6052 14900
rect 6380 14822 6408 15574
rect 6472 14822 6500 15846
rect 6932 15570 6960 15846
rect 7024 15706 7052 18090
rect 8772 17882 8800 18566
rect 9140 18426 9168 18702
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9416 18290 9444 18566
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 8956 17980 9252 18000
rect 9012 17978 9036 17980
rect 9092 17978 9116 17980
rect 9172 17978 9196 17980
rect 9034 17926 9036 17978
rect 9098 17926 9110 17978
rect 9172 17926 9174 17978
rect 9012 17924 9036 17926
rect 9092 17924 9116 17926
rect 9172 17924 9196 17926
rect 8956 17904 9252 17924
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 8772 17270 8800 17818
rect 9416 17610 9444 18226
rect 9508 18154 9536 19246
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 9784 18902 9812 19178
rect 9772 18896 9824 18902
rect 9772 18838 9824 18844
rect 9784 18426 9812 18838
rect 10060 18766 10088 19654
rect 10244 19514 10272 19926
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 11348 19310 11376 19926
rect 12544 19854 12572 20198
rect 12624 19984 12676 19990
rect 12624 19926 12676 19932
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12544 19514 12572 19790
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12636 19378 12664 19926
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 10060 18290 10088 18702
rect 11348 18630 11376 19246
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12452 18970 12480 19110
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9416 17270 9444 17546
rect 9508 17542 9536 18090
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 9312 17060 9364 17066
rect 9312 17002 9364 17008
rect 8956 16892 9252 16912
rect 9012 16890 9036 16892
rect 9092 16890 9116 16892
rect 9172 16890 9196 16892
rect 9034 16838 9036 16890
rect 9098 16838 9110 16890
rect 9172 16838 9174 16890
rect 9012 16836 9036 16838
rect 9092 16836 9116 16838
rect 9172 16836 9196 16838
rect 8956 16816 9252 16836
rect 9324 16726 9352 17002
rect 9784 16998 9812 17750
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9876 17202 9904 17614
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10244 17105 10272 17138
rect 10230 17096 10286 17105
rect 10230 17031 10286 17040
rect 10692 17060 10744 17066
rect 10692 17002 10744 17008
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 9312 16720 9364 16726
rect 9312 16662 9364 16668
rect 9784 16658 9812 16934
rect 10152 16794 10180 16934
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 8128 16250 8156 16594
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 8588 16114 8616 16526
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 7300 15434 7328 15982
rect 8588 15706 8616 16050
rect 8680 16046 8708 16594
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8680 15570 8708 15982
rect 9508 15910 9536 16594
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 8956 15804 9252 15824
rect 9012 15802 9036 15804
rect 9092 15802 9116 15804
rect 9172 15802 9196 15804
rect 9034 15750 9036 15802
rect 9098 15750 9110 15802
rect 9172 15750 9174 15802
rect 9012 15748 9036 15750
rect 9092 15748 9116 15750
rect 9172 15748 9196 15750
rect 8956 15728 9252 15748
rect 9508 15706 9536 15846
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 6736 15428 6788 15434
rect 6736 15370 6788 15376
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6380 14550 6408 14758
rect 6368 14544 6420 14550
rect 6368 14486 6420 14492
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 5920 14074 5948 14350
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 5920 13530 5948 14010
rect 6380 13734 6408 14486
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 6104 12646 6132 13330
rect 6472 13326 6500 14758
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 5908 11620 5960 11626
rect 5908 11562 5960 11568
rect 5920 11150 5948 11562
rect 6104 11558 6132 12582
rect 6196 12306 6224 12718
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 6012 10810 6040 11222
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 9926 6040 10406
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 5920 8498 5948 9046
rect 6104 9042 6132 11494
rect 6196 10470 6224 12242
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6288 9926 6316 12854
rect 6472 12646 6500 13262
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6472 11914 6500 12582
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6564 12102 6592 12242
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6472 11886 6592 11914
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6380 10062 6408 10610
rect 6564 10198 6592 11886
rect 6656 11830 6684 12174
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6748 10198 6776 15370
rect 8036 14822 8064 15506
rect 8680 14822 8708 15506
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7484 13530 7512 13806
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12782 7328 13126
rect 7484 12850 7512 13466
rect 7944 13394 7972 13670
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7300 12170 7328 12718
rect 7944 12442 7972 13330
rect 8128 12986 8156 14350
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8496 12986 8524 13126
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8496 12646 8524 12922
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7012 11620 7064 11626
rect 7012 11562 7064 11568
rect 7024 11354 7052 11562
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7024 10606 7052 11290
rect 7116 11014 7144 12038
rect 7392 11626 7420 12038
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 8128 11286 8156 12174
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8312 11558 8340 12038
rect 8404 11762 8432 12174
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8404 11354 8432 11698
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8116 11280 8168 11286
rect 8116 11222 8168 11228
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7116 10810 7144 10950
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 7024 10266 7052 10542
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6564 10062 6592 10134
rect 7208 10130 7236 10950
rect 7392 10266 7420 11086
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8312 10470 8340 10950
rect 8588 10742 8616 12922
rect 8680 12442 8708 14758
rect 8956 14716 9252 14736
rect 9012 14714 9036 14716
rect 9092 14714 9116 14716
rect 9172 14714 9196 14716
rect 9034 14662 9036 14714
rect 9098 14662 9110 14714
rect 9172 14662 9174 14714
rect 9012 14660 9036 14662
rect 9092 14660 9116 14662
rect 9172 14660 9196 14662
rect 8956 14640 9252 14660
rect 10152 14482 10180 16730
rect 10704 16454 10732 17002
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10244 15162 10272 15914
rect 10336 15638 10364 15982
rect 10324 15632 10376 15638
rect 10324 15574 10376 15580
rect 10704 15366 10732 16390
rect 11256 16250 11284 17478
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10244 14890 10272 15098
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10232 14884 10284 14890
rect 10232 14826 10284 14832
rect 10336 14618 10364 14894
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 10152 14006 10180 14418
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 8956 13628 9252 13648
rect 9012 13626 9036 13628
rect 9092 13626 9116 13628
rect 9172 13626 9196 13628
rect 9034 13574 9036 13626
rect 9098 13574 9110 13626
rect 9172 13574 9174 13626
rect 9012 13572 9036 13574
rect 9092 13572 9116 13574
rect 9172 13572 9196 13574
rect 8956 13552 9252 13572
rect 9324 13530 9352 13874
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9968 12782 9996 13738
rect 10244 13734 10272 14350
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 10152 12714 10180 13466
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10428 12782 10456 13126
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 8956 12540 9252 12560
rect 9012 12538 9036 12540
rect 9092 12538 9116 12540
rect 9172 12538 9196 12540
rect 9034 12486 9036 12538
rect 9098 12486 9110 12538
rect 9172 12486 9174 12538
rect 9012 12484 9036 12486
rect 9092 12484 9116 12486
rect 9172 12484 9196 12486
rect 8956 12464 9252 12484
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 9600 12374 9628 12582
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 10244 12306 10272 12718
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 9126 12200 9182 12209
rect 9126 12135 9182 12144
rect 9140 12102 9168 12135
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9140 11626 9168 12038
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 8956 11452 9252 11472
rect 9012 11450 9036 11452
rect 9092 11450 9116 11452
rect 9172 11450 9196 11452
rect 9034 11398 9036 11450
rect 9098 11398 9110 11450
rect 9172 11398 9174 11450
rect 9012 11396 9036 11398
rect 9092 11396 9116 11398
rect 9172 11396 9196 11398
rect 8956 11376 9252 11396
rect 9416 11286 9444 12038
rect 9508 11626 9536 12242
rect 10336 12102 10364 12582
rect 10428 12238 10456 12718
rect 10520 12646 10548 13330
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9416 10810 9444 11222
rect 9508 11218 9536 11562
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9508 11014 9536 11154
rect 9692 11014 9720 11494
rect 10060 11286 10088 11834
rect 10244 11830 10272 12038
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8404 10266 8432 10474
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8496 10130 8524 10406
rect 8588 10198 8616 10678
rect 8956 10364 9252 10384
rect 9012 10362 9036 10364
rect 9092 10362 9116 10364
rect 9172 10362 9196 10364
rect 9034 10310 9036 10362
rect 9098 10310 9110 10362
rect 9172 10310 9174 10362
rect 9012 10308 9036 10310
rect 9092 10308 9116 10310
rect 9172 10308 9196 10310
rect 8956 10288 9252 10308
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6288 9722 6316 9862
rect 6380 9722 6408 9998
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6276 9716 6328 9722
rect 6196 9676 6276 9704
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 6012 6934 6040 7278
rect 6104 7002 6132 8978
rect 6196 7478 6224 9676
rect 6276 9658 6328 9664
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6472 9450 6500 9930
rect 8312 9722 8340 10066
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 6472 9178 6500 9386
rect 7208 9178 7236 9454
rect 8496 9450 8524 10066
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6288 7546 6316 7822
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6196 6458 6224 6802
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6380 6458 6408 6734
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6196 6254 6224 6394
rect 6472 6390 6500 9114
rect 7852 9042 7880 9386
rect 8772 9042 8800 9998
rect 8956 9276 9252 9296
rect 9012 9274 9036 9276
rect 9092 9274 9116 9276
rect 9172 9274 9196 9276
rect 9034 9222 9036 9274
rect 9098 9222 9110 9274
rect 9172 9222 9174 9274
rect 9012 9220 9036 9222
rect 9092 9220 9116 9222
rect 9172 9220 9196 9222
rect 8956 9200 9252 9220
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 7852 8634 7880 8978
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7300 8022 7328 8230
rect 7288 8016 7340 8022
rect 6734 7984 6790 7993
rect 7288 7958 7340 7964
rect 6734 7919 6790 7928
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 6012 4826 6040 5714
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6012 3738 6040 4762
rect 6196 4758 6224 5510
rect 6472 5370 6500 6326
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6472 5166 6500 5306
rect 6748 5166 6776 7919
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6840 7342 6868 7686
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6840 7002 6868 7278
rect 7300 7002 7328 7958
rect 7760 7546 7788 8366
rect 8128 8294 8156 8910
rect 8772 8634 8800 8978
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 8036 6934 8064 7482
rect 8024 6928 8076 6934
rect 8024 6870 8076 6876
rect 6920 6860 6972 6866
rect 6972 6820 7052 6848
rect 6920 6802 6972 6808
rect 7024 6662 7052 6820
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 6118 7052 6598
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7024 5846 7052 6054
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 7024 4826 7052 5782
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 6196 4282 6224 4694
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5722 3088 5778 3097
rect 5722 3023 5778 3032
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 6012 2514 6040 3674
rect 6472 3398 6500 4558
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6840 4078 6868 4422
rect 7484 4078 7512 6054
rect 7760 5710 7788 6190
rect 8036 5914 8064 6870
rect 8128 6118 8156 8230
rect 8956 8188 9252 8208
rect 9012 8186 9036 8188
rect 9092 8186 9116 8188
rect 9172 8186 9196 8188
rect 9034 8134 9036 8186
rect 9098 8134 9110 8186
rect 9172 8134 9174 8186
rect 9012 8132 9036 8134
rect 9092 8132 9116 8134
rect 9172 8132 9196 8134
rect 8956 8112 9252 8132
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8220 6798 8248 7822
rect 8760 7744 8812 7750
rect 8760 7686 8812 7692
rect 8772 7410 8800 7686
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 6840 3534 6868 4014
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7300 3602 7328 3878
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 4956 2204 5252 2224
rect 5012 2202 5036 2204
rect 5092 2202 5116 2204
rect 5172 2202 5196 2204
rect 5034 2150 5036 2202
rect 5098 2150 5110 2202
rect 5172 2150 5174 2202
rect 5012 2148 5036 2150
rect 5092 2148 5116 2150
rect 5172 2148 5196 2150
rect 4956 2128 5252 2148
rect 4894 82 4950 480
rect 4632 54 4950 82
rect 6196 82 6224 2790
rect 6472 2650 6500 3334
rect 7300 3194 7328 3538
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 7668 2446 7696 4490
rect 7760 4146 7788 4694
rect 7852 4690 7880 5510
rect 8220 5030 8248 5714
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7760 3738 7788 4082
rect 8128 3942 8156 4150
rect 8404 4010 8432 4626
rect 8588 4570 8616 5102
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8496 4542 8616 4570
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 8128 3670 8156 3878
rect 8496 3738 8524 4542
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8128 3194 8156 3606
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8496 2922 8524 3674
rect 8680 3602 8708 5034
rect 8772 4826 8800 7346
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 8956 7100 9252 7120
rect 9012 7098 9036 7100
rect 9092 7098 9116 7100
rect 9172 7098 9196 7100
rect 9034 7046 9036 7098
rect 9098 7046 9110 7098
rect 9172 7046 9174 7098
rect 9012 7044 9036 7046
rect 9092 7044 9116 7046
rect 9172 7044 9196 7046
rect 8956 7024 9252 7044
rect 9324 7002 9352 7210
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9324 6730 9352 6938
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 8956 6012 9252 6032
rect 9012 6010 9036 6012
rect 9092 6010 9116 6012
rect 9172 6010 9196 6012
rect 9034 5958 9036 6010
rect 9098 5958 9110 6010
rect 9172 5958 9174 6010
rect 9012 5956 9036 5958
rect 9092 5956 9116 5958
rect 9172 5956 9196 5958
rect 8956 5936 9252 5956
rect 9324 5914 9352 6666
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9416 5846 9444 10746
rect 9508 10266 9536 10950
rect 9692 10470 9720 10950
rect 10060 10742 10088 11222
rect 10152 11150 10180 11698
rect 10336 11558 10364 12038
rect 10428 11694 10456 12174
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10152 10810 10180 11086
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10048 10736 10100 10742
rect 10048 10678 10100 10684
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9692 10130 9720 10406
rect 10060 10266 10088 10678
rect 10520 10606 10548 12582
rect 10612 11898 10640 13670
rect 10704 12442 10732 15302
rect 10888 14890 10916 15506
rect 11348 15162 11376 18566
rect 11900 18426 11928 18702
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 12452 18358 12480 18906
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 12268 17814 12296 18022
rect 12256 17808 12308 17814
rect 12256 17750 12308 17756
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11532 16590 11560 17002
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11532 15706 11560 16526
rect 11900 15978 11928 16730
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 12072 15972 12124 15978
rect 12072 15914 12124 15920
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 12084 15162 12112 15914
rect 12452 15638 12480 15982
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 12084 14890 12112 15098
rect 12360 14958 12388 15302
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 10784 14340 10836 14346
rect 10784 14282 10836 14288
rect 10796 13870 10824 14282
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10796 13530 10824 13806
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10888 13462 10916 14826
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 14074 11100 14214
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10876 13456 10928 13462
rect 10876 13398 10928 13404
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10796 12986 10824 13330
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10796 12442 10824 12922
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10612 10606 10640 11834
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10796 11665 10824 11698
rect 10782 11656 10838 11665
rect 10782 11591 10838 11600
rect 11072 11286 11100 14010
rect 11900 13938 11928 14418
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11164 11898 11192 13874
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11532 13530 11560 13806
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11532 12986 11560 13466
rect 12084 13462 12112 14826
rect 12360 14550 12388 14894
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12176 14074 12204 14418
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 12084 12986 12112 13398
rect 12176 13394 12204 14010
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12636 12986 12664 13262
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 11520 12164 11572 12170
rect 11520 12106 11572 12112
rect 11532 11898 11560 12106
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 12084 11830 12112 12922
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12084 11286 12112 11766
rect 12452 11694 12480 12378
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11348 10674 11376 11086
rect 11532 10810 11560 11222
rect 12268 11014 12296 11222
rect 12728 11150 12756 19790
rect 12820 19514 12848 23520
rect 12956 21788 13252 21808
rect 13012 21786 13036 21788
rect 13092 21786 13116 21788
rect 13172 21786 13196 21788
rect 13034 21734 13036 21786
rect 13098 21734 13110 21786
rect 13172 21734 13174 21786
rect 13012 21732 13036 21734
rect 13092 21732 13116 21734
rect 13172 21732 13196 21734
rect 12956 21712 13252 21732
rect 12956 20700 13252 20720
rect 13012 20698 13036 20700
rect 13092 20698 13116 20700
rect 13172 20698 13196 20700
rect 13034 20646 13036 20698
rect 13098 20646 13110 20698
rect 13172 20646 13174 20698
rect 13012 20644 13036 20646
rect 13092 20644 13116 20646
rect 13172 20644 13196 20646
rect 12956 20624 13252 20644
rect 14292 20602 14320 23582
rect 14554 23520 14610 23582
rect 15856 23582 16266 23610
rect 15856 20602 15884 23582
rect 16210 23520 16266 23582
rect 17696 23582 18014 23610
rect 16956 21244 17252 21264
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17034 21190 17036 21242
rect 17098 21190 17110 21242
rect 17172 21190 17174 21242
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 16956 21168 17252 21188
rect 17696 20602 17724 23582
rect 17958 23520 18014 23582
rect 19444 23582 19762 23610
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 14556 20392 14608 20398
rect 14556 20334 14608 20340
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 12956 19612 13252 19632
rect 13012 19610 13036 19612
rect 13092 19610 13116 19612
rect 13172 19610 13196 19612
rect 13034 19558 13036 19610
rect 13098 19558 13110 19610
rect 13172 19558 13174 19610
rect 13012 19556 13036 19558
rect 13092 19556 13116 19558
rect 13172 19556 13196 19558
rect 12956 19536 13252 19556
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 12820 19310 12848 19450
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12820 18766 12848 19110
rect 12900 18896 12952 18902
rect 12900 18838 12952 18844
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12912 18612 12940 18838
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 12820 18584 12940 18612
rect 12820 18068 12848 18584
rect 12956 18524 13252 18544
rect 13012 18522 13036 18524
rect 13092 18522 13116 18524
rect 13172 18522 13196 18524
rect 13034 18470 13036 18522
rect 13098 18470 13110 18522
rect 13172 18470 13174 18522
rect 13012 18468 13036 18470
rect 13092 18468 13116 18470
rect 13172 18468 13196 18470
rect 12956 18448 13252 18468
rect 13280 18290 13308 18702
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 12900 18080 12952 18086
rect 12820 18040 12900 18068
rect 12900 18022 12952 18028
rect 12912 17746 12940 18022
rect 12900 17740 12952 17746
rect 12820 17700 12900 17728
rect 12820 17338 12848 17700
rect 12900 17682 12952 17688
rect 12956 17436 13252 17456
rect 13012 17434 13036 17436
rect 13092 17434 13116 17436
rect 13172 17434 13196 17436
rect 13034 17382 13036 17434
rect 13098 17382 13110 17434
rect 13172 17382 13174 17434
rect 13012 17380 13036 17382
rect 13092 17380 13116 17382
rect 13172 17380 13196 17382
rect 12956 17360 13252 17380
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12820 16794 12848 17274
rect 13280 17202 13308 18226
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 13004 16794 13032 16934
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 12956 16348 13252 16368
rect 13012 16346 13036 16348
rect 13092 16346 13116 16348
rect 13172 16346 13196 16348
rect 13034 16294 13036 16346
rect 13098 16294 13110 16346
rect 13172 16294 13174 16346
rect 13012 16292 13036 16294
rect 13092 16292 13116 16294
rect 13172 16292 13196 16294
rect 12956 16272 13252 16292
rect 13280 16182 13308 16934
rect 13268 16176 13320 16182
rect 13268 16118 13320 16124
rect 13372 15706 13400 20198
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13464 16250 13492 16662
rect 13648 16590 13676 17002
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13648 16046 13676 16526
rect 13740 16522 13768 17614
rect 14464 17060 14516 17066
rect 14464 17002 14516 17008
rect 14476 16726 14504 17002
rect 14464 16720 14516 16726
rect 14464 16662 14516 16668
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13740 16250 13768 16458
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 12956 15260 13252 15280
rect 13012 15258 13036 15260
rect 13092 15258 13116 15260
rect 13172 15258 13196 15260
rect 13034 15206 13036 15258
rect 13098 15206 13110 15258
rect 13172 15206 13174 15258
rect 13012 15204 13036 15206
rect 13092 15204 13116 15206
rect 13172 15204 13196 15206
rect 12956 15184 13252 15204
rect 13464 15094 13492 15370
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 13870 12848 14214
rect 12956 14172 13252 14192
rect 13012 14170 13036 14172
rect 13092 14170 13116 14172
rect 13172 14170 13196 14172
rect 13034 14118 13036 14170
rect 13098 14118 13110 14170
rect 13172 14118 13174 14170
rect 13012 14116 13036 14118
rect 13092 14116 13116 14118
rect 13172 14116 13196 14118
rect 12956 14096 13252 14116
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12820 13530 12848 13806
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12820 12986 12848 13466
rect 12956 13084 13252 13104
rect 13012 13082 13036 13084
rect 13092 13082 13116 13084
rect 13172 13082 13196 13084
rect 13034 13030 13036 13082
rect 13098 13030 13110 13082
rect 13172 13030 13174 13082
rect 13012 13028 13036 13030
rect 13092 13028 13116 13030
rect 13172 13028 13196 13030
rect 12956 13008 13252 13028
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 13280 12374 13308 13670
rect 13464 13530 13492 15030
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13464 12850 13492 13466
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 12956 11996 13252 12016
rect 13012 11994 13036 11996
rect 13092 11994 13116 11996
rect 13172 11994 13196 11996
rect 13034 11942 13036 11994
rect 13098 11942 13110 11994
rect 13172 11942 13174 11994
rect 13012 11940 13036 11942
rect 13092 11940 13116 11942
rect 13172 11940 13196 11942
rect 12956 11920 13252 11940
rect 13280 11830 13308 12310
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13372 11898 13400 12174
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13464 11558 13492 12582
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9692 9994 9720 10066
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9692 9382 9720 9930
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9968 9518 9996 9590
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9404 5840 9456 5846
rect 9404 5782 9456 5788
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8772 4146 8800 4422
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8772 3738 8800 4082
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8680 3058 8708 3538
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7668 1329 7696 2382
rect 7852 1970 7880 2790
rect 8496 2650 8524 2858
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8024 2100 8076 2106
rect 8024 2042 8076 2048
rect 7840 1964 7892 1970
rect 7840 1906 7892 1912
rect 7654 1320 7710 1329
rect 7654 1255 7710 1264
rect 6274 82 6330 480
rect 6196 54 6330 82
rect 662 0 718 54
rect 2042 0 2098 54
rect 3422 0 3478 54
rect 4894 0 4950 54
rect 6274 0 6330 54
rect 7654 82 7710 480
rect 8036 82 8064 2042
rect 7654 54 8064 82
rect 8864 82 8892 4966
rect 8956 4924 9252 4944
rect 9012 4922 9036 4924
rect 9092 4922 9116 4924
rect 9172 4922 9196 4924
rect 9034 4870 9036 4922
rect 9098 4870 9110 4922
rect 9172 4870 9174 4922
rect 9012 4868 9036 4870
rect 9092 4868 9116 4870
rect 9172 4868 9196 4870
rect 8956 4848 9252 4868
rect 8956 3836 9252 3856
rect 9012 3834 9036 3836
rect 9092 3834 9116 3836
rect 9172 3834 9196 3836
rect 9034 3782 9036 3834
rect 9098 3782 9110 3834
rect 9172 3782 9174 3834
rect 9012 3780 9036 3782
rect 9092 3780 9116 3782
rect 9172 3780 9196 3782
rect 8956 3760 9252 3780
rect 9324 3194 9352 5034
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9416 3126 9444 5578
rect 9508 5098 9536 5646
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9692 4154 9720 9318
rect 9784 9110 9812 9318
rect 9968 9178 9996 9454
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9968 8634 9996 9114
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9876 6934 9904 7278
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9876 6458 9904 6870
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9968 6186 9996 8570
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9968 5370 9996 5646
rect 10060 5642 10088 10202
rect 10520 9926 10548 10542
rect 10612 10266 10640 10542
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10520 9722 10548 9862
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 11532 9654 11560 10746
rect 12268 10130 12296 10950
rect 12728 10674 12756 10950
rect 12956 10908 13252 10928
rect 13012 10906 13036 10908
rect 13092 10906 13116 10908
rect 13172 10906 13196 10908
rect 13034 10854 13036 10906
rect 13098 10854 13110 10906
rect 13172 10854 13174 10906
rect 13012 10852 13036 10854
rect 13092 10852 13116 10854
rect 13172 10852 13196 10854
rect 12956 10832 13252 10852
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12544 10266 12572 10474
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10244 9450 10272 9522
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 10244 9178 10272 9386
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10244 7954 10272 9114
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10888 8498 10916 8774
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 11164 8362 11192 9386
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10336 8090 10364 8230
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 11164 8022 11192 8298
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10244 7546 10272 7890
rect 11716 7886 11744 9862
rect 12268 9722 12296 10066
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12728 9586 12756 10610
rect 13280 10266 13308 11086
rect 13372 10674 13400 11086
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13372 10130 13400 10610
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 12956 9820 13252 9840
rect 13012 9818 13036 9820
rect 13092 9818 13116 9820
rect 13172 9818 13196 9820
rect 13034 9766 13036 9818
rect 13098 9766 13110 9818
rect 13172 9766 13174 9818
rect 13012 9764 13036 9766
rect 13092 9764 13116 9766
rect 13172 9764 13196 9766
rect 12956 9744 13252 9764
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 13464 8956 13492 11494
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13556 10810 13584 11222
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13544 8968 13596 8974
rect 13464 8928 13544 8956
rect 13544 8910 13596 8916
rect 12956 8732 13252 8752
rect 13012 8730 13036 8732
rect 13092 8730 13116 8732
rect 13172 8730 13196 8732
rect 13034 8678 13036 8730
rect 13098 8678 13110 8730
rect 13172 8678 13174 8730
rect 13012 8676 13036 8678
rect 13092 8676 13116 8678
rect 13172 8676 13196 8678
rect 12956 8656 13252 8676
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11716 7546 11744 7822
rect 12084 7546 12112 7890
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 11704 7268 11756 7274
rect 11704 7210 11756 7216
rect 11716 7002 11744 7210
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11256 6322 11284 6734
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 10060 5370 10088 5578
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 9864 5296 9916 5302
rect 10060 5250 10088 5306
rect 9916 5244 10088 5250
rect 9864 5238 10088 5244
rect 9876 5222 10088 5238
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9784 4758 9812 5102
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 10428 4690 10456 5306
rect 10520 5234 10548 5646
rect 10784 5296 10836 5302
rect 10784 5238 10836 5244
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10796 4758 10824 5238
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 11072 4690 11100 6258
rect 11256 6225 11284 6258
rect 11242 6216 11298 6225
rect 11242 6151 11298 6160
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11440 5302 11468 5714
rect 11428 5296 11480 5302
rect 11428 5238 11480 5244
rect 11808 4758 11836 6054
rect 12084 5370 12112 7482
rect 12360 7002 12388 7822
rect 13556 7818 13584 8910
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12728 7274 12756 7686
rect 12956 7644 13252 7664
rect 13012 7642 13036 7644
rect 13092 7642 13116 7644
rect 13172 7642 13196 7644
rect 13034 7590 13036 7642
rect 13098 7590 13110 7642
rect 13172 7590 13174 7642
rect 13012 7588 13036 7590
rect 13092 7588 13116 7590
rect 13172 7588 13196 7590
rect 12956 7568 13252 7588
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12256 6928 12308 6934
rect 12256 6870 12308 6876
rect 12268 6186 12296 6870
rect 12360 6322 12388 6938
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12728 6322 12756 6666
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12256 6180 12308 6186
rect 12256 6122 12308 6128
rect 12268 5778 12296 6122
rect 12256 5772 12308 5778
rect 12256 5714 12308 5720
rect 12268 5370 12296 5714
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 10060 4282 10088 4626
rect 10428 4282 10456 4626
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11164 4282 11192 4558
rect 11808 4282 11836 4694
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 9692 4126 9812 4154
rect 10060 4146 10088 4218
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9416 2922 9444 3062
rect 9508 2990 9536 3606
rect 9496 2984 9548 2990
rect 9784 2961 9812 4126
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3670 10088 3878
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10060 3058 10088 3470
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10704 2990 10732 3606
rect 11164 3398 11192 4014
rect 11992 3534 12020 5034
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 10692 2984 10744 2990
rect 9496 2926 9548 2932
rect 9770 2952 9826 2961
rect 9404 2916 9456 2922
rect 10692 2926 10744 2932
rect 9770 2887 9826 2896
rect 10784 2916 10836 2922
rect 9404 2858 9456 2864
rect 10784 2858 10836 2864
rect 8956 2748 9252 2768
rect 9012 2746 9036 2748
rect 9092 2746 9116 2748
rect 9172 2746 9196 2748
rect 9034 2694 9036 2746
rect 9098 2694 9110 2746
rect 9172 2694 9174 2746
rect 9012 2692 9036 2694
rect 9092 2692 9116 2694
rect 9172 2692 9196 2694
rect 8956 2672 9252 2692
rect 10796 2582 10824 2858
rect 11164 2582 11192 3334
rect 11992 2650 12020 3470
rect 12084 3194 12112 3606
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 10232 1964 10284 1970
rect 10232 1906 10284 1912
rect 9126 82 9182 480
rect 8864 54 9182 82
rect 10244 82 10272 1906
rect 10506 82 10562 480
rect 10244 54 10562 82
rect 7654 0 7710 54
rect 9126 0 9182 54
rect 10506 0 10562 54
rect 11886 82 11942 480
rect 12176 82 12204 5102
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12268 3738 12296 4422
rect 12544 4146 12572 4626
rect 12728 4154 12756 6258
rect 12820 5914 12848 7142
rect 13464 6934 13492 7346
rect 13452 6928 13504 6934
rect 13452 6870 13504 6876
rect 12956 6556 13252 6576
rect 13012 6554 13036 6556
rect 13092 6554 13116 6556
rect 13172 6554 13196 6556
rect 13034 6502 13036 6554
rect 13098 6502 13110 6554
rect 13172 6502 13174 6554
rect 13012 6500 13036 6502
rect 13092 6500 13116 6502
rect 13172 6500 13196 6502
rect 12956 6480 13252 6500
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12956 5468 13252 5488
rect 13012 5466 13036 5468
rect 13092 5466 13116 5468
rect 13172 5466 13196 5468
rect 13034 5414 13036 5466
rect 13098 5414 13110 5466
rect 13172 5414 13174 5466
rect 13012 5412 13036 5414
rect 13092 5412 13116 5414
rect 13172 5412 13196 5414
rect 12956 5392 13252 5412
rect 13556 5166 13584 7754
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 12956 4380 13252 4400
rect 13012 4378 13036 4380
rect 13092 4378 13116 4380
rect 13172 4378 13196 4380
rect 13034 4326 13036 4378
rect 13098 4326 13110 4378
rect 13172 4326 13174 4378
rect 13012 4324 13036 4326
rect 13092 4324 13116 4326
rect 13172 4324 13196 4326
rect 12956 4304 13252 4324
rect 12728 4146 12848 4154
rect 12532 4140 12584 4146
rect 12728 4140 12860 4146
rect 12728 4126 12808 4140
rect 12532 4082 12584 4088
rect 12808 4082 12860 4088
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12544 2514 12572 3878
rect 12820 3670 12848 4082
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12912 3670 12940 3946
rect 13464 3942 13492 4626
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 12808 3664 12860 3670
rect 12808 3606 12860 3612
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 12956 3292 13252 3312
rect 13012 3290 13036 3292
rect 13092 3290 13116 3292
rect 13172 3290 13196 3292
rect 13034 3238 13036 3290
rect 13098 3238 13110 3290
rect 13172 3238 13174 3290
rect 13012 3236 13036 3238
rect 13092 3236 13116 3238
rect 13172 3236 13196 3238
rect 12956 3216 13252 3236
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12820 1193 12848 2246
rect 12956 2204 13252 2224
rect 13012 2202 13036 2204
rect 13092 2202 13116 2204
rect 13172 2202 13196 2204
rect 13034 2150 13036 2202
rect 13098 2150 13110 2202
rect 13172 2150 13174 2202
rect 13012 2148 13036 2150
rect 13092 2148 13116 2150
rect 13172 2148 13196 2150
rect 12956 2128 13252 2148
rect 12806 1184 12862 1193
rect 12806 1119 12862 1128
rect 11886 54 12204 82
rect 13280 82 13308 2314
rect 13464 2106 13492 3878
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13556 3194 13584 3538
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13648 2514 13676 15846
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13740 15162 13768 15574
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13740 14482 13768 15098
rect 14292 15026 14320 15642
rect 14476 15502 14504 16390
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 14550 14136 14758
rect 14476 14618 14504 15438
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13740 14074 13768 14418
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13740 12374 13768 12786
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13832 12238 13860 13262
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 14016 11694 14044 12038
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 14016 11354 14044 11630
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14016 10266 14044 11290
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13832 9722 13860 10066
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13740 8294 13768 8978
rect 13728 8288 13780 8294
rect 13728 8230 13780 8236
rect 13740 6254 13768 8230
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13832 4282 13860 6190
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 14108 4154 14136 9862
rect 14476 9042 14504 10610
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14568 7546 14596 20334
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 14936 14929 14964 20198
rect 16956 20156 17252 20176
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17034 20102 17036 20154
rect 17098 20102 17110 20154
rect 17172 20102 17174 20154
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 16956 20080 17252 20100
rect 16956 19068 17252 19088
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17034 19014 17036 19066
rect 17098 19014 17110 19066
rect 17172 19014 17174 19066
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 16956 18992 17252 19012
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 15382 17640 15438 17649
rect 15382 17575 15438 17584
rect 15396 16658 15424 17575
rect 16408 17105 16436 18566
rect 16956 17980 17252 18000
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17034 17926 17036 17978
rect 17098 17926 17110 17978
rect 17172 17926 17174 17978
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 16956 17904 17252 17924
rect 16394 17096 16450 17105
rect 16394 17031 16450 17040
rect 16956 16892 17252 16912
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17034 16838 17036 16890
rect 17098 16838 17110 16890
rect 17172 16838 17174 16890
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 16956 16816 17252 16836
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15396 16250 15424 16594
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 16956 15804 17252 15824
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17034 15750 17036 15802
rect 17098 15750 17110 15802
rect 17172 15750 17174 15802
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 16956 15728 17252 15748
rect 16670 15056 16726 15065
rect 16670 14991 16726 15000
rect 14922 14920 14978 14929
rect 14922 14855 14978 14864
rect 16684 14414 16712 14991
rect 16956 14716 17252 14736
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17034 14662 17036 14714
rect 17098 14662 17110 14714
rect 17172 14662 17174 14714
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 16956 14640 17252 14660
rect 16764 14544 16816 14550
rect 16764 14486 16816 14492
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15488 13938 15516 14214
rect 16684 14006 16712 14350
rect 16776 14074 16804 14486
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 14740 13796 14792 13802
rect 14740 13738 14792 13744
rect 14752 12764 14780 13738
rect 14832 12776 14884 12782
rect 14752 12736 14832 12764
rect 14752 12442 14780 12736
rect 14832 12718 14884 12724
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 15212 12306 15240 13874
rect 15488 13814 15516 13874
rect 15396 13786 15516 13814
rect 15396 12850 15424 13786
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15948 13462 15976 13670
rect 16776 13530 16804 14010
rect 16956 13628 17252 13648
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17034 13574 17036 13626
rect 17098 13574 17110 13626
rect 17172 13574 17174 13626
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 16956 13552 17252 13572
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 15936 13456 15988 13462
rect 15936 13398 15988 13404
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15488 12442 15516 13262
rect 15948 12646 15976 13398
rect 16776 12986 16804 13466
rect 17328 13326 17356 14350
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17420 13462 17448 13670
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17420 12986 17448 13398
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 16776 12782 16804 12922
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15212 11898 15240 12242
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15212 10674 15240 11834
rect 15948 11626 15976 12582
rect 16956 12540 17252 12560
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17034 12486 17036 12538
rect 17098 12486 17110 12538
rect 17172 12486 17174 12538
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 16956 12464 17252 12484
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16684 11898 16712 12242
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 15936 11620 15988 11626
rect 15936 11562 15988 11568
rect 15948 11354 15976 11562
rect 16956 11452 17252 11472
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17034 11398 17036 11450
rect 17098 11398 17110 11450
rect 17172 11398 17174 11450
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 16956 11376 17252 11396
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15580 10674 15608 11086
rect 15948 10810 15976 11290
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17420 11014 17448 11222
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17420 10810 17448 10950
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15120 10266 15148 10542
rect 16956 10364 17252 10384
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17034 10310 17036 10362
rect 17098 10310 17110 10362
rect 17172 10310 17174 10362
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 16956 10288 17252 10308
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 17420 10130 17448 10746
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17420 9654 17448 10066
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 16956 9276 17252 9296
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17034 9222 17036 9274
rect 17098 9222 17110 9274
rect 17172 9222 17174 9274
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 16956 9200 17252 9220
rect 16956 8188 17252 8208
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17034 8134 17036 8186
rect 17098 8134 17110 8186
rect 17172 8134 17174 8186
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 16956 8112 17252 8132
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 16956 7100 17252 7120
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17034 7046 17036 7098
rect 17098 7046 17110 7098
rect 17172 7046 17174 7098
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 16956 7024 17252 7044
rect 14464 6248 14516 6254
rect 17328 6225 17356 7142
rect 14464 6190 14516 6196
rect 17314 6216 17370 6225
rect 14476 5914 14504 6190
rect 15108 6180 15160 6186
rect 17314 6151 17370 6160
rect 15108 6122 15160 6128
rect 15120 5914 15148 6122
rect 16956 6012 17252 6032
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17034 5958 17036 6010
rect 17098 5958 17110 6010
rect 17172 5958 17174 6010
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 16956 5936 17252 5956
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 14476 5710 14504 5850
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14476 5166 14504 5646
rect 15580 5234 15608 5850
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14200 4826 14228 5102
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14384 4826 14412 5034
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14016 4126 14136 4154
rect 14384 4146 14412 4762
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14372 4140 14424 4146
rect 14016 2582 14044 4126
rect 14372 4082 14424 4088
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 14004 2576 14056 2582
rect 14004 2518 14056 2524
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 13452 2100 13504 2106
rect 13452 2042 13504 2048
rect 13358 82 13414 480
rect 13280 54 13414 82
rect 14384 82 14412 2790
rect 14660 1737 14688 4218
rect 15396 4010 15424 4966
rect 16500 4758 16528 4966
rect 16956 4924 17252 4944
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17034 4870 17036 4922
rect 17098 4870 17110 4922
rect 17172 4870 17174 4922
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 16956 4848 17252 4868
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 17224 4752 17276 4758
rect 17224 4694 17276 4700
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15580 3670 15608 4422
rect 16132 4214 16160 4626
rect 17236 4282 17264 4694
rect 17224 4276 17276 4282
rect 17276 4236 17356 4264
rect 17224 4218 17276 4224
rect 16120 4208 16172 4214
rect 16120 4150 16172 4156
rect 16132 4010 16160 4150
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16316 3670 16344 4082
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15752 3664 15804 3670
rect 15752 3606 15804 3612
rect 16028 3664 16080 3670
rect 16028 3606 16080 3612
rect 16304 3664 16356 3670
rect 16304 3606 16356 3612
rect 15764 3194 15792 3606
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 16040 3126 16068 3606
rect 16408 3534 16436 3878
rect 16956 3836 17252 3856
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17034 3782 17036 3834
rect 17098 3782 17110 3834
rect 17172 3782 17174 3834
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 16956 3760 17252 3780
rect 17328 3602 17356 4236
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16132 3194 16160 3470
rect 17328 3194 17356 3538
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 16956 2748 17252 2768
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17034 2694 17036 2746
rect 17098 2694 17110 2746
rect 17172 2694 17174 2746
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 16956 2672 17252 2692
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 15936 2304 15988 2310
rect 15936 2246 15988 2252
rect 14646 1728 14702 1737
rect 14646 1663 14702 1672
rect 14738 82 14794 480
rect 14384 54 14794 82
rect 15948 82 15976 2246
rect 16960 1329 16988 2450
rect 16946 1320 17002 1329
rect 16946 1255 17002 1264
rect 16118 82 16174 480
rect 15948 54 16174 82
rect 17420 82 17448 9318
rect 17512 4622 17540 20198
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 17868 19712 17920 19718
rect 17868 19654 17920 19660
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17696 11558 17724 12242
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17696 6361 17724 11494
rect 17880 11150 17908 19654
rect 18708 19242 18736 19858
rect 19444 19514 19472 23582
rect 19706 23520 19762 23582
rect 21284 23582 21418 23610
rect 20956 21788 21252 21808
rect 21012 21786 21036 21788
rect 21092 21786 21116 21788
rect 21172 21786 21196 21788
rect 21034 21734 21036 21786
rect 21098 21734 21110 21786
rect 21172 21734 21174 21786
rect 21012 21732 21036 21734
rect 21092 21732 21116 21734
rect 21172 21732 21196 21734
rect 20956 21712 21252 21732
rect 20956 20700 21252 20720
rect 21012 20698 21036 20700
rect 21092 20698 21116 20700
rect 21172 20698 21196 20700
rect 21034 20646 21036 20698
rect 21098 20646 21110 20698
rect 21172 20646 21174 20698
rect 21012 20644 21036 20646
rect 21092 20644 21116 20646
rect 21172 20644 21196 20646
rect 20956 20624 21252 20644
rect 21284 20602 21312 23582
rect 21362 23520 21418 23582
rect 22848 23582 23166 23610
rect 21454 22128 21510 22137
rect 21454 22063 21510 22072
rect 21468 20602 21496 22063
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21468 20398 21496 20538
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 18696 19236 18748 19242
rect 18696 19178 18748 19184
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 19890 14920 19946 14929
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 18064 13462 18092 14010
rect 18432 13802 18460 14214
rect 18524 13802 18552 14894
rect 19890 14855 19946 14864
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19720 14482 19748 14758
rect 19904 14618 19932 14855
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 18800 14074 18828 14418
rect 19720 14074 19748 14418
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 18800 13462 18828 13738
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18708 12918 18736 13262
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18156 12442 18184 12786
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11830 18460 12038
rect 18420 11824 18472 11830
rect 18420 11766 18472 11772
rect 18432 11626 18460 11766
rect 18708 11626 18736 12174
rect 18984 11762 19012 12174
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 18328 11620 18380 11626
rect 18328 11562 18380 11568
rect 18420 11620 18472 11626
rect 18420 11562 18472 11568
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18340 11286 18368 11562
rect 18328 11280 18380 11286
rect 18328 11222 18380 11228
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17880 10742 17908 11086
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 18340 10674 18368 11222
rect 18432 11218 18460 11562
rect 18708 11354 18736 11562
rect 19444 11558 19472 12310
rect 20640 12209 20668 20198
rect 21270 19816 21326 19825
rect 21270 19751 21326 19760
rect 20956 19612 21252 19632
rect 21012 19610 21036 19612
rect 21092 19610 21116 19612
rect 21172 19610 21196 19612
rect 21034 19558 21036 19610
rect 21098 19558 21110 19610
rect 21172 19558 21174 19610
rect 21012 19556 21036 19558
rect 21092 19556 21116 19558
rect 21172 19556 21196 19558
rect 20956 19536 21252 19556
rect 21284 18834 21312 19751
rect 22848 19242 22876 23582
rect 23110 23520 23166 23582
rect 22836 19236 22888 19242
rect 22836 19178 22888 19184
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 20956 18524 21252 18544
rect 21012 18522 21036 18524
rect 21092 18522 21116 18524
rect 21172 18522 21196 18524
rect 21034 18470 21036 18522
rect 21098 18470 21110 18522
rect 21172 18470 21174 18522
rect 21012 18468 21036 18470
rect 21092 18468 21116 18470
rect 21172 18468 21196 18470
rect 20956 18448 21252 18468
rect 21284 18426 21312 18770
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 20956 17436 21252 17456
rect 21012 17434 21036 17436
rect 21092 17434 21116 17436
rect 21172 17434 21196 17436
rect 21034 17382 21036 17434
rect 21098 17382 21110 17434
rect 21172 17382 21174 17434
rect 21012 17380 21036 17382
rect 21092 17380 21116 17382
rect 21172 17380 21196 17382
rect 20956 17360 21252 17380
rect 20956 16348 21252 16368
rect 21012 16346 21036 16348
rect 21092 16346 21116 16348
rect 21172 16346 21196 16348
rect 21034 16294 21036 16346
rect 21098 16294 21110 16346
rect 21172 16294 21174 16346
rect 21012 16292 21036 16294
rect 21092 16292 21116 16294
rect 21172 16292 21196 16294
rect 20956 16272 21252 16292
rect 20956 15260 21252 15280
rect 21012 15258 21036 15260
rect 21092 15258 21116 15260
rect 21172 15258 21196 15260
rect 21034 15206 21036 15258
rect 21098 15206 21110 15258
rect 21172 15206 21174 15258
rect 21012 15204 21036 15206
rect 21092 15204 21116 15206
rect 21172 15204 21196 15206
rect 20956 15184 21252 15204
rect 20956 14172 21252 14192
rect 21012 14170 21036 14172
rect 21092 14170 21116 14172
rect 21172 14170 21196 14172
rect 21034 14118 21036 14170
rect 21098 14118 21110 14170
rect 21172 14118 21174 14170
rect 21012 14116 21036 14118
rect 21092 14116 21116 14118
rect 21172 14116 21196 14118
rect 20956 14096 21252 14116
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 21086 12608 21142 12617
rect 21086 12543 21142 12552
rect 21100 12442 21128 12543
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20626 12200 20682 12209
rect 20626 12135 20682 12144
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19444 11354 19472 11494
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 20732 11218 20760 12106
rect 20824 11830 20852 12242
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 19168 10810 19196 11154
rect 20732 10810 20760 11154
rect 23572 11008 23624 11014
rect 23572 10950 23624 10956
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 23584 10713 23612 10950
rect 23570 10704 23626 10713
rect 18328 10668 18380 10674
rect 23570 10639 23626 10648
rect 18328 10610 18380 10616
rect 18144 10532 18196 10538
rect 18064 10492 18144 10520
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17788 10198 17816 10406
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 18064 9926 18092 10492
rect 18144 10474 18196 10480
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 18064 9722 18092 9862
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19260 7546 19288 7890
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 21454 7712 21510 7721
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 17682 6352 17738 6361
rect 17682 6287 17738 6296
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 17512 3738 17540 4558
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 18064 3942 18092 4422
rect 18432 4146 18460 4558
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17788 3670 17816 3878
rect 17776 3664 17828 3670
rect 17776 3606 17828 3612
rect 18064 3194 18092 3878
rect 18248 3670 18276 3946
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18432 3534 18460 4082
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 17590 82 17646 480
rect 17420 54 17646 82
rect 18616 82 18644 2790
rect 19996 2514 20024 7686
rect 20956 7644 21252 7664
rect 21454 7647 21510 7656
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21468 7546 21496 7647
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21468 7342 21496 7482
rect 21456 7336 21508 7342
rect 21456 7278 21508 7284
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 21548 2304 21600 2310
rect 21548 2246 21600 2252
rect 18970 82 19026 480
rect 18616 54 19026 82
rect 20088 82 20116 2246
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 20350 82 20406 480
rect 20088 54 20406 82
rect 21560 82 21588 2246
rect 23294 1184 23350 1193
rect 23294 1119 23350 1128
rect 21822 82 21878 480
rect 21560 54 21878 82
rect 11886 0 11942 54
rect 13358 0 13414 54
rect 14738 0 14794 54
rect 16118 0 16174 54
rect 17590 0 17646 54
rect 18970 0 19026 54
rect 20350 0 20406 54
rect 21822 0 21878 54
rect 23202 82 23258 480
rect 23308 82 23336 1119
rect 23202 54 23336 82
rect 23202 0 23258 54
<< via2 >>
rect 110 23296 166 23352
rect 1214 21664 1270 21720
rect 1582 20440 1638 20496
rect 1582 19488 1638 19544
rect 110 18808 166 18864
rect 110 11872 166 11928
rect 110 10784 166 10840
rect 110 9696 166 9752
rect 1582 17040 1638 17096
rect 4956 21786 5012 21788
rect 5036 21786 5092 21788
rect 5116 21786 5172 21788
rect 5196 21786 5252 21788
rect 4956 21734 4982 21786
rect 4982 21734 5012 21786
rect 5036 21734 5046 21786
rect 5046 21734 5092 21786
rect 5116 21734 5162 21786
rect 5162 21734 5172 21786
rect 5196 21734 5226 21786
rect 5226 21734 5252 21786
rect 4956 21732 5012 21734
rect 5036 21732 5092 21734
rect 5116 21732 5172 21734
rect 5196 21732 5252 21734
rect 4956 20698 5012 20700
rect 5036 20698 5092 20700
rect 5116 20698 5172 20700
rect 5196 20698 5252 20700
rect 4956 20646 4982 20698
rect 4982 20646 5012 20698
rect 5036 20646 5046 20698
rect 5046 20646 5092 20698
rect 5116 20646 5162 20698
rect 5162 20646 5172 20698
rect 5196 20646 5226 20698
rect 5226 20646 5252 20698
rect 4956 20644 5012 20646
rect 5036 20644 5092 20646
rect 5116 20644 5172 20646
rect 5196 20644 5252 20646
rect 8956 21242 9012 21244
rect 9036 21242 9092 21244
rect 9116 21242 9172 21244
rect 9196 21242 9252 21244
rect 8956 21190 8982 21242
rect 8982 21190 9012 21242
rect 9036 21190 9046 21242
rect 9046 21190 9092 21242
rect 9116 21190 9162 21242
rect 9162 21190 9172 21242
rect 9196 21190 9226 21242
rect 9226 21190 9252 21242
rect 8956 21188 9012 21190
rect 9036 21188 9092 21190
rect 9116 21188 9172 21190
rect 9196 21188 9252 21190
rect 2134 14728 2190 14784
rect 1490 12552 1546 12608
rect 4956 19610 5012 19612
rect 5036 19610 5092 19612
rect 5116 19610 5172 19612
rect 5196 19610 5252 19612
rect 4956 19558 4982 19610
rect 4982 19558 5012 19610
rect 5036 19558 5046 19610
rect 5046 19558 5092 19610
rect 5116 19558 5162 19610
rect 5162 19558 5172 19610
rect 5196 19558 5226 19610
rect 5226 19558 5252 19610
rect 4956 19556 5012 19558
rect 5036 19556 5092 19558
rect 5116 19556 5172 19558
rect 5196 19556 5252 19558
rect 4956 18522 5012 18524
rect 5036 18522 5092 18524
rect 5116 18522 5172 18524
rect 5196 18522 5252 18524
rect 4956 18470 4982 18522
rect 4982 18470 5012 18522
rect 5036 18470 5046 18522
rect 5046 18470 5092 18522
rect 5116 18470 5162 18522
rect 5162 18470 5172 18522
rect 5196 18470 5226 18522
rect 5226 18470 5252 18522
rect 4956 18468 5012 18470
rect 5036 18468 5092 18470
rect 5116 18468 5172 18470
rect 5196 18468 5252 18470
rect 4956 17434 5012 17436
rect 5036 17434 5092 17436
rect 5116 17434 5172 17436
rect 5196 17434 5252 17436
rect 4956 17382 4982 17434
rect 4982 17382 5012 17434
rect 5036 17382 5046 17434
rect 5046 17382 5092 17434
rect 5116 17382 5162 17434
rect 5162 17382 5172 17434
rect 5196 17382 5226 17434
rect 5226 17382 5252 17434
rect 4956 17380 5012 17382
rect 5036 17380 5092 17382
rect 5116 17380 5172 17382
rect 5196 17380 5252 17382
rect 4956 16346 5012 16348
rect 5036 16346 5092 16348
rect 5116 16346 5172 16348
rect 5196 16346 5252 16348
rect 4956 16294 4982 16346
rect 4982 16294 5012 16346
rect 5036 16294 5046 16346
rect 5046 16294 5092 16346
rect 5116 16294 5162 16346
rect 5162 16294 5172 16346
rect 5196 16294 5226 16346
rect 5226 16294 5252 16346
rect 4956 16292 5012 16294
rect 5036 16292 5092 16294
rect 5116 16292 5172 16294
rect 5196 16292 5252 16294
rect 5722 15952 5778 16008
rect 4066 14864 4122 14920
rect 4956 15258 5012 15260
rect 5036 15258 5092 15260
rect 5116 15258 5172 15260
rect 5196 15258 5252 15260
rect 4956 15206 4982 15258
rect 4982 15206 5012 15258
rect 5036 15206 5046 15258
rect 5046 15206 5092 15258
rect 5116 15206 5162 15258
rect 5162 15206 5172 15258
rect 5196 15206 5226 15258
rect 5226 15206 5252 15258
rect 4956 15204 5012 15206
rect 5036 15204 5092 15206
rect 5116 15204 5172 15206
rect 5196 15204 5252 15206
rect 3974 11600 4030 11656
rect 110 7384 166 7440
rect 1214 3440 1270 3496
rect 1582 4528 1638 4584
rect 3606 5072 3662 5128
rect 1858 1944 1914 2000
rect 2134 1128 2190 1184
rect 4158 7112 4214 7168
rect 4956 14170 5012 14172
rect 5036 14170 5092 14172
rect 5116 14170 5172 14172
rect 5196 14170 5252 14172
rect 4956 14118 4982 14170
rect 4982 14118 5012 14170
rect 5036 14118 5046 14170
rect 5046 14118 5092 14170
rect 5116 14118 5162 14170
rect 5162 14118 5172 14170
rect 5196 14118 5226 14170
rect 5226 14118 5252 14170
rect 4956 14116 5012 14118
rect 5036 14116 5092 14118
rect 5116 14116 5172 14118
rect 5196 14116 5252 14118
rect 4956 13082 5012 13084
rect 5036 13082 5092 13084
rect 5116 13082 5172 13084
rect 5196 13082 5252 13084
rect 4956 13030 4982 13082
rect 4982 13030 5012 13082
rect 5036 13030 5046 13082
rect 5046 13030 5092 13082
rect 5116 13030 5162 13082
rect 5162 13030 5172 13082
rect 5196 13030 5226 13082
rect 5226 13030 5252 13082
rect 4956 13028 5012 13030
rect 5036 13028 5092 13030
rect 5116 13028 5172 13030
rect 5196 13028 5252 13030
rect 4956 11994 5012 11996
rect 5036 11994 5092 11996
rect 5116 11994 5172 11996
rect 5196 11994 5252 11996
rect 4956 11942 4982 11994
rect 4982 11942 5012 11994
rect 5036 11942 5046 11994
rect 5046 11942 5092 11994
rect 5116 11942 5162 11994
rect 5162 11942 5172 11994
rect 5196 11942 5226 11994
rect 5226 11942 5252 11994
rect 4956 11940 5012 11942
rect 5036 11940 5092 11942
rect 5116 11940 5172 11942
rect 5196 11940 5252 11942
rect 4956 10906 5012 10908
rect 5036 10906 5092 10908
rect 5116 10906 5172 10908
rect 5196 10906 5252 10908
rect 4956 10854 4982 10906
rect 4982 10854 5012 10906
rect 5036 10854 5046 10906
rect 5046 10854 5092 10906
rect 5116 10854 5162 10906
rect 5162 10854 5172 10906
rect 5196 10854 5226 10906
rect 5226 10854 5252 10906
rect 4956 10852 5012 10854
rect 5036 10852 5092 10854
rect 5116 10852 5172 10854
rect 5196 10852 5252 10854
rect 4956 9818 5012 9820
rect 5036 9818 5092 9820
rect 5116 9818 5172 9820
rect 5196 9818 5252 9820
rect 4956 9766 4982 9818
rect 4982 9766 5012 9818
rect 5036 9766 5046 9818
rect 5046 9766 5092 9818
rect 5116 9766 5162 9818
rect 5162 9766 5172 9818
rect 5196 9766 5226 9818
rect 5226 9766 5252 9818
rect 4956 9764 5012 9766
rect 5036 9764 5092 9766
rect 5116 9764 5172 9766
rect 5196 9764 5252 9766
rect 4956 8730 5012 8732
rect 5036 8730 5092 8732
rect 5116 8730 5172 8732
rect 5196 8730 5252 8732
rect 4956 8678 4982 8730
rect 4982 8678 5012 8730
rect 5036 8678 5046 8730
rect 5046 8678 5092 8730
rect 5116 8678 5162 8730
rect 5162 8678 5172 8730
rect 5196 8678 5226 8730
rect 5226 8678 5252 8730
rect 4956 8676 5012 8678
rect 5036 8676 5092 8678
rect 5116 8676 5172 8678
rect 5196 8676 5252 8678
rect 4618 5072 4674 5128
rect 4956 7642 5012 7644
rect 5036 7642 5092 7644
rect 5116 7642 5172 7644
rect 5196 7642 5252 7644
rect 4956 7590 4982 7642
rect 4982 7590 5012 7642
rect 5036 7590 5046 7642
rect 5046 7590 5092 7642
rect 5116 7590 5162 7642
rect 5162 7590 5172 7642
rect 5196 7590 5226 7642
rect 5226 7590 5252 7642
rect 4956 7588 5012 7590
rect 5036 7588 5092 7590
rect 5116 7588 5172 7590
rect 5196 7588 5252 7590
rect 4956 6554 5012 6556
rect 5036 6554 5092 6556
rect 5116 6554 5172 6556
rect 5196 6554 5252 6556
rect 4956 6502 4982 6554
rect 4982 6502 5012 6554
rect 5036 6502 5046 6554
rect 5046 6502 5092 6554
rect 5116 6502 5162 6554
rect 5162 6502 5172 6554
rect 5196 6502 5226 6554
rect 5226 6502 5252 6554
rect 4956 6500 5012 6502
rect 5036 6500 5092 6502
rect 5116 6500 5172 6502
rect 5196 6500 5252 6502
rect 5630 7148 5632 7168
rect 5632 7148 5684 7168
rect 5684 7148 5686 7168
rect 5630 7112 5686 7148
rect 4802 5616 4858 5672
rect 4956 5466 5012 5468
rect 5036 5466 5092 5468
rect 5116 5466 5172 5468
rect 5196 5466 5252 5468
rect 4956 5414 4982 5466
rect 4982 5414 5012 5466
rect 5036 5414 5046 5466
rect 5046 5414 5092 5466
rect 5116 5414 5162 5466
rect 5162 5414 5172 5466
rect 5196 5414 5226 5466
rect 5226 5414 5252 5466
rect 4956 5412 5012 5414
rect 5036 5412 5092 5414
rect 5116 5412 5172 5414
rect 5196 5412 5252 5414
rect 4986 5208 5042 5264
rect 5630 5208 5686 5264
rect 4956 4378 5012 4380
rect 5036 4378 5092 4380
rect 5116 4378 5172 4380
rect 5196 4378 5252 4380
rect 4956 4326 4982 4378
rect 4982 4326 5012 4378
rect 5036 4326 5046 4378
rect 5046 4326 5092 4378
rect 5116 4326 5162 4378
rect 5162 4326 5172 4378
rect 5196 4326 5226 4378
rect 5226 4326 5252 4378
rect 4956 4324 5012 4326
rect 5036 4324 5092 4326
rect 5116 4324 5172 4326
rect 5196 4324 5252 4326
rect 4956 3290 5012 3292
rect 5036 3290 5092 3292
rect 5116 3290 5172 3292
rect 5196 3290 5252 3292
rect 4956 3238 4982 3290
rect 4982 3238 5012 3290
rect 5036 3238 5046 3290
rect 5046 3238 5092 3290
rect 5116 3238 5162 3290
rect 5162 3238 5172 3290
rect 5196 3238 5226 3290
rect 5226 3238 5252 3290
rect 4956 3236 5012 3238
rect 5036 3236 5092 3238
rect 5116 3236 5172 3238
rect 5196 3236 5252 3238
rect 8956 20154 9012 20156
rect 9036 20154 9092 20156
rect 9116 20154 9172 20156
rect 9196 20154 9252 20156
rect 8956 20102 8982 20154
rect 8982 20102 9012 20154
rect 9036 20102 9046 20154
rect 9046 20102 9092 20154
rect 9116 20102 9162 20154
rect 9162 20102 9172 20154
rect 9196 20102 9226 20154
rect 9226 20102 9252 20154
rect 8956 20100 9012 20102
rect 9036 20100 9092 20102
rect 9116 20100 9172 20102
rect 9196 20100 9252 20102
rect 8956 19066 9012 19068
rect 9036 19066 9092 19068
rect 9116 19066 9172 19068
rect 9196 19066 9252 19068
rect 8956 19014 8982 19066
rect 8982 19014 9012 19066
rect 9036 19014 9046 19066
rect 9046 19014 9092 19066
rect 9116 19014 9162 19066
rect 9162 19014 9172 19066
rect 9196 19014 9226 19066
rect 9226 19014 9252 19066
rect 8956 19012 9012 19014
rect 9036 19012 9092 19014
rect 9116 19012 9172 19014
rect 9196 19012 9252 19014
rect 5998 15000 6054 15056
rect 6274 15000 6330 15056
rect 8956 17978 9012 17980
rect 9036 17978 9092 17980
rect 9116 17978 9172 17980
rect 9196 17978 9252 17980
rect 8956 17926 8982 17978
rect 8982 17926 9012 17978
rect 9036 17926 9046 17978
rect 9046 17926 9092 17978
rect 9116 17926 9162 17978
rect 9162 17926 9172 17978
rect 9196 17926 9226 17978
rect 9226 17926 9252 17978
rect 8956 17924 9012 17926
rect 9036 17924 9092 17926
rect 9116 17924 9172 17926
rect 9196 17924 9252 17926
rect 8956 16890 9012 16892
rect 9036 16890 9092 16892
rect 9116 16890 9172 16892
rect 9196 16890 9252 16892
rect 8956 16838 8982 16890
rect 8982 16838 9012 16890
rect 9036 16838 9046 16890
rect 9046 16838 9092 16890
rect 9116 16838 9162 16890
rect 9162 16838 9172 16890
rect 9196 16838 9226 16890
rect 9226 16838 9252 16890
rect 8956 16836 9012 16838
rect 9036 16836 9092 16838
rect 9116 16836 9172 16838
rect 9196 16836 9252 16838
rect 10230 17040 10286 17096
rect 8956 15802 9012 15804
rect 9036 15802 9092 15804
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 8956 15750 8982 15802
rect 8982 15750 9012 15802
rect 9036 15750 9046 15802
rect 9046 15750 9092 15802
rect 9116 15750 9162 15802
rect 9162 15750 9172 15802
rect 9196 15750 9226 15802
rect 9226 15750 9252 15802
rect 8956 15748 9012 15750
rect 9036 15748 9092 15750
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 8956 14714 9012 14716
rect 9036 14714 9092 14716
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 8956 14662 8982 14714
rect 8982 14662 9012 14714
rect 9036 14662 9046 14714
rect 9046 14662 9092 14714
rect 9116 14662 9162 14714
rect 9162 14662 9172 14714
rect 9196 14662 9226 14714
rect 9226 14662 9252 14714
rect 8956 14660 9012 14662
rect 9036 14660 9092 14662
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 8956 13626 9012 13628
rect 9036 13626 9092 13628
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 8956 13574 8982 13626
rect 8982 13574 9012 13626
rect 9036 13574 9046 13626
rect 9046 13574 9092 13626
rect 9116 13574 9162 13626
rect 9162 13574 9172 13626
rect 9196 13574 9226 13626
rect 9226 13574 9252 13626
rect 8956 13572 9012 13574
rect 9036 13572 9092 13574
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 8956 12538 9012 12540
rect 9036 12538 9092 12540
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 8956 12486 8982 12538
rect 8982 12486 9012 12538
rect 9036 12486 9046 12538
rect 9046 12486 9092 12538
rect 9116 12486 9162 12538
rect 9162 12486 9172 12538
rect 9196 12486 9226 12538
rect 9226 12486 9252 12538
rect 8956 12484 9012 12486
rect 9036 12484 9092 12486
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 9126 12144 9182 12200
rect 8956 11450 9012 11452
rect 9036 11450 9092 11452
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 8956 11398 8982 11450
rect 8982 11398 9012 11450
rect 9036 11398 9046 11450
rect 9046 11398 9092 11450
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9252 11450
rect 8956 11396 9012 11398
rect 9036 11396 9092 11398
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 8956 10362 9012 10364
rect 9036 10362 9092 10364
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 8956 10310 8982 10362
rect 8982 10310 9012 10362
rect 9036 10310 9046 10362
rect 9046 10310 9092 10362
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9252 10362
rect 8956 10308 9012 10310
rect 9036 10308 9092 10310
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 8956 9274 9012 9276
rect 9036 9274 9092 9276
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 8956 9222 8982 9274
rect 8982 9222 9012 9274
rect 9036 9222 9046 9274
rect 9046 9222 9092 9274
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9252 9274
rect 8956 9220 9012 9222
rect 9036 9220 9092 9222
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 6734 7928 6790 7984
rect 5722 3032 5778 3088
rect 8956 8186 9012 8188
rect 9036 8186 9092 8188
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 8956 8134 8982 8186
rect 8982 8134 9012 8186
rect 9036 8134 9046 8186
rect 9046 8134 9092 8186
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9252 8186
rect 8956 8132 9012 8134
rect 9036 8132 9092 8134
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 4956 2202 5012 2204
rect 5036 2202 5092 2204
rect 5116 2202 5172 2204
rect 5196 2202 5252 2204
rect 4956 2150 4982 2202
rect 4982 2150 5012 2202
rect 5036 2150 5046 2202
rect 5046 2150 5092 2202
rect 5116 2150 5162 2202
rect 5162 2150 5172 2202
rect 5196 2150 5226 2202
rect 5226 2150 5252 2202
rect 4956 2148 5012 2150
rect 5036 2148 5092 2150
rect 5116 2148 5172 2150
rect 5196 2148 5252 2150
rect 8956 7098 9012 7100
rect 9036 7098 9092 7100
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 8956 7046 8982 7098
rect 8982 7046 9012 7098
rect 9036 7046 9046 7098
rect 9046 7046 9092 7098
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9252 7098
rect 8956 7044 9012 7046
rect 9036 7044 9092 7046
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 8956 6010 9012 6012
rect 9036 6010 9092 6012
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 8956 5958 8982 6010
rect 8982 5958 9012 6010
rect 9036 5958 9046 6010
rect 9046 5958 9092 6010
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9252 6010
rect 8956 5956 9012 5958
rect 9036 5956 9092 5958
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 10782 11600 10838 11656
rect 12956 21786 13012 21788
rect 13036 21786 13092 21788
rect 13116 21786 13172 21788
rect 13196 21786 13252 21788
rect 12956 21734 12982 21786
rect 12982 21734 13012 21786
rect 13036 21734 13046 21786
rect 13046 21734 13092 21786
rect 13116 21734 13162 21786
rect 13162 21734 13172 21786
rect 13196 21734 13226 21786
rect 13226 21734 13252 21786
rect 12956 21732 13012 21734
rect 13036 21732 13092 21734
rect 13116 21732 13172 21734
rect 13196 21732 13252 21734
rect 12956 20698 13012 20700
rect 13036 20698 13092 20700
rect 13116 20698 13172 20700
rect 13196 20698 13252 20700
rect 12956 20646 12982 20698
rect 12982 20646 13012 20698
rect 13036 20646 13046 20698
rect 13046 20646 13092 20698
rect 13116 20646 13162 20698
rect 13162 20646 13172 20698
rect 13196 20646 13226 20698
rect 13226 20646 13252 20698
rect 12956 20644 13012 20646
rect 13036 20644 13092 20646
rect 13116 20644 13172 20646
rect 13196 20644 13252 20646
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 16982 21242
rect 16982 21190 17012 21242
rect 17036 21190 17046 21242
rect 17046 21190 17092 21242
rect 17116 21190 17162 21242
rect 17162 21190 17172 21242
rect 17196 21190 17226 21242
rect 17226 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 12956 19610 13012 19612
rect 13036 19610 13092 19612
rect 13116 19610 13172 19612
rect 13196 19610 13252 19612
rect 12956 19558 12982 19610
rect 12982 19558 13012 19610
rect 13036 19558 13046 19610
rect 13046 19558 13092 19610
rect 13116 19558 13162 19610
rect 13162 19558 13172 19610
rect 13196 19558 13226 19610
rect 13226 19558 13252 19610
rect 12956 19556 13012 19558
rect 13036 19556 13092 19558
rect 13116 19556 13172 19558
rect 13196 19556 13252 19558
rect 12956 18522 13012 18524
rect 13036 18522 13092 18524
rect 13116 18522 13172 18524
rect 13196 18522 13252 18524
rect 12956 18470 12982 18522
rect 12982 18470 13012 18522
rect 13036 18470 13046 18522
rect 13046 18470 13092 18522
rect 13116 18470 13162 18522
rect 13162 18470 13172 18522
rect 13196 18470 13226 18522
rect 13226 18470 13252 18522
rect 12956 18468 13012 18470
rect 13036 18468 13092 18470
rect 13116 18468 13172 18470
rect 13196 18468 13252 18470
rect 12956 17434 13012 17436
rect 13036 17434 13092 17436
rect 13116 17434 13172 17436
rect 13196 17434 13252 17436
rect 12956 17382 12982 17434
rect 12982 17382 13012 17434
rect 13036 17382 13046 17434
rect 13046 17382 13092 17434
rect 13116 17382 13162 17434
rect 13162 17382 13172 17434
rect 13196 17382 13226 17434
rect 13226 17382 13252 17434
rect 12956 17380 13012 17382
rect 13036 17380 13092 17382
rect 13116 17380 13172 17382
rect 13196 17380 13252 17382
rect 12956 16346 13012 16348
rect 13036 16346 13092 16348
rect 13116 16346 13172 16348
rect 13196 16346 13252 16348
rect 12956 16294 12982 16346
rect 12982 16294 13012 16346
rect 13036 16294 13046 16346
rect 13046 16294 13092 16346
rect 13116 16294 13162 16346
rect 13162 16294 13172 16346
rect 13196 16294 13226 16346
rect 13226 16294 13252 16346
rect 12956 16292 13012 16294
rect 13036 16292 13092 16294
rect 13116 16292 13172 16294
rect 13196 16292 13252 16294
rect 12956 15258 13012 15260
rect 13036 15258 13092 15260
rect 13116 15258 13172 15260
rect 13196 15258 13252 15260
rect 12956 15206 12982 15258
rect 12982 15206 13012 15258
rect 13036 15206 13046 15258
rect 13046 15206 13092 15258
rect 13116 15206 13162 15258
rect 13162 15206 13172 15258
rect 13196 15206 13226 15258
rect 13226 15206 13252 15258
rect 12956 15204 13012 15206
rect 13036 15204 13092 15206
rect 13116 15204 13172 15206
rect 13196 15204 13252 15206
rect 12956 14170 13012 14172
rect 13036 14170 13092 14172
rect 13116 14170 13172 14172
rect 13196 14170 13252 14172
rect 12956 14118 12982 14170
rect 12982 14118 13012 14170
rect 13036 14118 13046 14170
rect 13046 14118 13092 14170
rect 13116 14118 13162 14170
rect 13162 14118 13172 14170
rect 13196 14118 13226 14170
rect 13226 14118 13252 14170
rect 12956 14116 13012 14118
rect 13036 14116 13092 14118
rect 13116 14116 13172 14118
rect 13196 14116 13252 14118
rect 12956 13082 13012 13084
rect 13036 13082 13092 13084
rect 13116 13082 13172 13084
rect 13196 13082 13252 13084
rect 12956 13030 12982 13082
rect 12982 13030 13012 13082
rect 13036 13030 13046 13082
rect 13046 13030 13092 13082
rect 13116 13030 13162 13082
rect 13162 13030 13172 13082
rect 13196 13030 13226 13082
rect 13226 13030 13252 13082
rect 12956 13028 13012 13030
rect 13036 13028 13092 13030
rect 13116 13028 13172 13030
rect 13196 13028 13252 13030
rect 12956 11994 13012 11996
rect 13036 11994 13092 11996
rect 13116 11994 13172 11996
rect 13196 11994 13252 11996
rect 12956 11942 12982 11994
rect 12982 11942 13012 11994
rect 13036 11942 13046 11994
rect 13046 11942 13092 11994
rect 13116 11942 13162 11994
rect 13162 11942 13172 11994
rect 13196 11942 13226 11994
rect 13226 11942 13252 11994
rect 12956 11940 13012 11942
rect 13036 11940 13092 11942
rect 13116 11940 13172 11942
rect 13196 11940 13252 11942
rect 7654 1264 7710 1320
rect 8956 4922 9012 4924
rect 9036 4922 9092 4924
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 8956 4870 8982 4922
rect 8982 4870 9012 4922
rect 9036 4870 9046 4922
rect 9046 4870 9092 4922
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9252 4922
rect 8956 4868 9012 4870
rect 9036 4868 9092 4870
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 8956 3834 9012 3836
rect 9036 3834 9092 3836
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 8956 3782 8982 3834
rect 8982 3782 9012 3834
rect 9036 3782 9046 3834
rect 9046 3782 9092 3834
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9252 3834
rect 8956 3780 9012 3782
rect 9036 3780 9092 3782
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 12956 10906 13012 10908
rect 13036 10906 13092 10908
rect 13116 10906 13172 10908
rect 13196 10906 13252 10908
rect 12956 10854 12982 10906
rect 12982 10854 13012 10906
rect 13036 10854 13046 10906
rect 13046 10854 13092 10906
rect 13116 10854 13162 10906
rect 13162 10854 13172 10906
rect 13196 10854 13226 10906
rect 13226 10854 13252 10906
rect 12956 10852 13012 10854
rect 13036 10852 13092 10854
rect 13116 10852 13172 10854
rect 13196 10852 13252 10854
rect 12956 9818 13012 9820
rect 13036 9818 13092 9820
rect 13116 9818 13172 9820
rect 13196 9818 13252 9820
rect 12956 9766 12982 9818
rect 12982 9766 13012 9818
rect 13036 9766 13046 9818
rect 13046 9766 13092 9818
rect 13116 9766 13162 9818
rect 13162 9766 13172 9818
rect 13196 9766 13226 9818
rect 13226 9766 13252 9818
rect 12956 9764 13012 9766
rect 13036 9764 13092 9766
rect 13116 9764 13172 9766
rect 13196 9764 13252 9766
rect 12956 8730 13012 8732
rect 13036 8730 13092 8732
rect 13116 8730 13172 8732
rect 13196 8730 13252 8732
rect 12956 8678 12982 8730
rect 12982 8678 13012 8730
rect 13036 8678 13046 8730
rect 13046 8678 13092 8730
rect 13116 8678 13162 8730
rect 13162 8678 13172 8730
rect 13196 8678 13226 8730
rect 13226 8678 13252 8730
rect 12956 8676 13012 8678
rect 13036 8676 13092 8678
rect 13116 8676 13172 8678
rect 13196 8676 13252 8678
rect 11242 6160 11298 6216
rect 12956 7642 13012 7644
rect 13036 7642 13092 7644
rect 13116 7642 13172 7644
rect 13196 7642 13252 7644
rect 12956 7590 12982 7642
rect 12982 7590 13012 7642
rect 13036 7590 13046 7642
rect 13046 7590 13092 7642
rect 13116 7590 13162 7642
rect 13162 7590 13172 7642
rect 13196 7590 13226 7642
rect 13226 7590 13252 7642
rect 12956 7588 13012 7590
rect 13036 7588 13092 7590
rect 13116 7588 13172 7590
rect 13196 7588 13252 7590
rect 9770 2896 9826 2952
rect 8956 2746 9012 2748
rect 9036 2746 9092 2748
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 8956 2694 8982 2746
rect 8982 2694 9012 2746
rect 9036 2694 9046 2746
rect 9046 2694 9092 2746
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9252 2746
rect 8956 2692 9012 2694
rect 9036 2692 9092 2694
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 12956 6554 13012 6556
rect 13036 6554 13092 6556
rect 13116 6554 13172 6556
rect 13196 6554 13252 6556
rect 12956 6502 12982 6554
rect 12982 6502 13012 6554
rect 13036 6502 13046 6554
rect 13046 6502 13092 6554
rect 13116 6502 13162 6554
rect 13162 6502 13172 6554
rect 13196 6502 13226 6554
rect 13226 6502 13252 6554
rect 12956 6500 13012 6502
rect 13036 6500 13092 6502
rect 13116 6500 13172 6502
rect 13196 6500 13252 6502
rect 12956 5466 13012 5468
rect 13036 5466 13092 5468
rect 13116 5466 13172 5468
rect 13196 5466 13252 5468
rect 12956 5414 12982 5466
rect 12982 5414 13012 5466
rect 13036 5414 13046 5466
rect 13046 5414 13092 5466
rect 13116 5414 13162 5466
rect 13162 5414 13172 5466
rect 13196 5414 13226 5466
rect 13226 5414 13252 5466
rect 12956 5412 13012 5414
rect 13036 5412 13092 5414
rect 13116 5412 13172 5414
rect 13196 5412 13252 5414
rect 12956 4378 13012 4380
rect 13036 4378 13092 4380
rect 13116 4378 13172 4380
rect 13196 4378 13252 4380
rect 12956 4326 12982 4378
rect 12982 4326 13012 4378
rect 13036 4326 13046 4378
rect 13046 4326 13092 4378
rect 13116 4326 13162 4378
rect 13162 4326 13172 4378
rect 13196 4326 13226 4378
rect 13226 4326 13252 4378
rect 12956 4324 13012 4326
rect 13036 4324 13092 4326
rect 13116 4324 13172 4326
rect 13196 4324 13252 4326
rect 12956 3290 13012 3292
rect 13036 3290 13092 3292
rect 13116 3290 13172 3292
rect 13196 3290 13252 3292
rect 12956 3238 12982 3290
rect 12982 3238 13012 3290
rect 13036 3238 13046 3290
rect 13046 3238 13092 3290
rect 13116 3238 13162 3290
rect 13162 3238 13172 3290
rect 13196 3238 13226 3290
rect 13226 3238 13252 3290
rect 12956 3236 13012 3238
rect 13036 3236 13092 3238
rect 13116 3236 13172 3238
rect 13196 3236 13252 3238
rect 12956 2202 13012 2204
rect 13036 2202 13092 2204
rect 13116 2202 13172 2204
rect 13196 2202 13252 2204
rect 12956 2150 12982 2202
rect 12982 2150 13012 2202
rect 13036 2150 13046 2202
rect 13046 2150 13092 2202
rect 13116 2150 13162 2202
rect 13162 2150 13172 2202
rect 13196 2150 13226 2202
rect 13226 2150 13252 2202
rect 12956 2148 13012 2150
rect 13036 2148 13092 2150
rect 13116 2148 13172 2150
rect 13196 2148 13252 2150
rect 12806 1128 12862 1184
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 16982 20154
rect 16982 20102 17012 20154
rect 17036 20102 17046 20154
rect 17046 20102 17092 20154
rect 17116 20102 17162 20154
rect 17162 20102 17172 20154
rect 17196 20102 17226 20154
rect 17226 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 16982 19066
rect 16982 19014 17012 19066
rect 17036 19014 17046 19066
rect 17046 19014 17092 19066
rect 17116 19014 17162 19066
rect 17162 19014 17172 19066
rect 17196 19014 17226 19066
rect 17226 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 15382 17584 15438 17640
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 16982 17978
rect 16982 17926 17012 17978
rect 17036 17926 17046 17978
rect 17046 17926 17092 17978
rect 17116 17926 17162 17978
rect 17162 17926 17172 17978
rect 17196 17926 17226 17978
rect 17226 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 16394 17040 16450 17096
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 16982 16890
rect 16982 16838 17012 16890
rect 17036 16838 17046 16890
rect 17046 16838 17092 16890
rect 17116 16838 17162 16890
rect 17162 16838 17172 16890
rect 17196 16838 17226 16890
rect 17226 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 16982 15802
rect 16982 15750 17012 15802
rect 17036 15750 17046 15802
rect 17046 15750 17092 15802
rect 17116 15750 17162 15802
rect 17162 15750 17172 15802
rect 17196 15750 17226 15802
rect 17226 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16670 15000 16726 15056
rect 14922 14864 14978 14920
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 16982 14714
rect 16982 14662 17012 14714
rect 17036 14662 17046 14714
rect 17046 14662 17092 14714
rect 17116 14662 17162 14714
rect 17162 14662 17172 14714
rect 17196 14662 17226 14714
rect 17226 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 16982 13626
rect 16982 13574 17012 13626
rect 17036 13574 17046 13626
rect 17046 13574 17092 13626
rect 17116 13574 17162 13626
rect 17162 13574 17172 13626
rect 17196 13574 17226 13626
rect 17226 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 16982 12538
rect 16982 12486 17012 12538
rect 17036 12486 17046 12538
rect 17046 12486 17092 12538
rect 17116 12486 17162 12538
rect 17162 12486 17172 12538
rect 17196 12486 17226 12538
rect 17226 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 16982 11450
rect 16982 11398 17012 11450
rect 17036 11398 17046 11450
rect 17046 11398 17092 11450
rect 17116 11398 17162 11450
rect 17162 11398 17172 11450
rect 17196 11398 17226 11450
rect 17226 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 16982 10362
rect 16982 10310 17012 10362
rect 17036 10310 17046 10362
rect 17046 10310 17092 10362
rect 17116 10310 17162 10362
rect 17162 10310 17172 10362
rect 17196 10310 17226 10362
rect 17226 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 16982 9274
rect 16982 9222 17012 9274
rect 17036 9222 17046 9274
rect 17046 9222 17092 9274
rect 17116 9222 17162 9274
rect 17162 9222 17172 9274
rect 17196 9222 17226 9274
rect 17226 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 16982 8186
rect 16982 8134 17012 8186
rect 17036 8134 17046 8186
rect 17046 8134 17092 8186
rect 17116 8134 17162 8186
rect 17162 8134 17172 8186
rect 17196 8134 17226 8186
rect 17226 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 16982 7098
rect 16982 7046 17012 7098
rect 17036 7046 17046 7098
rect 17046 7046 17092 7098
rect 17116 7046 17162 7098
rect 17162 7046 17172 7098
rect 17196 7046 17226 7098
rect 17226 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 17314 6160 17370 6216
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 16982 6010
rect 16982 5958 17012 6010
rect 17036 5958 17046 6010
rect 17046 5958 17092 6010
rect 17116 5958 17162 6010
rect 17162 5958 17172 6010
rect 17196 5958 17226 6010
rect 17226 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 16982 4922
rect 16982 4870 17012 4922
rect 17036 4870 17046 4922
rect 17046 4870 17092 4922
rect 17116 4870 17162 4922
rect 17162 4870 17172 4922
rect 17196 4870 17226 4922
rect 17226 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 16982 3834
rect 16982 3782 17012 3834
rect 17036 3782 17046 3834
rect 17046 3782 17092 3834
rect 17116 3782 17162 3834
rect 17162 3782 17172 3834
rect 17196 3782 17226 3834
rect 17226 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 16982 2746
rect 16982 2694 17012 2746
rect 17036 2694 17046 2746
rect 17046 2694 17092 2746
rect 17116 2694 17162 2746
rect 17162 2694 17172 2746
rect 17196 2694 17226 2746
rect 17226 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 14646 1672 14702 1728
rect 16946 1264 17002 1320
rect 20956 21786 21012 21788
rect 21036 21786 21092 21788
rect 21116 21786 21172 21788
rect 21196 21786 21252 21788
rect 20956 21734 20982 21786
rect 20982 21734 21012 21786
rect 21036 21734 21046 21786
rect 21046 21734 21092 21786
rect 21116 21734 21162 21786
rect 21162 21734 21172 21786
rect 21196 21734 21226 21786
rect 21226 21734 21252 21786
rect 20956 21732 21012 21734
rect 21036 21732 21092 21734
rect 21116 21732 21172 21734
rect 21196 21732 21252 21734
rect 20956 20698 21012 20700
rect 21036 20698 21092 20700
rect 21116 20698 21172 20700
rect 21196 20698 21252 20700
rect 20956 20646 20982 20698
rect 20982 20646 21012 20698
rect 21036 20646 21046 20698
rect 21046 20646 21092 20698
rect 21116 20646 21162 20698
rect 21162 20646 21172 20698
rect 21196 20646 21226 20698
rect 21226 20646 21252 20698
rect 20956 20644 21012 20646
rect 21036 20644 21092 20646
rect 21116 20644 21172 20646
rect 21196 20644 21252 20646
rect 21454 22072 21510 22128
rect 19890 14864 19946 14920
rect 21270 19760 21326 19816
rect 20956 19610 21012 19612
rect 21036 19610 21092 19612
rect 21116 19610 21172 19612
rect 21196 19610 21252 19612
rect 20956 19558 20982 19610
rect 20982 19558 21012 19610
rect 21036 19558 21046 19610
rect 21046 19558 21092 19610
rect 21116 19558 21162 19610
rect 21162 19558 21172 19610
rect 21196 19558 21226 19610
rect 21226 19558 21252 19610
rect 20956 19556 21012 19558
rect 21036 19556 21092 19558
rect 21116 19556 21172 19558
rect 21196 19556 21252 19558
rect 20956 18522 21012 18524
rect 21036 18522 21092 18524
rect 21116 18522 21172 18524
rect 21196 18522 21252 18524
rect 20956 18470 20982 18522
rect 20982 18470 21012 18522
rect 21036 18470 21046 18522
rect 21046 18470 21092 18522
rect 21116 18470 21162 18522
rect 21162 18470 21172 18522
rect 21196 18470 21226 18522
rect 21226 18470 21252 18522
rect 20956 18468 21012 18470
rect 21036 18468 21092 18470
rect 21116 18468 21172 18470
rect 21196 18468 21252 18470
rect 20956 17434 21012 17436
rect 21036 17434 21092 17436
rect 21116 17434 21172 17436
rect 21196 17434 21252 17436
rect 20956 17382 20982 17434
rect 20982 17382 21012 17434
rect 21036 17382 21046 17434
rect 21046 17382 21092 17434
rect 21116 17382 21162 17434
rect 21162 17382 21172 17434
rect 21196 17382 21226 17434
rect 21226 17382 21252 17434
rect 20956 17380 21012 17382
rect 21036 17380 21092 17382
rect 21116 17380 21172 17382
rect 21196 17380 21252 17382
rect 20956 16346 21012 16348
rect 21036 16346 21092 16348
rect 21116 16346 21172 16348
rect 21196 16346 21252 16348
rect 20956 16294 20982 16346
rect 20982 16294 21012 16346
rect 21036 16294 21046 16346
rect 21046 16294 21092 16346
rect 21116 16294 21162 16346
rect 21162 16294 21172 16346
rect 21196 16294 21226 16346
rect 21226 16294 21252 16346
rect 20956 16292 21012 16294
rect 21036 16292 21092 16294
rect 21116 16292 21172 16294
rect 21196 16292 21252 16294
rect 20956 15258 21012 15260
rect 21036 15258 21092 15260
rect 21116 15258 21172 15260
rect 21196 15258 21252 15260
rect 20956 15206 20982 15258
rect 20982 15206 21012 15258
rect 21036 15206 21046 15258
rect 21046 15206 21092 15258
rect 21116 15206 21162 15258
rect 21162 15206 21172 15258
rect 21196 15206 21226 15258
rect 21226 15206 21252 15258
rect 20956 15204 21012 15206
rect 21036 15204 21092 15206
rect 21116 15204 21172 15206
rect 21196 15204 21252 15206
rect 20956 14170 21012 14172
rect 21036 14170 21092 14172
rect 21116 14170 21172 14172
rect 21196 14170 21252 14172
rect 20956 14118 20982 14170
rect 20982 14118 21012 14170
rect 21036 14118 21046 14170
rect 21046 14118 21092 14170
rect 21116 14118 21162 14170
rect 21162 14118 21172 14170
rect 21196 14118 21226 14170
rect 21226 14118 21252 14170
rect 20956 14116 21012 14118
rect 21036 14116 21092 14118
rect 21116 14116 21172 14118
rect 21196 14116 21252 14118
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 21086 12552 21142 12608
rect 20626 12144 20682 12200
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 23570 10648 23626 10704
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 17682 6296 17738 6352
rect 21454 7656 21510 7712
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 23294 1128 23350 1184
<< metal3 >>
rect 0 23352 480 23384
rect 0 23296 110 23352
rect 166 23296 480 23352
rect 0 23264 480 23296
rect 23520 22584 24000 22704
rect 0 22176 480 22296
rect 62 21722 122 22176
rect 21449 22130 21515 22133
rect 23614 22130 23674 22584
rect 21449 22128 23674 22130
rect 21449 22072 21454 22128
rect 21510 22072 23674 22128
rect 21449 22070 23674 22072
rect 21449 22067 21515 22070
rect 4944 21792 5264 21793
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 21727 5264 21728
rect 12944 21792 13264 21793
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 21727 13264 21728
rect 20944 21792 21264 21793
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 21727 21264 21728
rect 1209 21722 1275 21725
rect 62 21720 1275 21722
rect 62 21664 1214 21720
rect 1270 21664 1275 21720
rect 62 21662 1275 21664
rect 1209 21659 1275 21662
rect 8944 21248 9264 21249
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 21183 9264 21184
rect 16944 21248 17264 21249
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 21183 17264 21184
rect 0 20952 480 21072
rect 62 20498 122 20952
rect 4944 20704 5264 20705
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 20639 5264 20640
rect 12944 20704 13264 20705
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 20639 13264 20640
rect 20944 20704 21264 20705
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 20639 21264 20640
rect 1577 20498 1643 20501
rect 62 20496 1643 20498
rect 62 20440 1582 20496
rect 1638 20440 1643 20496
rect 62 20438 1643 20440
rect 1577 20435 1643 20438
rect 8944 20160 9264 20161
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 20095 9264 20096
rect 16944 20160 17264 20161
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 23520 20136 24000 20256
rect 16944 20095 17264 20096
rect 0 19864 480 19984
rect 62 19546 122 19864
rect 21265 19818 21331 19821
rect 23614 19818 23674 20136
rect 21265 19816 23674 19818
rect 21265 19760 21270 19816
rect 21326 19760 23674 19816
rect 21265 19758 23674 19760
rect 21265 19755 21331 19758
rect 4944 19616 5264 19617
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 19551 5264 19552
rect 12944 19616 13264 19617
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 19551 13264 19552
rect 20944 19616 21264 19617
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 19551 21264 19552
rect 1577 19546 1643 19549
rect 62 19544 1643 19546
rect 62 19488 1582 19544
rect 1638 19488 1643 19544
rect 62 19486 1643 19488
rect 1577 19483 1643 19486
rect 8944 19072 9264 19073
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 19007 9264 19008
rect 16944 19072 17264 19073
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 19007 17264 19008
rect 0 18864 480 18896
rect 0 18808 110 18864
rect 166 18808 480 18864
rect 0 18776 480 18808
rect 4944 18528 5264 18529
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 18463 5264 18464
rect 12944 18528 13264 18529
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 18463 13264 18464
rect 20944 18528 21264 18529
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 18463 21264 18464
rect 8944 17984 9264 17985
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 17919 9264 17920
rect 16944 17984 17264 17985
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 17919 17264 17920
rect 23520 17824 24000 17944
rect 0 17552 480 17672
rect 15377 17642 15443 17645
rect 23614 17642 23674 17824
rect 15377 17640 23674 17642
rect 15377 17584 15382 17640
rect 15438 17584 23674 17640
rect 15377 17582 23674 17584
rect 15377 17579 15443 17582
rect 62 17098 122 17552
rect 4944 17440 5264 17441
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 17375 5264 17376
rect 12944 17440 13264 17441
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 17375 13264 17376
rect 20944 17440 21264 17441
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 17375 21264 17376
rect 1577 17098 1643 17101
rect 62 17096 1643 17098
rect 62 17040 1582 17096
rect 1638 17040 1643 17096
rect 62 17038 1643 17040
rect 1577 17035 1643 17038
rect 10225 17098 10291 17101
rect 16389 17098 16455 17101
rect 10225 17096 16455 17098
rect 10225 17040 10230 17096
rect 10286 17040 16394 17096
rect 16450 17040 16455 17096
rect 10225 17038 16455 17040
rect 10225 17035 10291 17038
rect 16389 17035 16455 17038
rect 8944 16896 9264 16897
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 16831 9264 16832
rect 16944 16896 17264 16897
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 16831 17264 16832
rect 0 16464 480 16584
rect 62 16010 122 16464
rect 4944 16352 5264 16353
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 16287 5264 16288
rect 12944 16352 13264 16353
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 16287 13264 16288
rect 20944 16352 21264 16353
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 16287 21264 16288
rect 5717 16010 5783 16013
rect 62 16008 5783 16010
rect 62 15952 5722 16008
rect 5778 15952 5783 16008
rect 62 15950 5783 15952
rect 5717 15947 5783 15950
rect 8944 15808 9264 15809
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 15743 9264 15744
rect 16944 15808 17264 15809
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 15743 17264 15744
rect 23520 15376 24000 15496
rect 0 15240 480 15360
rect 4944 15264 5264 15265
rect 62 15058 122 15240
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 15199 5264 15200
rect 12944 15264 13264 15265
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 15199 13264 15200
rect 20944 15264 21264 15265
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 15199 21264 15200
rect 5993 15058 6059 15061
rect 62 15056 6059 15058
rect 62 15000 5998 15056
rect 6054 15000 6059 15056
rect 62 14998 6059 15000
rect 5993 14995 6059 14998
rect 6269 15058 6335 15061
rect 16665 15058 16731 15061
rect 6269 15056 16731 15058
rect 6269 15000 6274 15056
rect 6330 15000 16670 15056
rect 16726 15000 16731 15056
rect 6269 14998 16731 15000
rect 6269 14995 6335 14998
rect 16665 14995 16731 14998
rect 4061 14922 4127 14925
rect 14917 14922 14983 14925
rect 4061 14920 14983 14922
rect 4061 14864 4066 14920
rect 4122 14864 14922 14920
rect 14978 14864 14983 14920
rect 4061 14862 14983 14864
rect 4061 14859 4127 14862
rect 14917 14859 14983 14862
rect 19885 14922 19951 14925
rect 23614 14922 23674 15376
rect 19885 14920 23674 14922
rect 19885 14864 19890 14920
rect 19946 14864 23674 14920
rect 19885 14862 23674 14864
rect 19885 14859 19951 14862
rect 2129 14786 2195 14789
rect 62 14784 2195 14786
rect 62 14728 2134 14784
rect 2190 14728 2195 14784
rect 62 14726 2195 14728
rect 62 14272 122 14726
rect 2129 14723 2195 14726
rect 8944 14720 9264 14721
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 14655 9264 14656
rect 16944 14720 17264 14721
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 14655 17264 14656
rect 0 14152 480 14272
rect 4944 14176 5264 14177
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 14111 5264 14112
rect 12944 14176 13264 14177
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 14111 13264 14112
rect 20944 14176 21264 14177
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 14111 21264 14112
rect 8944 13632 9264 13633
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 13567 9264 13568
rect 16944 13632 17264 13633
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13567 17264 13568
rect 0 13064 480 13184
rect 4944 13088 5264 13089
rect 62 12610 122 13064
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 13023 5264 13024
rect 12944 13088 13264 13089
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 13023 13264 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 23520 13064 24000 13184
rect 20944 13023 21264 13024
rect 1485 12610 1551 12613
rect 62 12608 1551 12610
rect 62 12552 1490 12608
rect 1546 12552 1551 12608
rect 62 12550 1551 12552
rect 1485 12547 1551 12550
rect 21081 12610 21147 12613
rect 23614 12610 23674 13064
rect 21081 12608 23674 12610
rect 21081 12552 21086 12608
rect 21142 12552 23674 12608
rect 21081 12550 23674 12552
rect 21081 12547 21147 12550
rect 8944 12544 9264 12545
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 12479 9264 12480
rect 16944 12544 17264 12545
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 12479 17264 12480
rect 9121 12202 9187 12205
rect 20621 12202 20687 12205
rect 9121 12200 20687 12202
rect 9121 12144 9126 12200
rect 9182 12144 20626 12200
rect 20682 12144 20687 12200
rect 9121 12142 20687 12144
rect 9121 12139 9187 12142
rect 20621 12139 20687 12142
rect 4944 12000 5264 12001
rect 0 11928 480 11960
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 11935 5264 11936
rect 12944 12000 13264 12001
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 11935 13264 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 0 11872 110 11928
rect 166 11872 480 11928
rect 0 11840 480 11872
rect 3969 11658 4035 11661
rect 10777 11658 10843 11661
rect 3969 11656 10843 11658
rect 3969 11600 3974 11656
rect 4030 11600 10782 11656
rect 10838 11600 10843 11656
rect 3969 11598 10843 11600
rect 3969 11595 4035 11598
rect 10777 11595 10843 11598
rect 8944 11456 9264 11457
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 11391 9264 11392
rect 16944 11456 17264 11457
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 11391 17264 11392
rect 4944 10912 5264 10913
rect 0 10840 480 10872
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 10847 5264 10848
rect 12944 10912 13264 10913
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 10847 13264 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 0 10784 110 10840
rect 166 10784 480 10840
rect 0 10752 480 10784
rect 23520 10706 24000 10736
rect 23484 10704 24000 10706
rect 23484 10648 23570 10704
rect 23626 10648 24000 10704
rect 23484 10646 24000 10648
rect 23520 10616 24000 10646
rect 8944 10368 9264 10369
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 10303 9264 10304
rect 16944 10368 17264 10369
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 10303 17264 10304
rect 4944 9824 5264 9825
rect 0 9752 480 9784
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 9759 5264 9760
rect 12944 9824 13264 9825
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 9759 13264 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 0 9696 110 9752
rect 166 9696 480 9752
rect 0 9664 480 9696
rect 8944 9280 9264 9281
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 9215 9264 9216
rect 16944 9280 17264 9281
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 9215 17264 9216
rect 4944 8736 5264 8737
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 8671 5264 8672
rect 12944 8736 13264 8737
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 8671 13264 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 0 8440 480 8560
rect 62 7986 122 8440
rect 8944 8192 9264 8193
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 8127 9264 8128
rect 16944 8192 17264 8193
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 23520 8168 24000 8288
rect 16944 8127 17264 8128
rect 6729 7986 6795 7989
rect 62 7984 6795 7986
rect 62 7928 6734 7984
rect 6790 7928 6795 7984
rect 62 7926 6795 7928
rect 6729 7923 6795 7926
rect 21449 7714 21515 7717
rect 23614 7714 23674 8168
rect 21449 7712 23674 7714
rect 21449 7656 21454 7712
rect 21510 7656 23674 7712
rect 21449 7654 23674 7656
rect 21449 7651 21515 7654
rect 4944 7648 5264 7649
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 7583 5264 7584
rect 12944 7648 13264 7649
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 7583 13264 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 0 7440 480 7472
rect 0 7384 110 7440
rect 166 7384 480 7440
rect 0 7352 480 7384
rect 4153 7170 4219 7173
rect 5625 7170 5691 7173
rect 4153 7168 5691 7170
rect 4153 7112 4158 7168
rect 4214 7112 5630 7168
rect 5686 7112 5691 7168
rect 4153 7110 5691 7112
rect 4153 7107 4219 7110
rect 5625 7107 5691 7110
rect 8944 7104 9264 7105
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 7039 9264 7040
rect 16944 7104 17264 7105
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 7039 17264 7040
rect 4944 6560 5264 6561
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 6495 5264 6496
rect 12944 6560 13264 6561
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 6495 13264 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 17677 6354 17743 6357
rect 17677 6352 23674 6354
rect 17677 6296 17682 6352
rect 17738 6296 23674 6352
rect 17677 6294 23674 6296
rect 17677 6291 17743 6294
rect 0 6128 480 6248
rect 11237 6218 11303 6221
rect 17309 6218 17375 6221
rect 11237 6216 17375 6218
rect 11237 6160 11242 6216
rect 11298 6160 17314 6216
rect 17370 6160 17375 6216
rect 11237 6158 17375 6160
rect 11237 6155 11303 6158
rect 17309 6155 17375 6158
rect 62 5674 122 6128
rect 8944 6016 9264 6017
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 5951 9264 5952
rect 16944 6016 17264 6017
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 23614 5976 23674 6294
rect 16944 5951 17264 5952
rect 23520 5856 24000 5976
rect 4797 5674 4863 5677
rect 62 5672 4863 5674
rect 62 5616 4802 5672
rect 4858 5616 4863 5672
rect 62 5614 4863 5616
rect 4797 5611 4863 5614
rect 4944 5472 5264 5473
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 5407 5264 5408
rect 12944 5472 13264 5473
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 5407 13264 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 4981 5266 5047 5269
rect 5625 5266 5691 5269
rect 4981 5264 5691 5266
rect 4981 5208 4986 5264
rect 5042 5208 5630 5264
rect 5686 5208 5691 5264
rect 4981 5206 5691 5208
rect 4981 5203 5047 5206
rect 5625 5203 5691 5206
rect 0 5040 480 5160
rect 3601 5130 3667 5133
rect 4613 5130 4679 5133
rect 3601 5128 4679 5130
rect 3601 5072 3606 5128
rect 3662 5072 4618 5128
rect 4674 5072 4679 5128
rect 3601 5070 4679 5072
rect 3601 5067 3667 5070
rect 4613 5067 4679 5070
rect 62 4586 122 5040
rect 8944 4928 9264 4929
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 4863 9264 4864
rect 16944 4928 17264 4929
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 4863 17264 4864
rect 1577 4586 1643 4589
rect 62 4584 1643 4586
rect 62 4528 1582 4584
rect 1638 4528 1643 4584
rect 62 4526 1643 4528
rect 1577 4523 1643 4526
rect 4944 4384 5264 4385
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 4319 5264 4320
rect 12944 4384 13264 4385
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 4319 13264 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 0 3952 480 4072
rect 62 3498 122 3952
rect 8944 3840 9264 3841
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 3775 9264 3776
rect 16944 3840 17264 3841
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3775 17264 3776
rect 1209 3498 1275 3501
rect 62 3496 1275 3498
rect 62 3440 1214 3496
rect 1270 3440 1275 3496
rect 62 3438 1275 3440
rect 1209 3435 1275 3438
rect 23520 3408 24000 3528
rect 4944 3296 5264 3297
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 3231 5264 3232
rect 12944 3296 13264 3297
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 3231 13264 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 5717 3090 5783 3093
rect 62 3088 5783 3090
rect 62 3032 5722 3088
rect 5778 3032 5783 3088
rect 62 3030 5783 3032
rect 62 2848 122 3030
rect 5717 3027 5783 3030
rect 9765 2954 9831 2957
rect 23614 2954 23674 3408
rect 9765 2952 23674 2954
rect 9765 2896 9770 2952
rect 9826 2896 23674 2952
rect 9765 2894 23674 2896
rect 9765 2891 9831 2894
rect 0 2728 480 2848
rect 8944 2752 9264 2753
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2687 9264 2688
rect 16944 2752 17264 2753
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2687 17264 2688
rect 4944 2208 5264 2209
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2143 5264 2144
rect 12944 2208 13264 2209
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2143 13264 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 1853 2002 1919 2005
rect 62 2000 1919 2002
rect 62 1944 1858 2000
rect 1914 1944 1919 2000
rect 62 1942 1919 1944
rect 62 1760 122 1942
rect 1853 1939 1919 1942
rect 0 1640 480 1760
rect 14641 1730 14707 1733
rect 14641 1728 23674 1730
rect 14641 1672 14646 1728
rect 14702 1672 23674 1728
rect 14641 1670 23674 1672
rect 14641 1667 14707 1670
rect 7649 1322 7715 1325
rect 16941 1322 17007 1325
rect 7649 1320 17007 1322
rect 7649 1264 7654 1320
rect 7710 1264 16946 1320
rect 17002 1264 17007 1320
rect 7649 1262 17007 1264
rect 7649 1259 7715 1262
rect 16941 1259 17007 1262
rect 23614 1216 23674 1670
rect 2129 1186 2195 1189
rect 62 1184 2195 1186
rect 62 1128 2134 1184
rect 2190 1128 2195 1184
rect 62 1126 2195 1128
rect 62 672 122 1126
rect 2129 1123 2195 1126
rect 12801 1186 12867 1189
rect 23289 1186 23355 1189
rect 12801 1184 23355 1186
rect 12801 1128 12806 1184
rect 12862 1128 23294 1184
rect 23350 1128 23355 1184
rect 12801 1126 23355 1128
rect 12801 1123 12867 1126
rect 23289 1123 23355 1126
rect 23520 1096 24000 1216
rect 0 552 480 672
<< via3 >>
rect 4952 21788 5016 21792
rect 4952 21732 4956 21788
rect 4956 21732 5012 21788
rect 5012 21732 5016 21788
rect 4952 21728 5016 21732
rect 5032 21788 5096 21792
rect 5032 21732 5036 21788
rect 5036 21732 5092 21788
rect 5092 21732 5096 21788
rect 5032 21728 5096 21732
rect 5112 21788 5176 21792
rect 5112 21732 5116 21788
rect 5116 21732 5172 21788
rect 5172 21732 5176 21788
rect 5112 21728 5176 21732
rect 5192 21788 5256 21792
rect 5192 21732 5196 21788
rect 5196 21732 5252 21788
rect 5252 21732 5256 21788
rect 5192 21728 5256 21732
rect 12952 21788 13016 21792
rect 12952 21732 12956 21788
rect 12956 21732 13012 21788
rect 13012 21732 13016 21788
rect 12952 21728 13016 21732
rect 13032 21788 13096 21792
rect 13032 21732 13036 21788
rect 13036 21732 13092 21788
rect 13092 21732 13096 21788
rect 13032 21728 13096 21732
rect 13112 21788 13176 21792
rect 13112 21732 13116 21788
rect 13116 21732 13172 21788
rect 13172 21732 13176 21788
rect 13112 21728 13176 21732
rect 13192 21788 13256 21792
rect 13192 21732 13196 21788
rect 13196 21732 13252 21788
rect 13252 21732 13256 21788
rect 13192 21728 13256 21732
rect 20952 21788 21016 21792
rect 20952 21732 20956 21788
rect 20956 21732 21012 21788
rect 21012 21732 21016 21788
rect 20952 21728 21016 21732
rect 21032 21788 21096 21792
rect 21032 21732 21036 21788
rect 21036 21732 21092 21788
rect 21092 21732 21096 21788
rect 21032 21728 21096 21732
rect 21112 21788 21176 21792
rect 21112 21732 21116 21788
rect 21116 21732 21172 21788
rect 21172 21732 21176 21788
rect 21112 21728 21176 21732
rect 21192 21788 21256 21792
rect 21192 21732 21196 21788
rect 21196 21732 21252 21788
rect 21252 21732 21256 21788
rect 21192 21728 21256 21732
rect 8952 21244 9016 21248
rect 8952 21188 8956 21244
rect 8956 21188 9012 21244
rect 9012 21188 9016 21244
rect 8952 21184 9016 21188
rect 9032 21244 9096 21248
rect 9032 21188 9036 21244
rect 9036 21188 9092 21244
rect 9092 21188 9096 21244
rect 9032 21184 9096 21188
rect 9112 21244 9176 21248
rect 9112 21188 9116 21244
rect 9116 21188 9172 21244
rect 9172 21188 9176 21244
rect 9112 21184 9176 21188
rect 9192 21244 9256 21248
rect 9192 21188 9196 21244
rect 9196 21188 9252 21244
rect 9252 21188 9256 21244
rect 9192 21184 9256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 4952 20700 5016 20704
rect 4952 20644 4956 20700
rect 4956 20644 5012 20700
rect 5012 20644 5016 20700
rect 4952 20640 5016 20644
rect 5032 20700 5096 20704
rect 5032 20644 5036 20700
rect 5036 20644 5092 20700
rect 5092 20644 5096 20700
rect 5032 20640 5096 20644
rect 5112 20700 5176 20704
rect 5112 20644 5116 20700
rect 5116 20644 5172 20700
rect 5172 20644 5176 20700
rect 5112 20640 5176 20644
rect 5192 20700 5256 20704
rect 5192 20644 5196 20700
rect 5196 20644 5252 20700
rect 5252 20644 5256 20700
rect 5192 20640 5256 20644
rect 12952 20700 13016 20704
rect 12952 20644 12956 20700
rect 12956 20644 13012 20700
rect 13012 20644 13016 20700
rect 12952 20640 13016 20644
rect 13032 20700 13096 20704
rect 13032 20644 13036 20700
rect 13036 20644 13092 20700
rect 13092 20644 13096 20700
rect 13032 20640 13096 20644
rect 13112 20700 13176 20704
rect 13112 20644 13116 20700
rect 13116 20644 13172 20700
rect 13172 20644 13176 20700
rect 13112 20640 13176 20644
rect 13192 20700 13256 20704
rect 13192 20644 13196 20700
rect 13196 20644 13252 20700
rect 13252 20644 13256 20700
rect 13192 20640 13256 20644
rect 20952 20700 21016 20704
rect 20952 20644 20956 20700
rect 20956 20644 21012 20700
rect 21012 20644 21016 20700
rect 20952 20640 21016 20644
rect 21032 20700 21096 20704
rect 21032 20644 21036 20700
rect 21036 20644 21092 20700
rect 21092 20644 21096 20700
rect 21032 20640 21096 20644
rect 21112 20700 21176 20704
rect 21112 20644 21116 20700
rect 21116 20644 21172 20700
rect 21172 20644 21176 20700
rect 21112 20640 21176 20644
rect 21192 20700 21256 20704
rect 21192 20644 21196 20700
rect 21196 20644 21252 20700
rect 21252 20644 21256 20700
rect 21192 20640 21256 20644
rect 8952 20156 9016 20160
rect 8952 20100 8956 20156
rect 8956 20100 9012 20156
rect 9012 20100 9016 20156
rect 8952 20096 9016 20100
rect 9032 20156 9096 20160
rect 9032 20100 9036 20156
rect 9036 20100 9092 20156
rect 9092 20100 9096 20156
rect 9032 20096 9096 20100
rect 9112 20156 9176 20160
rect 9112 20100 9116 20156
rect 9116 20100 9172 20156
rect 9172 20100 9176 20156
rect 9112 20096 9176 20100
rect 9192 20156 9256 20160
rect 9192 20100 9196 20156
rect 9196 20100 9252 20156
rect 9252 20100 9256 20156
rect 9192 20096 9256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 4952 19612 5016 19616
rect 4952 19556 4956 19612
rect 4956 19556 5012 19612
rect 5012 19556 5016 19612
rect 4952 19552 5016 19556
rect 5032 19612 5096 19616
rect 5032 19556 5036 19612
rect 5036 19556 5092 19612
rect 5092 19556 5096 19612
rect 5032 19552 5096 19556
rect 5112 19612 5176 19616
rect 5112 19556 5116 19612
rect 5116 19556 5172 19612
rect 5172 19556 5176 19612
rect 5112 19552 5176 19556
rect 5192 19612 5256 19616
rect 5192 19556 5196 19612
rect 5196 19556 5252 19612
rect 5252 19556 5256 19612
rect 5192 19552 5256 19556
rect 12952 19612 13016 19616
rect 12952 19556 12956 19612
rect 12956 19556 13012 19612
rect 13012 19556 13016 19612
rect 12952 19552 13016 19556
rect 13032 19612 13096 19616
rect 13032 19556 13036 19612
rect 13036 19556 13092 19612
rect 13092 19556 13096 19612
rect 13032 19552 13096 19556
rect 13112 19612 13176 19616
rect 13112 19556 13116 19612
rect 13116 19556 13172 19612
rect 13172 19556 13176 19612
rect 13112 19552 13176 19556
rect 13192 19612 13256 19616
rect 13192 19556 13196 19612
rect 13196 19556 13252 19612
rect 13252 19556 13256 19612
rect 13192 19552 13256 19556
rect 20952 19612 21016 19616
rect 20952 19556 20956 19612
rect 20956 19556 21012 19612
rect 21012 19556 21016 19612
rect 20952 19552 21016 19556
rect 21032 19612 21096 19616
rect 21032 19556 21036 19612
rect 21036 19556 21092 19612
rect 21092 19556 21096 19612
rect 21032 19552 21096 19556
rect 21112 19612 21176 19616
rect 21112 19556 21116 19612
rect 21116 19556 21172 19612
rect 21172 19556 21176 19612
rect 21112 19552 21176 19556
rect 21192 19612 21256 19616
rect 21192 19556 21196 19612
rect 21196 19556 21252 19612
rect 21252 19556 21256 19612
rect 21192 19552 21256 19556
rect 8952 19068 9016 19072
rect 8952 19012 8956 19068
rect 8956 19012 9012 19068
rect 9012 19012 9016 19068
rect 8952 19008 9016 19012
rect 9032 19068 9096 19072
rect 9032 19012 9036 19068
rect 9036 19012 9092 19068
rect 9092 19012 9096 19068
rect 9032 19008 9096 19012
rect 9112 19068 9176 19072
rect 9112 19012 9116 19068
rect 9116 19012 9172 19068
rect 9172 19012 9176 19068
rect 9112 19008 9176 19012
rect 9192 19068 9256 19072
rect 9192 19012 9196 19068
rect 9196 19012 9252 19068
rect 9252 19012 9256 19068
rect 9192 19008 9256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 4952 18524 5016 18528
rect 4952 18468 4956 18524
rect 4956 18468 5012 18524
rect 5012 18468 5016 18524
rect 4952 18464 5016 18468
rect 5032 18524 5096 18528
rect 5032 18468 5036 18524
rect 5036 18468 5092 18524
rect 5092 18468 5096 18524
rect 5032 18464 5096 18468
rect 5112 18524 5176 18528
rect 5112 18468 5116 18524
rect 5116 18468 5172 18524
rect 5172 18468 5176 18524
rect 5112 18464 5176 18468
rect 5192 18524 5256 18528
rect 5192 18468 5196 18524
rect 5196 18468 5252 18524
rect 5252 18468 5256 18524
rect 5192 18464 5256 18468
rect 12952 18524 13016 18528
rect 12952 18468 12956 18524
rect 12956 18468 13012 18524
rect 13012 18468 13016 18524
rect 12952 18464 13016 18468
rect 13032 18524 13096 18528
rect 13032 18468 13036 18524
rect 13036 18468 13092 18524
rect 13092 18468 13096 18524
rect 13032 18464 13096 18468
rect 13112 18524 13176 18528
rect 13112 18468 13116 18524
rect 13116 18468 13172 18524
rect 13172 18468 13176 18524
rect 13112 18464 13176 18468
rect 13192 18524 13256 18528
rect 13192 18468 13196 18524
rect 13196 18468 13252 18524
rect 13252 18468 13256 18524
rect 13192 18464 13256 18468
rect 20952 18524 21016 18528
rect 20952 18468 20956 18524
rect 20956 18468 21012 18524
rect 21012 18468 21016 18524
rect 20952 18464 21016 18468
rect 21032 18524 21096 18528
rect 21032 18468 21036 18524
rect 21036 18468 21092 18524
rect 21092 18468 21096 18524
rect 21032 18464 21096 18468
rect 21112 18524 21176 18528
rect 21112 18468 21116 18524
rect 21116 18468 21172 18524
rect 21172 18468 21176 18524
rect 21112 18464 21176 18468
rect 21192 18524 21256 18528
rect 21192 18468 21196 18524
rect 21196 18468 21252 18524
rect 21252 18468 21256 18524
rect 21192 18464 21256 18468
rect 8952 17980 9016 17984
rect 8952 17924 8956 17980
rect 8956 17924 9012 17980
rect 9012 17924 9016 17980
rect 8952 17920 9016 17924
rect 9032 17980 9096 17984
rect 9032 17924 9036 17980
rect 9036 17924 9092 17980
rect 9092 17924 9096 17980
rect 9032 17920 9096 17924
rect 9112 17980 9176 17984
rect 9112 17924 9116 17980
rect 9116 17924 9172 17980
rect 9172 17924 9176 17980
rect 9112 17920 9176 17924
rect 9192 17980 9256 17984
rect 9192 17924 9196 17980
rect 9196 17924 9252 17980
rect 9252 17924 9256 17980
rect 9192 17920 9256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 4952 17436 5016 17440
rect 4952 17380 4956 17436
rect 4956 17380 5012 17436
rect 5012 17380 5016 17436
rect 4952 17376 5016 17380
rect 5032 17436 5096 17440
rect 5032 17380 5036 17436
rect 5036 17380 5092 17436
rect 5092 17380 5096 17436
rect 5032 17376 5096 17380
rect 5112 17436 5176 17440
rect 5112 17380 5116 17436
rect 5116 17380 5172 17436
rect 5172 17380 5176 17436
rect 5112 17376 5176 17380
rect 5192 17436 5256 17440
rect 5192 17380 5196 17436
rect 5196 17380 5252 17436
rect 5252 17380 5256 17436
rect 5192 17376 5256 17380
rect 12952 17436 13016 17440
rect 12952 17380 12956 17436
rect 12956 17380 13012 17436
rect 13012 17380 13016 17436
rect 12952 17376 13016 17380
rect 13032 17436 13096 17440
rect 13032 17380 13036 17436
rect 13036 17380 13092 17436
rect 13092 17380 13096 17436
rect 13032 17376 13096 17380
rect 13112 17436 13176 17440
rect 13112 17380 13116 17436
rect 13116 17380 13172 17436
rect 13172 17380 13176 17436
rect 13112 17376 13176 17380
rect 13192 17436 13256 17440
rect 13192 17380 13196 17436
rect 13196 17380 13252 17436
rect 13252 17380 13256 17436
rect 13192 17376 13256 17380
rect 20952 17436 21016 17440
rect 20952 17380 20956 17436
rect 20956 17380 21012 17436
rect 21012 17380 21016 17436
rect 20952 17376 21016 17380
rect 21032 17436 21096 17440
rect 21032 17380 21036 17436
rect 21036 17380 21092 17436
rect 21092 17380 21096 17436
rect 21032 17376 21096 17380
rect 21112 17436 21176 17440
rect 21112 17380 21116 17436
rect 21116 17380 21172 17436
rect 21172 17380 21176 17436
rect 21112 17376 21176 17380
rect 21192 17436 21256 17440
rect 21192 17380 21196 17436
rect 21196 17380 21252 17436
rect 21252 17380 21256 17436
rect 21192 17376 21256 17380
rect 8952 16892 9016 16896
rect 8952 16836 8956 16892
rect 8956 16836 9012 16892
rect 9012 16836 9016 16892
rect 8952 16832 9016 16836
rect 9032 16892 9096 16896
rect 9032 16836 9036 16892
rect 9036 16836 9092 16892
rect 9092 16836 9096 16892
rect 9032 16832 9096 16836
rect 9112 16892 9176 16896
rect 9112 16836 9116 16892
rect 9116 16836 9172 16892
rect 9172 16836 9176 16892
rect 9112 16832 9176 16836
rect 9192 16892 9256 16896
rect 9192 16836 9196 16892
rect 9196 16836 9252 16892
rect 9252 16836 9256 16892
rect 9192 16832 9256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 4952 16348 5016 16352
rect 4952 16292 4956 16348
rect 4956 16292 5012 16348
rect 5012 16292 5016 16348
rect 4952 16288 5016 16292
rect 5032 16348 5096 16352
rect 5032 16292 5036 16348
rect 5036 16292 5092 16348
rect 5092 16292 5096 16348
rect 5032 16288 5096 16292
rect 5112 16348 5176 16352
rect 5112 16292 5116 16348
rect 5116 16292 5172 16348
rect 5172 16292 5176 16348
rect 5112 16288 5176 16292
rect 5192 16348 5256 16352
rect 5192 16292 5196 16348
rect 5196 16292 5252 16348
rect 5252 16292 5256 16348
rect 5192 16288 5256 16292
rect 12952 16348 13016 16352
rect 12952 16292 12956 16348
rect 12956 16292 13012 16348
rect 13012 16292 13016 16348
rect 12952 16288 13016 16292
rect 13032 16348 13096 16352
rect 13032 16292 13036 16348
rect 13036 16292 13092 16348
rect 13092 16292 13096 16348
rect 13032 16288 13096 16292
rect 13112 16348 13176 16352
rect 13112 16292 13116 16348
rect 13116 16292 13172 16348
rect 13172 16292 13176 16348
rect 13112 16288 13176 16292
rect 13192 16348 13256 16352
rect 13192 16292 13196 16348
rect 13196 16292 13252 16348
rect 13252 16292 13256 16348
rect 13192 16288 13256 16292
rect 20952 16348 21016 16352
rect 20952 16292 20956 16348
rect 20956 16292 21012 16348
rect 21012 16292 21016 16348
rect 20952 16288 21016 16292
rect 21032 16348 21096 16352
rect 21032 16292 21036 16348
rect 21036 16292 21092 16348
rect 21092 16292 21096 16348
rect 21032 16288 21096 16292
rect 21112 16348 21176 16352
rect 21112 16292 21116 16348
rect 21116 16292 21172 16348
rect 21172 16292 21176 16348
rect 21112 16288 21176 16292
rect 21192 16348 21256 16352
rect 21192 16292 21196 16348
rect 21196 16292 21252 16348
rect 21252 16292 21256 16348
rect 21192 16288 21256 16292
rect 8952 15804 9016 15808
rect 8952 15748 8956 15804
rect 8956 15748 9012 15804
rect 9012 15748 9016 15804
rect 8952 15744 9016 15748
rect 9032 15804 9096 15808
rect 9032 15748 9036 15804
rect 9036 15748 9092 15804
rect 9092 15748 9096 15804
rect 9032 15744 9096 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 4952 15260 5016 15264
rect 4952 15204 4956 15260
rect 4956 15204 5012 15260
rect 5012 15204 5016 15260
rect 4952 15200 5016 15204
rect 5032 15260 5096 15264
rect 5032 15204 5036 15260
rect 5036 15204 5092 15260
rect 5092 15204 5096 15260
rect 5032 15200 5096 15204
rect 5112 15260 5176 15264
rect 5112 15204 5116 15260
rect 5116 15204 5172 15260
rect 5172 15204 5176 15260
rect 5112 15200 5176 15204
rect 5192 15260 5256 15264
rect 5192 15204 5196 15260
rect 5196 15204 5252 15260
rect 5252 15204 5256 15260
rect 5192 15200 5256 15204
rect 12952 15260 13016 15264
rect 12952 15204 12956 15260
rect 12956 15204 13012 15260
rect 13012 15204 13016 15260
rect 12952 15200 13016 15204
rect 13032 15260 13096 15264
rect 13032 15204 13036 15260
rect 13036 15204 13092 15260
rect 13092 15204 13096 15260
rect 13032 15200 13096 15204
rect 13112 15260 13176 15264
rect 13112 15204 13116 15260
rect 13116 15204 13172 15260
rect 13172 15204 13176 15260
rect 13112 15200 13176 15204
rect 13192 15260 13256 15264
rect 13192 15204 13196 15260
rect 13196 15204 13252 15260
rect 13252 15204 13256 15260
rect 13192 15200 13256 15204
rect 20952 15260 21016 15264
rect 20952 15204 20956 15260
rect 20956 15204 21012 15260
rect 21012 15204 21016 15260
rect 20952 15200 21016 15204
rect 21032 15260 21096 15264
rect 21032 15204 21036 15260
rect 21036 15204 21092 15260
rect 21092 15204 21096 15260
rect 21032 15200 21096 15204
rect 21112 15260 21176 15264
rect 21112 15204 21116 15260
rect 21116 15204 21172 15260
rect 21172 15204 21176 15260
rect 21112 15200 21176 15204
rect 21192 15260 21256 15264
rect 21192 15204 21196 15260
rect 21196 15204 21252 15260
rect 21252 15204 21256 15260
rect 21192 15200 21256 15204
rect 8952 14716 9016 14720
rect 8952 14660 8956 14716
rect 8956 14660 9012 14716
rect 9012 14660 9016 14716
rect 8952 14656 9016 14660
rect 9032 14716 9096 14720
rect 9032 14660 9036 14716
rect 9036 14660 9092 14716
rect 9092 14660 9096 14716
rect 9032 14656 9096 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 4952 14172 5016 14176
rect 4952 14116 4956 14172
rect 4956 14116 5012 14172
rect 5012 14116 5016 14172
rect 4952 14112 5016 14116
rect 5032 14172 5096 14176
rect 5032 14116 5036 14172
rect 5036 14116 5092 14172
rect 5092 14116 5096 14172
rect 5032 14112 5096 14116
rect 5112 14172 5176 14176
rect 5112 14116 5116 14172
rect 5116 14116 5172 14172
rect 5172 14116 5176 14172
rect 5112 14112 5176 14116
rect 5192 14172 5256 14176
rect 5192 14116 5196 14172
rect 5196 14116 5252 14172
rect 5252 14116 5256 14172
rect 5192 14112 5256 14116
rect 12952 14172 13016 14176
rect 12952 14116 12956 14172
rect 12956 14116 13012 14172
rect 13012 14116 13016 14172
rect 12952 14112 13016 14116
rect 13032 14172 13096 14176
rect 13032 14116 13036 14172
rect 13036 14116 13092 14172
rect 13092 14116 13096 14172
rect 13032 14112 13096 14116
rect 13112 14172 13176 14176
rect 13112 14116 13116 14172
rect 13116 14116 13172 14172
rect 13172 14116 13176 14172
rect 13112 14112 13176 14116
rect 13192 14172 13256 14176
rect 13192 14116 13196 14172
rect 13196 14116 13252 14172
rect 13252 14116 13256 14172
rect 13192 14112 13256 14116
rect 20952 14172 21016 14176
rect 20952 14116 20956 14172
rect 20956 14116 21012 14172
rect 21012 14116 21016 14172
rect 20952 14112 21016 14116
rect 21032 14172 21096 14176
rect 21032 14116 21036 14172
rect 21036 14116 21092 14172
rect 21092 14116 21096 14172
rect 21032 14112 21096 14116
rect 21112 14172 21176 14176
rect 21112 14116 21116 14172
rect 21116 14116 21172 14172
rect 21172 14116 21176 14172
rect 21112 14112 21176 14116
rect 21192 14172 21256 14176
rect 21192 14116 21196 14172
rect 21196 14116 21252 14172
rect 21252 14116 21256 14172
rect 21192 14112 21256 14116
rect 8952 13628 9016 13632
rect 8952 13572 8956 13628
rect 8956 13572 9012 13628
rect 9012 13572 9016 13628
rect 8952 13568 9016 13572
rect 9032 13628 9096 13632
rect 9032 13572 9036 13628
rect 9036 13572 9092 13628
rect 9092 13572 9096 13628
rect 9032 13568 9096 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 4952 13084 5016 13088
rect 4952 13028 4956 13084
rect 4956 13028 5012 13084
rect 5012 13028 5016 13084
rect 4952 13024 5016 13028
rect 5032 13084 5096 13088
rect 5032 13028 5036 13084
rect 5036 13028 5092 13084
rect 5092 13028 5096 13084
rect 5032 13024 5096 13028
rect 5112 13084 5176 13088
rect 5112 13028 5116 13084
rect 5116 13028 5172 13084
rect 5172 13028 5176 13084
rect 5112 13024 5176 13028
rect 5192 13084 5256 13088
rect 5192 13028 5196 13084
rect 5196 13028 5252 13084
rect 5252 13028 5256 13084
rect 5192 13024 5256 13028
rect 12952 13084 13016 13088
rect 12952 13028 12956 13084
rect 12956 13028 13012 13084
rect 13012 13028 13016 13084
rect 12952 13024 13016 13028
rect 13032 13084 13096 13088
rect 13032 13028 13036 13084
rect 13036 13028 13092 13084
rect 13092 13028 13096 13084
rect 13032 13024 13096 13028
rect 13112 13084 13176 13088
rect 13112 13028 13116 13084
rect 13116 13028 13172 13084
rect 13172 13028 13176 13084
rect 13112 13024 13176 13028
rect 13192 13084 13256 13088
rect 13192 13028 13196 13084
rect 13196 13028 13252 13084
rect 13252 13028 13256 13084
rect 13192 13024 13256 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 8952 12540 9016 12544
rect 8952 12484 8956 12540
rect 8956 12484 9012 12540
rect 9012 12484 9016 12540
rect 8952 12480 9016 12484
rect 9032 12540 9096 12544
rect 9032 12484 9036 12540
rect 9036 12484 9092 12540
rect 9092 12484 9096 12540
rect 9032 12480 9096 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 4952 11996 5016 12000
rect 4952 11940 4956 11996
rect 4956 11940 5012 11996
rect 5012 11940 5016 11996
rect 4952 11936 5016 11940
rect 5032 11996 5096 12000
rect 5032 11940 5036 11996
rect 5036 11940 5092 11996
rect 5092 11940 5096 11996
rect 5032 11936 5096 11940
rect 5112 11996 5176 12000
rect 5112 11940 5116 11996
rect 5116 11940 5172 11996
rect 5172 11940 5176 11996
rect 5112 11936 5176 11940
rect 5192 11996 5256 12000
rect 5192 11940 5196 11996
rect 5196 11940 5252 11996
rect 5252 11940 5256 11996
rect 5192 11936 5256 11940
rect 12952 11996 13016 12000
rect 12952 11940 12956 11996
rect 12956 11940 13012 11996
rect 13012 11940 13016 11996
rect 12952 11936 13016 11940
rect 13032 11996 13096 12000
rect 13032 11940 13036 11996
rect 13036 11940 13092 11996
rect 13092 11940 13096 11996
rect 13032 11936 13096 11940
rect 13112 11996 13176 12000
rect 13112 11940 13116 11996
rect 13116 11940 13172 11996
rect 13172 11940 13176 11996
rect 13112 11936 13176 11940
rect 13192 11996 13256 12000
rect 13192 11940 13196 11996
rect 13196 11940 13252 11996
rect 13252 11940 13256 11996
rect 13192 11936 13256 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 8952 11452 9016 11456
rect 8952 11396 8956 11452
rect 8956 11396 9012 11452
rect 9012 11396 9016 11452
rect 8952 11392 9016 11396
rect 9032 11452 9096 11456
rect 9032 11396 9036 11452
rect 9036 11396 9092 11452
rect 9092 11396 9096 11452
rect 9032 11392 9096 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 4952 10908 5016 10912
rect 4952 10852 4956 10908
rect 4956 10852 5012 10908
rect 5012 10852 5016 10908
rect 4952 10848 5016 10852
rect 5032 10908 5096 10912
rect 5032 10852 5036 10908
rect 5036 10852 5092 10908
rect 5092 10852 5096 10908
rect 5032 10848 5096 10852
rect 5112 10908 5176 10912
rect 5112 10852 5116 10908
rect 5116 10852 5172 10908
rect 5172 10852 5176 10908
rect 5112 10848 5176 10852
rect 5192 10908 5256 10912
rect 5192 10852 5196 10908
rect 5196 10852 5252 10908
rect 5252 10852 5256 10908
rect 5192 10848 5256 10852
rect 12952 10908 13016 10912
rect 12952 10852 12956 10908
rect 12956 10852 13012 10908
rect 13012 10852 13016 10908
rect 12952 10848 13016 10852
rect 13032 10908 13096 10912
rect 13032 10852 13036 10908
rect 13036 10852 13092 10908
rect 13092 10852 13096 10908
rect 13032 10848 13096 10852
rect 13112 10908 13176 10912
rect 13112 10852 13116 10908
rect 13116 10852 13172 10908
rect 13172 10852 13176 10908
rect 13112 10848 13176 10852
rect 13192 10908 13256 10912
rect 13192 10852 13196 10908
rect 13196 10852 13252 10908
rect 13252 10852 13256 10908
rect 13192 10848 13256 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 8952 10364 9016 10368
rect 8952 10308 8956 10364
rect 8956 10308 9012 10364
rect 9012 10308 9016 10364
rect 8952 10304 9016 10308
rect 9032 10364 9096 10368
rect 9032 10308 9036 10364
rect 9036 10308 9092 10364
rect 9092 10308 9096 10364
rect 9032 10304 9096 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 4952 9820 5016 9824
rect 4952 9764 4956 9820
rect 4956 9764 5012 9820
rect 5012 9764 5016 9820
rect 4952 9760 5016 9764
rect 5032 9820 5096 9824
rect 5032 9764 5036 9820
rect 5036 9764 5092 9820
rect 5092 9764 5096 9820
rect 5032 9760 5096 9764
rect 5112 9820 5176 9824
rect 5112 9764 5116 9820
rect 5116 9764 5172 9820
rect 5172 9764 5176 9820
rect 5112 9760 5176 9764
rect 5192 9820 5256 9824
rect 5192 9764 5196 9820
rect 5196 9764 5252 9820
rect 5252 9764 5256 9820
rect 5192 9760 5256 9764
rect 12952 9820 13016 9824
rect 12952 9764 12956 9820
rect 12956 9764 13012 9820
rect 13012 9764 13016 9820
rect 12952 9760 13016 9764
rect 13032 9820 13096 9824
rect 13032 9764 13036 9820
rect 13036 9764 13092 9820
rect 13092 9764 13096 9820
rect 13032 9760 13096 9764
rect 13112 9820 13176 9824
rect 13112 9764 13116 9820
rect 13116 9764 13172 9820
rect 13172 9764 13176 9820
rect 13112 9760 13176 9764
rect 13192 9820 13256 9824
rect 13192 9764 13196 9820
rect 13196 9764 13252 9820
rect 13252 9764 13256 9820
rect 13192 9760 13256 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 8952 9276 9016 9280
rect 8952 9220 8956 9276
rect 8956 9220 9012 9276
rect 9012 9220 9016 9276
rect 8952 9216 9016 9220
rect 9032 9276 9096 9280
rect 9032 9220 9036 9276
rect 9036 9220 9092 9276
rect 9092 9220 9096 9276
rect 9032 9216 9096 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 4952 8732 5016 8736
rect 4952 8676 4956 8732
rect 4956 8676 5012 8732
rect 5012 8676 5016 8732
rect 4952 8672 5016 8676
rect 5032 8732 5096 8736
rect 5032 8676 5036 8732
rect 5036 8676 5092 8732
rect 5092 8676 5096 8732
rect 5032 8672 5096 8676
rect 5112 8732 5176 8736
rect 5112 8676 5116 8732
rect 5116 8676 5172 8732
rect 5172 8676 5176 8732
rect 5112 8672 5176 8676
rect 5192 8732 5256 8736
rect 5192 8676 5196 8732
rect 5196 8676 5252 8732
rect 5252 8676 5256 8732
rect 5192 8672 5256 8676
rect 12952 8732 13016 8736
rect 12952 8676 12956 8732
rect 12956 8676 13012 8732
rect 13012 8676 13016 8732
rect 12952 8672 13016 8676
rect 13032 8732 13096 8736
rect 13032 8676 13036 8732
rect 13036 8676 13092 8732
rect 13092 8676 13096 8732
rect 13032 8672 13096 8676
rect 13112 8732 13176 8736
rect 13112 8676 13116 8732
rect 13116 8676 13172 8732
rect 13172 8676 13176 8732
rect 13112 8672 13176 8676
rect 13192 8732 13256 8736
rect 13192 8676 13196 8732
rect 13196 8676 13252 8732
rect 13252 8676 13256 8732
rect 13192 8672 13256 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 8952 8188 9016 8192
rect 8952 8132 8956 8188
rect 8956 8132 9012 8188
rect 9012 8132 9016 8188
rect 8952 8128 9016 8132
rect 9032 8188 9096 8192
rect 9032 8132 9036 8188
rect 9036 8132 9092 8188
rect 9092 8132 9096 8188
rect 9032 8128 9096 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 4952 7644 5016 7648
rect 4952 7588 4956 7644
rect 4956 7588 5012 7644
rect 5012 7588 5016 7644
rect 4952 7584 5016 7588
rect 5032 7644 5096 7648
rect 5032 7588 5036 7644
rect 5036 7588 5092 7644
rect 5092 7588 5096 7644
rect 5032 7584 5096 7588
rect 5112 7644 5176 7648
rect 5112 7588 5116 7644
rect 5116 7588 5172 7644
rect 5172 7588 5176 7644
rect 5112 7584 5176 7588
rect 5192 7644 5256 7648
rect 5192 7588 5196 7644
rect 5196 7588 5252 7644
rect 5252 7588 5256 7644
rect 5192 7584 5256 7588
rect 12952 7644 13016 7648
rect 12952 7588 12956 7644
rect 12956 7588 13012 7644
rect 13012 7588 13016 7644
rect 12952 7584 13016 7588
rect 13032 7644 13096 7648
rect 13032 7588 13036 7644
rect 13036 7588 13092 7644
rect 13092 7588 13096 7644
rect 13032 7584 13096 7588
rect 13112 7644 13176 7648
rect 13112 7588 13116 7644
rect 13116 7588 13172 7644
rect 13172 7588 13176 7644
rect 13112 7584 13176 7588
rect 13192 7644 13256 7648
rect 13192 7588 13196 7644
rect 13196 7588 13252 7644
rect 13252 7588 13256 7644
rect 13192 7584 13256 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 8952 7100 9016 7104
rect 8952 7044 8956 7100
rect 8956 7044 9012 7100
rect 9012 7044 9016 7100
rect 8952 7040 9016 7044
rect 9032 7100 9096 7104
rect 9032 7044 9036 7100
rect 9036 7044 9092 7100
rect 9092 7044 9096 7100
rect 9032 7040 9096 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 4952 6556 5016 6560
rect 4952 6500 4956 6556
rect 4956 6500 5012 6556
rect 5012 6500 5016 6556
rect 4952 6496 5016 6500
rect 5032 6556 5096 6560
rect 5032 6500 5036 6556
rect 5036 6500 5092 6556
rect 5092 6500 5096 6556
rect 5032 6496 5096 6500
rect 5112 6556 5176 6560
rect 5112 6500 5116 6556
rect 5116 6500 5172 6556
rect 5172 6500 5176 6556
rect 5112 6496 5176 6500
rect 5192 6556 5256 6560
rect 5192 6500 5196 6556
rect 5196 6500 5252 6556
rect 5252 6500 5256 6556
rect 5192 6496 5256 6500
rect 12952 6556 13016 6560
rect 12952 6500 12956 6556
rect 12956 6500 13012 6556
rect 13012 6500 13016 6556
rect 12952 6496 13016 6500
rect 13032 6556 13096 6560
rect 13032 6500 13036 6556
rect 13036 6500 13092 6556
rect 13092 6500 13096 6556
rect 13032 6496 13096 6500
rect 13112 6556 13176 6560
rect 13112 6500 13116 6556
rect 13116 6500 13172 6556
rect 13172 6500 13176 6556
rect 13112 6496 13176 6500
rect 13192 6556 13256 6560
rect 13192 6500 13196 6556
rect 13196 6500 13252 6556
rect 13252 6500 13256 6556
rect 13192 6496 13256 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 8952 6012 9016 6016
rect 8952 5956 8956 6012
rect 8956 5956 9012 6012
rect 9012 5956 9016 6012
rect 8952 5952 9016 5956
rect 9032 6012 9096 6016
rect 9032 5956 9036 6012
rect 9036 5956 9092 6012
rect 9092 5956 9096 6012
rect 9032 5952 9096 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 4952 5468 5016 5472
rect 4952 5412 4956 5468
rect 4956 5412 5012 5468
rect 5012 5412 5016 5468
rect 4952 5408 5016 5412
rect 5032 5468 5096 5472
rect 5032 5412 5036 5468
rect 5036 5412 5092 5468
rect 5092 5412 5096 5468
rect 5032 5408 5096 5412
rect 5112 5468 5176 5472
rect 5112 5412 5116 5468
rect 5116 5412 5172 5468
rect 5172 5412 5176 5468
rect 5112 5408 5176 5412
rect 5192 5468 5256 5472
rect 5192 5412 5196 5468
rect 5196 5412 5252 5468
rect 5252 5412 5256 5468
rect 5192 5408 5256 5412
rect 12952 5468 13016 5472
rect 12952 5412 12956 5468
rect 12956 5412 13012 5468
rect 13012 5412 13016 5468
rect 12952 5408 13016 5412
rect 13032 5468 13096 5472
rect 13032 5412 13036 5468
rect 13036 5412 13092 5468
rect 13092 5412 13096 5468
rect 13032 5408 13096 5412
rect 13112 5468 13176 5472
rect 13112 5412 13116 5468
rect 13116 5412 13172 5468
rect 13172 5412 13176 5468
rect 13112 5408 13176 5412
rect 13192 5468 13256 5472
rect 13192 5412 13196 5468
rect 13196 5412 13252 5468
rect 13252 5412 13256 5468
rect 13192 5408 13256 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 8952 4924 9016 4928
rect 8952 4868 8956 4924
rect 8956 4868 9012 4924
rect 9012 4868 9016 4924
rect 8952 4864 9016 4868
rect 9032 4924 9096 4928
rect 9032 4868 9036 4924
rect 9036 4868 9092 4924
rect 9092 4868 9096 4924
rect 9032 4864 9096 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 4952 4380 5016 4384
rect 4952 4324 4956 4380
rect 4956 4324 5012 4380
rect 5012 4324 5016 4380
rect 4952 4320 5016 4324
rect 5032 4380 5096 4384
rect 5032 4324 5036 4380
rect 5036 4324 5092 4380
rect 5092 4324 5096 4380
rect 5032 4320 5096 4324
rect 5112 4380 5176 4384
rect 5112 4324 5116 4380
rect 5116 4324 5172 4380
rect 5172 4324 5176 4380
rect 5112 4320 5176 4324
rect 5192 4380 5256 4384
rect 5192 4324 5196 4380
rect 5196 4324 5252 4380
rect 5252 4324 5256 4380
rect 5192 4320 5256 4324
rect 12952 4380 13016 4384
rect 12952 4324 12956 4380
rect 12956 4324 13012 4380
rect 13012 4324 13016 4380
rect 12952 4320 13016 4324
rect 13032 4380 13096 4384
rect 13032 4324 13036 4380
rect 13036 4324 13092 4380
rect 13092 4324 13096 4380
rect 13032 4320 13096 4324
rect 13112 4380 13176 4384
rect 13112 4324 13116 4380
rect 13116 4324 13172 4380
rect 13172 4324 13176 4380
rect 13112 4320 13176 4324
rect 13192 4380 13256 4384
rect 13192 4324 13196 4380
rect 13196 4324 13252 4380
rect 13252 4324 13256 4380
rect 13192 4320 13256 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 8952 3836 9016 3840
rect 8952 3780 8956 3836
rect 8956 3780 9012 3836
rect 9012 3780 9016 3836
rect 8952 3776 9016 3780
rect 9032 3836 9096 3840
rect 9032 3780 9036 3836
rect 9036 3780 9092 3836
rect 9092 3780 9096 3836
rect 9032 3776 9096 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 4952 3292 5016 3296
rect 4952 3236 4956 3292
rect 4956 3236 5012 3292
rect 5012 3236 5016 3292
rect 4952 3232 5016 3236
rect 5032 3292 5096 3296
rect 5032 3236 5036 3292
rect 5036 3236 5092 3292
rect 5092 3236 5096 3292
rect 5032 3232 5096 3236
rect 5112 3292 5176 3296
rect 5112 3236 5116 3292
rect 5116 3236 5172 3292
rect 5172 3236 5176 3292
rect 5112 3232 5176 3236
rect 5192 3292 5256 3296
rect 5192 3236 5196 3292
rect 5196 3236 5252 3292
rect 5252 3236 5256 3292
rect 5192 3232 5256 3236
rect 12952 3292 13016 3296
rect 12952 3236 12956 3292
rect 12956 3236 13012 3292
rect 13012 3236 13016 3292
rect 12952 3232 13016 3236
rect 13032 3292 13096 3296
rect 13032 3236 13036 3292
rect 13036 3236 13092 3292
rect 13092 3236 13096 3292
rect 13032 3232 13096 3236
rect 13112 3292 13176 3296
rect 13112 3236 13116 3292
rect 13116 3236 13172 3292
rect 13172 3236 13176 3292
rect 13112 3232 13176 3236
rect 13192 3292 13256 3296
rect 13192 3236 13196 3292
rect 13196 3236 13252 3292
rect 13252 3236 13256 3292
rect 13192 3232 13256 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 8952 2748 9016 2752
rect 8952 2692 8956 2748
rect 8956 2692 9012 2748
rect 9012 2692 9016 2748
rect 8952 2688 9016 2692
rect 9032 2748 9096 2752
rect 9032 2692 9036 2748
rect 9036 2692 9092 2748
rect 9092 2692 9096 2748
rect 9032 2688 9096 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 4952 2204 5016 2208
rect 4952 2148 4956 2204
rect 4956 2148 5012 2204
rect 5012 2148 5016 2204
rect 4952 2144 5016 2148
rect 5032 2204 5096 2208
rect 5032 2148 5036 2204
rect 5036 2148 5092 2204
rect 5092 2148 5096 2204
rect 5032 2144 5096 2148
rect 5112 2204 5176 2208
rect 5112 2148 5116 2204
rect 5116 2148 5172 2204
rect 5172 2148 5176 2204
rect 5112 2144 5176 2148
rect 5192 2204 5256 2208
rect 5192 2148 5196 2204
rect 5196 2148 5252 2204
rect 5252 2148 5256 2204
rect 5192 2144 5256 2148
rect 12952 2204 13016 2208
rect 12952 2148 12956 2204
rect 12956 2148 13012 2204
rect 13012 2148 13016 2204
rect 12952 2144 13016 2148
rect 13032 2204 13096 2208
rect 13032 2148 13036 2204
rect 13036 2148 13092 2204
rect 13092 2148 13096 2204
rect 13032 2144 13096 2148
rect 13112 2204 13176 2208
rect 13112 2148 13116 2204
rect 13116 2148 13172 2204
rect 13172 2148 13176 2204
rect 13112 2144 13176 2148
rect 13192 2204 13256 2208
rect 13192 2148 13196 2204
rect 13196 2148 13252 2204
rect 13252 2148 13256 2204
rect 13192 2144 13256 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
<< metal4 >>
rect 4944 21792 5264 21808
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 20704 5264 21728
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 19616 5264 20640
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 18528 5264 19552
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 17440 5264 18464
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 16352 5264 17376
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 15264 5264 16288
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 14176 5264 15200
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 13088 5264 14112
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 12000 5264 13024
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 10912 5264 11936
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 9824 5264 10848
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 8736 5264 9760
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 7648 5264 8672
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 6560 5264 7584
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 5472 5264 6496
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 4384 5264 5408
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 3296 5264 4320
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 2208 5264 3232
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2128 5264 2144
rect 8944 21248 9264 21808
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 20160 9264 21184
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 19072 9264 20096
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 17984 9264 19008
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 16896 9264 17920
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 15808 9264 16832
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 14720 9264 15744
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 13632 9264 14656
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 12544 9264 13568
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 11456 9264 12480
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 10368 9264 11392
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 9280 9264 10304
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 8192 9264 9216
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 7104 9264 8128
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 6016 9264 7040
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 4928 9264 5952
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 3840 9264 4864
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 2752 9264 3776
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2128 9264 2688
rect 12944 21792 13264 21808
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 20704 13264 21728
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 19616 13264 20640
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 18528 13264 19552
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 17440 13264 18464
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 16352 13264 17376
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 15264 13264 16288
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 14176 13264 15200
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 13088 13264 14112
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 12000 13264 13024
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 10912 13264 11936
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 9824 13264 10848
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 8736 13264 9760
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 7648 13264 8672
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 6560 13264 7584
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 5472 13264 6496
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 4384 13264 5408
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 3296 13264 4320
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 2208 13264 3232
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2128 13264 2144
rect 16944 21248 17264 21808
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 17984 17264 19008
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 12544 17264 13568
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8192 17264 9216
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 7104 17264 8128
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 2752 17264 3776
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2128 17264 2688
rect 20944 21792 21264 21808
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 20704 21264 21728
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 19616 21264 20640
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 18528 21264 19552
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 17440 21264 18464
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 16352 21264 17376
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 15264 21264 16288
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 14176 21264 15200
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 13088 21264 14112
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
use scs8hd_fill_2  FILLER_1_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_10
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_9
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use scs8hd_nand2_4  _126_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_22
timestamp 1586364061
transform 1 0 3128 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_23
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_44 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_43
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_47
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_47
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_52
timestamp 1586364061
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _184_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_60
timestamp 1586364061
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_56
timestamp 1586364061
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_80
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_70
timestamp 1586364061
transform 1 0 7544 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_4  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_87
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_91
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_110
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_104
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_108
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_123
timestamp 1586364061
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_119
timestamp 1586364061
transform 1 0 12052 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_8  _119_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _203_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 590 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_141
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_145 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_146
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_150
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_153
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_161
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _194_
timestamp 1586364061
transform 1 0 16284 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_164
timestamp 1586364061
transform 1 0 16192 0 -1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_172
timestamp 1586364061
transform 1 0 16928 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_168
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_173
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_181
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_187
timestamp 1586364061
transform 1 0 18308 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _211_
timestamp 1586364061
transform 1 0 18584 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_191 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_194
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_198
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_204
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_203
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_215
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 22816 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 22816 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_227
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 590 592
use scs8hd_inv_8  _083_
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 4508 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_35
timestamp 1586364061
transform 1 0 4324 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_39
timestamp 1586364061
transform 1 0 4692 0 -1 3808
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_66
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_81
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_85
timestamp 1586364061
transform 1 0 8924 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_89
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_113
timestamp 1586364061
transform 1 0 11500 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_8  _106_
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_143
timestamp 1586364061
transform 1 0 14260 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _092_
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_4  FILLER_2_167
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_180
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_184
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_196
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_208
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 22816 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 590 592
use scs8hd_or2_4  _122_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 1 3808
box -38 -48 682 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_20
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_24
timestamp 1586364061
transform 1 0 3312 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_50
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_54
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 406 592
use scs8hd_nor3_4  _177_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__177__C
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_58
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__C
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_81
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_102
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_106
timestamp 1586364061
transform 1 0 10856 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_153
timestamp 1586364061
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_157
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_170
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_205
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 22816 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_229
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _160_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 4508 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__173__C
timestamp 1586364061
transform 1 0 4324 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_46
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_63
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_nor3_4  _176_
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 1234 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 9752 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_103
timestamp 1586364061
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_122
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_126
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_4_133
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_138
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_152
timestamp 1586364061
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_8  _091_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  FILLER_4_171
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_183
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_187
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_211
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 22816 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 590 592
use scs8hd_or2_4  _121_
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 682 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 3404 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_17
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_21
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_or4_4  _158_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__173__D
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_55
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__C
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_65
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_69
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _120_
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_73
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_90
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_93
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_or4_4  _155_
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_106
timestamp 1586364061
transform 1 0 10856 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__C
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__D
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_126
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_130
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_5_145
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_168
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_180
timestamp 1586364061
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 22816 0 1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 130 592
use scs8hd_inv_8  _104_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 5984
box -38 -48 866 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_12
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_13
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_17
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_16
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _178_
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_21
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use scs8hd_nand2_4  _148_
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 866 592
use scs8hd_or4_4  _173_
timestamp 1586364061
transform 1 0 4324 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_44
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_48
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_55
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__D
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _107_
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 6992 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_61
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_69
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 314 592
use scs8hd_nor3_4  _175_
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 1234 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_73
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__D
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_84
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_or4_4  _133_
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_106
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_103
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_107
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _105_
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_118
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_4  FILLER_7_111
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_115
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_133
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_6_146
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_159
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_153
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_165
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_171
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_177
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_183
timestamp 1586364061
transform 1 0 17940 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_195
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_6_207
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 22816 0 1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_17
timestamp 1586364061
transform 1 0 2668 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_21
timestamp 1586364061
transform 1 0 3036 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__C
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 774 592
use scs8hd_nor3_4  _174_
timestamp 1586364061
transform 1 0 5888 0 -1 7072
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_49
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_82
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_90
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 11684 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_114
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_118
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_122
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_1  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_135
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_147
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 22816 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_13
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_17
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_24
timestamp 1586364061
transform 1 0 3312 0 1 7072
box -38 -48 314 592
use scs8hd_or4_4  _152_
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_29
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__D
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_42
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_46
timestamp 1586364061
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_90
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _118_
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 866 592
use scs8hd_decap_6  FILLER_9_107
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_116
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_120
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_137
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_148
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_152
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_164
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_176
timestamp 1586364061
transform 1 0 17296 0 1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_182
timestamp 1586364061
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_211
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_218
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_222
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_230
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_16
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_20
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_24
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_28
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use scs8hd_conb_1  _181_
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_43
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_47
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_51
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_57
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_61
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_74
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_8  _115_
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_106
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 11592 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_10_123
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_130
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_142
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_150
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_200
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_212
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 22816 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_13
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_17
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_21
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_35
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _117_
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_73
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_77
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 774 592
use scs8hd_conb_1  _180_
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_85
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_97
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_150
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_162
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_182
timestamp 1586364061
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 22816 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 130 592
use scs8hd_inv_8  _103_
timestamp 1586364061
transform 1 0 1472 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_13
timestamp 1586364061
transform 1 0 2300 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_19
timestamp 1586364061
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_35
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_39
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__D
timestamp 1586364061
transform 1 0 6072 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_52
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _172_
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_60
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_12_77
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_89
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_104
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_108
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_120
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 1142 592
use scs8hd_inv_8  _084_
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_12_132
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use scs8hd_inv_8  _097_
timestamp 1586364061
transform 1 0 2668 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_26
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__D
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_38
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_8  _116_
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 866 592
use scs8hd_or4_4  _164_
timestamp 1586364061
transform 1 0 5980 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__D
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_42
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_52
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_45
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_49
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_62
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_60
timestamp 1586364061
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_56
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_66
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 1050 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_81
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_70
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_85
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_91
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_8  _082_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_106
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_106
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_110
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_8  _099_
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 866 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_126
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_130
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_130
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_134
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_152
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_4  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_164
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 590 592
use scs8hd_inv_8  _096_
timestamp 1586364061
transform 1 0 17020 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_172
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_182
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_198
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 22816 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 590 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_32
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_37
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_41
timestamp 1586364061
transform 1 0 4876 0 1 10336
box -38 -48 130 592
use scs8hd_or4_4  _142_
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _098_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _170_
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_88
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_92
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_96
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _146_
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_100
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_134
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 590 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_144
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_172
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_198
timestamp 1586364061
transform 1 0 19320 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_210
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 22816 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use scs8hd_or4_4  _161_
timestamp 1586364061
transform 1 0 4324 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__C
timestamp 1586364061
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_48
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_63
timestamp 1586364061
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_67
timestamp 1586364061
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__C
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_74
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _139_
timestamp 1586364061
transform 1 0 9752 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__D
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__D
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_103
timestamp 1586364061
transform 1 0 10580 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_107
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_16_122
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_127
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_139
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15548 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_168
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_176
timestamp 1586364061
transform 1 0 17296 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_188
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_192
timestamp 1586364061
transform 1 0 18768 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 19136 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_205
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_219
timestamp 1586364061
transform 1 0 21252 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 22816 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_231
timestamp 1586364061
transform 1 0 22356 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_25
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_29
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_36
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_40
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_90
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_94
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _145_
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_107
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__C
timestamp 1586364061
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__D
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_111
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_115
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_119
timestamp 1586364061
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_127
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_131
timestamp 1586364061
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_148
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_167
timestamp 1586364061
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_195
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_199
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_17_206
timestamp 1586364061
transform 1 0 20056 0 1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_217
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_221
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 22816 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_225
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_19
timestamp 1586364061
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 590 592
use scs8hd_inv_8  _086_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_50
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_53
timestamp 1586364061
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_66
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _136_
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_70
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _127_
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_106
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_121
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_18_126
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_137
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 14720 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_147
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_150
timestamp 1586364061
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17572 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_182
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_188
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_211
timestamp 1586364061
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_219
timestamp 1586364061
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 22816 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_231
timestamp 1586364061
transform 1 0 22356 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_8
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_25
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_20
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_24
timestamp 1586364061
transform 1 0 3312 0 -1 13600
box -38 -48 406 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_29
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_28
timestamp 1586364061
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 866 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_46
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_62
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_66
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_90
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 406 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_97
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_100
timestamp 1586364061
transform 1 0 10304 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_115
timestamp 1586364061
transform 1 0 11684 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_111
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 1050 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_127
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_130
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_134
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_8  _114_
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_157
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_161
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_167
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_179
timestamp 1586364061
transform 1 0 17572 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17756 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_201
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_213
timestamp 1586364061
transform 1 0 20700 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 22816 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 22816 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_19_225
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 774 592
use scs8hd_decap_6  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 590 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_14
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_22
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_25
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_38
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_42
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_49
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7452 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_21_80
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_or4_4  _167_
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_101
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_139
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_21_151
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_167
timestamp 1586364061
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _179_
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_204
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 22816 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_22_43
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_51
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_63
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use scs8hd_conb_1  _193_
timestamp 1586364061
transform 1 0 8372 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_75
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_90
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_110
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__D
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_123
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_8  _102_
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_128
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_132
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_146
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_158
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_177
timestamp 1586364061
transform 1 0 17388 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 866 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_194
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 22816 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_16
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_20
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_24
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_44
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_55
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_93
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_134
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_138
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_151
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_163
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18768 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_195
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_199
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_211
timestamp 1586364061
transform 1 0 20516 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 22816 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_223
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_231
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__213__A
timestamp 1586364061
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_11
timestamp 1586364061
transform 1 0 2116 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_21
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _163_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_29
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5888 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_63
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10304 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_115
timestamp 1586364061
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_119
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 22816 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 590 592
use scs8hd_buf_2  _213_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _085_
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_38
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_111
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_134
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_138
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_153
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_168
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_180
timestamp 1586364061
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 22816 0 1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 130 592
use scs8hd_inv_8  _109_
timestamp 1586364061
transform 1 0 1656 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 1050 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_25
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_49
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_44
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_54
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _112_
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_27_58
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_74
timestamp 1586364061
transform 1 0 7912 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_71
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _094_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_27_100
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_124
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_6  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_130
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_127
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_137
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 590 592
use scs8hd_inv_8  _087_
timestamp 1586364061
transform 1 0 14444 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_157
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_154
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_166
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_169
timestamp 1586364061
transform 1 0 16652 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_178
timestamp 1586364061
transform 1 0 17480 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_181
timestamp 1586364061
transform 1 0 17756 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_193
timestamp 1586364061
transform 1 0 18860 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_182
timestamp 1586364061
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_205
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 22816 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 22816 0 1 16864
box -38 -48 314 592
use scs8hd_decap_6  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_8
timestamp 1586364061
transform 1 0 1840 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_20
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_28_26
timestamp 1586364061
transform 1 0 3496 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_41
timestamp 1586364061
transform 1 0 4876 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_28_53
timestamp 1586364061
transform 1 0 5980 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_65
timestamp 1586364061
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_81
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_85
timestamp 1586364061
transform 1 0 8924 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_91
timestamp 1586364061
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_8  _088_
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_6  FILLER_28_114
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_120
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 130 592
use scs8hd_conb_1  _192_
timestamp 1586364061
transform 1 0 13800 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_130
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 22816 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3312 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_19
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_33
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_37
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_44
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_48
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_102
timestamp 1586364061
transform 1 0 10488 0 1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_148
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_160
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_172
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_180
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_214
timestamp 1586364061
transform 1 0 20792 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 22816 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_229
timestamp 1586364061
transform 1 0 22172 0 1 17952
box -38 -48 406 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 2300 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_11
timestamp 1586364061
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_8  _110_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_53
timestamp 1586364061
transform 1 0 5980 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_conb_1  _195_
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_91
timestamp 1586364061
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_119
timestamp 1586364061
transform 1 0 12052 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_1  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_135
timestamp 1586364061
transform 1 0 13524 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_147
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_218
timestamp 1586364061
transform 1 0 21160 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_230
timestamp 1586364061
transform 1 0 22264 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 2300 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_18
timestamp 1586364061
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_22
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_31_34
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_38
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 130 592
use scs8hd_conb_1  _186_
timestamp 1586364061
transform 1 0 5704 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 5520 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_42
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_46
timestamp 1586364061
transform 1 0 5336 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_31_83
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 130 592
use scs8hd_inv_8  _093_
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 406 592
use scs8hd_inv_8  _100_
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_126
timestamp 1586364061
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_130
timestamp 1586364061
transform 1 0 13064 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_134
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_146
timestamp 1586364061
transform 1 0 14536 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_158
timestamp 1586364061
transform 1 0 15640 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_170
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_182
timestamp 1586364061
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_188
timestamp 1586364061
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_192
timestamp 1586364061
transform 1 0 18768 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 22816 0 1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 130 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_7
timestamp 1586364061
transform 1 0 1748 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_30
timestamp 1586364061
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_8  _111_
timestamp 1586364061
transform 1 0 5980 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_52
timestamp 1586364061
transform 1 0 5888 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_62
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_74
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_86
timestamp 1586364061
transform 1 0 9016 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_32_96
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10856 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_100
timestamp 1586364061
transform 1 0 10304 0 -1 20128
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_115
timestamp 1586364061
transform 1 0 11684 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_132
timestamp 1586364061
transform 1 0 13248 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_144
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17940 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_182
timestamp 1586364061
transform 1 0 17848 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_186
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_198
timestamp 1586364061
transform 1 0 19320 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_210
timestamp 1586364061
transform 1 0 20424 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 22816 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_6
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_10
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_22
timestamp 1586364061
transform 1 0 3128 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_30
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_35
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_47
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_52
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_56
timestamp 1586364061
transform 1 0 6256 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_60
timestamp 1586364061
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_65
timestamp 1586364061
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_69
timestamp 1586364061
transform 1 0 7452 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 8740 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_87
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_91
timestamp 1586364061
transform 1 0 9476 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_95
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_104
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_108
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_99
timestamp 1586364061
transform 1 0 10212 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_120
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_111
timestamp 1586364061
transform 1 0 11316 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_123
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_131
timestamp 1586364061
transform 1 0 13156 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_137
timestamp 1586364061
transform 1 0 13708 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_135
timestamp 1586364061
transform 1 0 13524 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _212_
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__212__A
timestamp 1586364061
transform 1 0 15088 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_141
timestamp 1586364061
transform 1 0 14076 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_145
timestamp 1586364061
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_150
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_147
timestamp 1586364061
transform 1 0 14628 0 -1 21216
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_154
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_169
timestamp 1586364061
transform 1 0 16652 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_173
timestamp 1586364061
transform 1 0 17020 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_181
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_187
timestamp 1586364061
transform 1 0 18308 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_191
timestamp 1586364061
transform 1 0 18676 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_203
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_218
timestamp 1586364061
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 22816 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 22816 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_33_222
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_33_230
timestamp 1586364061
transform 1 0 22264 0 1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 22816 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 314 592
<< labels >>
rlabel metal3 s 23520 1096 24000 1216 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 552 480 672 6 address[1]
port 1 nsew default input
rlabel metal3 s 23520 3408 24000 3528 6 address[2]
port 2 nsew default input
rlabel metal2 s 3422 0 3478 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 846 23520 902 24000 6 address[4]
port 4 nsew default input
rlabel metal3 s 0 1640 480 1760 6 address[5]
port 5 nsew default input
rlabel metal2 s 4250 23520 4306 24000 6 bottom_left_grid_pin_11_
port 6 nsew default input
rlabel metal2 s 7654 0 7710 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 9126 0 9182 480 6 bottom_left_grid_pin_15_
port 8 nsew default input
rlabel metal3 s 0 2728 480 2848 6 bottom_left_grid_pin_1_
port 9 nsew default input
rlabel metal2 s 4894 0 4950 480 6 bottom_left_grid_pin_3_
port 10 nsew default input
rlabel metal2 s 2502 23520 2558 24000 6 bottom_left_grid_pin_5_
port 11 nsew default input
rlabel metal2 s 6274 0 6330 480 6 bottom_left_grid_pin_7_
port 12 nsew default input
rlabel metal3 s 23520 5856 24000 5976 6 bottom_left_grid_pin_9_
port 13 nsew default input
rlabel metal3 s 0 3952 480 4072 6 bottom_right_grid_pin_11_
port 14 nsew default input
rlabel metal3 s 23520 8168 24000 8288 6 chanx_right_in[0]
port 15 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_right_in[1]
port 16 nsew default input
rlabel metal2 s 5906 23520 5962 24000 6 chanx_right_in[2]
port 17 nsew default input
rlabel metal2 s 7654 23520 7710 24000 6 chanx_right_in[3]
port 18 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chanx_right_in[4]
port 19 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_right_in[5]
port 20 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chanx_right_in[6]
port 21 nsew default input
rlabel metal3 s 0 7352 480 7472 6 chanx_right_in[7]
port 22 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_right_in[8]
port 23 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_right_out[0]
port 24 nsew default tristate
rlabel metal2 s 13358 0 13414 480 6 chanx_right_out[1]
port 25 nsew default tristate
rlabel metal3 s 23520 10616 24000 10736 6 chanx_right_out[2]
port 26 nsew default tristate
rlabel metal2 s 14738 0 14794 480 6 chanx_right_out[3]
port 27 nsew default tristate
rlabel metal2 s 9402 23520 9458 24000 6 chanx_right_out[4]
port 28 nsew default tristate
rlabel metal3 s 23520 13064 24000 13184 6 chanx_right_out[5]
port 29 nsew default tristate
rlabel metal3 s 0 10752 480 10872 6 chanx_right_out[6]
port 30 nsew default tristate
rlabel metal2 s 16118 0 16174 480 6 chanx_right_out[7]
port 31 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 chanx_right_out[8]
port 32 nsew default tristate
rlabel metal2 s 11058 23520 11114 24000 6 chany_bottom_in[0]
port 33 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chany_bottom_in[1]
port 34 nsew default input
rlabel metal2 s 17590 0 17646 480 6 chany_bottom_in[2]
port 35 nsew default input
rlabel metal3 s 0 14152 480 14272 6 chany_bottom_in[3]
port 36 nsew default input
rlabel metal2 s 18970 0 19026 480 6 chany_bottom_in[4]
port 37 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chany_bottom_in[5]
port 38 nsew default input
rlabel metal2 s 12806 23520 12862 24000 6 chany_bottom_in[6]
port 39 nsew default input
rlabel metal3 s 0 16464 480 16584 6 chany_bottom_in[7]
port 40 nsew default input
rlabel metal2 s 14554 23520 14610 24000 6 chany_bottom_in[8]
port 41 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chany_bottom_out[0]
port 42 nsew default tristate
rlabel metal2 s 16210 23520 16266 24000 6 chany_bottom_out[1]
port 43 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 chany_bottom_out[2]
port 44 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chany_bottom_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 19864 480 19984 6 chany_bottom_out[4]
port 46 nsew default tristate
rlabel metal3 s 23520 15376 24000 15496 6 chany_bottom_out[5]
port 47 nsew default tristate
rlabel metal2 s 21822 0 21878 480 6 chany_bottom_out[6]
port 48 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 chany_bottom_out[7]
port 49 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_bottom_out[8]
port 50 nsew default tristate
rlabel metal2 s 2042 0 2098 480 6 data_in
port 51 nsew default input
rlabel metal2 s 662 0 718 480 6 enable
port 52 nsew default input
rlabel metal3 s 23520 17824 24000 17944 6 right_bottom_grid_pin_12_
port 53 nsew default input
rlabel metal2 s 23110 23520 23166 24000 6 right_top_grid_pin_11_
port 54 nsew default input
rlabel metal3 s 23520 22584 24000 22704 6 right_top_grid_pin_13_
port 55 nsew default input
rlabel metal3 s 0 23264 480 23384 6 right_top_grid_pin_15_
port 56 nsew default input
rlabel metal2 s 17958 23520 18014 24000 6 right_top_grid_pin_1_
port 57 nsew default input
rlabel metal2 s 19706 23520 19762 24000 6 right_top_grid_pin_3_
port 58 nsew default input
rlabel metal3 s 0 22176 480 22296 6 right_top_grid_pin_5_
port 59 nsew default input
rlabel metal2 s 21362 23520 21418 24000 6 right_top_grid_pin_7_
port 60 nsew default input
rlabel metal3 s 23520 20136 24000 20256 6 right_top_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 4944 2128 5264 21808 6 vpwr
port 62 nsew default input
rlabel metal4 s 8944 2128 9264 21808 6 vgnd
port 63 nsew default input
<< end >>
