magic
tech sky130A
magscale 1 2
timestamp 1605198272
<< locali >>
rect 10977 7259 11011 7497
rect 16589 2295 16623 2397
<< viali >>
rect 19073 20553 19107 20587
rect 18889 20349 18923 20383
rect 19993 20349 20027 20383
rect 20177 20213 20211 20247
rect 4261 20009 4295 20043
rect 18797 20009 18831 20043
rect 4077 19873 4111 19907
rect 18613 19873 18647 19907
rect 19717 19873 19751 19907
rect 17785 19805 17819 19839
rect 19901 19737 19935 19771
rect 4537 19669 4571 19703
rect 12449 19261 12483 19295
rect 14013 19261 14047 19295
rect 18797 19261 18831 19295
rect 19901 19261 19935 19295
rect 12725 19193 12759 19227
rect 14280 19193 14314 19227
rect 20177 19193 20211 19227
rect 15393 19125 15427 19159
rect 18981 19125 19015 19159
rect 14105 18853 14139 18887
rect 19809 18853 19843 18887
rect 10333 18785 10367 18819
rect 13829 18785 13863 18819
rect 19533 18785 19567 18819
rect 10609 18717 10643 18751
rect 13461 18377 13495 18411
rect 19625 18377 19659 18411
rect 20729 18377 20763 18411
rect 10425 18173 10459 18207
rect 13277 18173 13311 18207
rect 19441 18173 19475 18207
rect 20545 18173 20579 18207
rect 10701 18105 10735 18139
rect 19717 17697 19751 17731
rect 19901 17493 19935 17527
rect 18981 17289 19015 17323
rect 12817 17153 12851 17187
rect 20177 17153 20211 17187
rect 12541 17085 12575 17119
rect 18797 17085 18831 17119
rect 19901 17085 19935 17119
rect 18613 16745 18647 16779
rect 13001 16677 13035 16711
rect 19809 16677 19843 16711
rect 12725 16609 12759 16643
rect 18429 16609 18463 16643
rect 19533 16609 19567 16643
rect 18521 16201 18555 16235
rect 18337 15997 18371 16031
rect 19441 15997 19475 16031
rect 20545 15997 20579 16031
rect 19625 15861 19659 15895
rect 20729 15861 20763 15895
rect 18797 15657 18831 15691
rect 10793 15589 10827 15623
rect 10517 15521 10551 15555
rect 18613 15521 18647 15555
rect 19717 15521 19751 15555
rect 19901 15317 19935 15351
rect 19073 15113 19107 15147
rect 7757 14909 7791 14943
rect 9045 14909 9079 14943
rect 9321 14909 9355 14943
rect 18889 14909 18923 14943
rect 19993 14909 20027 14943
rect 8033 14841 8067 14875
rect 20269 14841 20303 14875
rect 16957 14773 16991 14807
rect 8309 14501 8343 14535
rect 19809 14501 19843 14535
rect 8033 14433 8067 14467
rect 17325 14433 17359 14467
rect 18429 14433 18463 14467
rect 19533 14433 19567 14467
rect 12541 14365 12575 14399
rect 15301 14365 15335 14399
rect 16313 14365 16347 14399
rect 17509 14229 17543 14263
rect 18613 14229 18647 14263
rect 12449 14025 12483 14059
rect 15577 14025 15611 14059
rect 13001 13889 13035 13923
rect 16221 13889 16255 13923
rect 18705 13889 18739 13923
rect 19993 13889 20027 13923
rect 12817 13821 12851 13855
rect 16037 13821 16071 13855
rect 18521 13821 18555 13855
rect 19809 13821 19843 13855
rect 12909 13685 12943 13719
rect 14565 13685 14599 13719
rect 15945 13685 15979 13719
rect 12725 13481 12759 13515
rect 14197 13481 14231 13515
rect 17969 13481 18003 13515
rect 19257 13481 19291 13515
rect 11612 13345 11646 13379
rect 15301 13345 15335 13379
rect 15557 13345 15591 13379
rect 19625 13345 19659 13379
rect 11345 13277 11379 13311
rect 18061 13277 18095 13311
rect 18153 13277 18187 13311
rect 19717 13277 19751 13311
rect 19809 13277 19843 13311
rect 17601 13209 17635 13243
rect 16681 13141 16715 13175
rect 15485 12937 15519 12971
rect 10149 12801 10183 12835
rect 15761 12801 15795 12835
rect 20545 12801 20579 12835
rect 12817 12733 12851 12767
rect 15669 12733 15703 12767
rect 16028 12733 16062 12767
rect 18061 12733 18095 12767
rect 20269 12733 20303 12767
rect 10416 12665 10450 12699
rect 13062 12665 13096 12699
rect 18306 12665 18340 12699
rect 11529 12597 11563 12631
rect 14197 12597 14231 12631
rect 17141 12597 17175 12631
rect 19441 12597 19475 12631
rect 9873 12393 9907 12427
rect 11437 12393 11471 12427
rect 15853 12393 15887 12427
rect 18153 12393 18187 12427
rect 11897 12325 11931 12359
rect 8585 12257 8619 12291
rect 10241 12257 10275 12291
rect 11805 12257 11839 12291
rect 13001 12257 13035 12291
rect 13268 12257 13302 12291
rect 15669 12257 15703 12291
rect 16773 12257 16807 12291
rect 17040 12257 17074 12291
rect 19625 12257 19659 12291
rect 19717 12257 19751 12291
rect 10333 12189 10367 12223
rect 10517 12189 10551 12223
rect 11989 12189 12023 12223
rect 19901 12189 19935 12223
rect 14381 12053 14415 12087
rect 19257 12053 19291 12087
rect 10609 11849 10643 11883
rect 13093 11849 13127 11883
rect 14657 11849 14691 11883
rect 16221 11849 16255 11883
rect 13737 11713 13771 11747
rect 15117 11713 15151 11747
rect 15301 11713 15335 11747
rect 16773 11713 16807 11747
rect 18061 11713 18095 11747
rect 19533 11713 19567 11747
rect 19717 11713 19751 11747
rect 9229 11645 9263 11679
rect 15025 11645 15059 11679
rect 16589 11645 16623 11679
rect 9496 11577 9530 11611
rect 19441 11577 19475 11611
rect 20637 11577 20671 11611
rect 13461 11509 13495 11543
rect 13553 11509 13587 11543
rect 16681 11509 16715 11543
rect 19073 11509 19107 11543
rect 9781 11305 9815 11339
rect 15301 11305 15335 11339
rect 16129 11305 16163 11339
rect 16773 11305 16807 11339
rect 19809 11305 19843 11339
rect 13093 11237 13127 11271
rect 16589 11237 16623 11271
rect 17141 11237 17175 11271
rect 10149 11169 10183 11203
rect 10241 11169 10275 11203
rect 11981 11169 12015 11203
rect 14657 11169 14691 11203
rect 16313 11169 16347 11203
rect 17233 11169 17267 11203
rect 18685 11169 18719 11203
rect 10333 11101 10367 11135
rect 17325 11101 17359 11135
rect 18429 11101 18463 11135
rect 11805 11033 11839 11067
rect 9873 10761 9907 10795
rect 10793 10761 10827 10795
rect 13829 10761 13863 10795
rect 15485 10761 15519 10795
rect 16405 10761 16439 10795
rect 20821 10761 20855 10795
rect 11437 10625 11471 10659
rect 14105 10625 14139 10659
rect 17049 10625 17083 10659
rect 19441 10625 19475 10659
rect 8493 10557 8527 10591
rect 12449 10557 12483 10591
rect 14361 10557 14395 10591
rect 18337 10557 18371 10591
rect 8760 10489 8794 10523
rect 11161 10489 11195 10523
rect 12694 10489 12728 10523
rect 16773 10489 16807 10523
rect 19708 10489 19742 10523
rect 11253 10421 11287 10455
rect 16865 10421 16899 10455
rect 18521 10421 18555 10455
rect 8033 10217 8067 10251
rect 9689 10217 9723 10251
rect 13093 10217 13127 10251
rect 14013 10217 14047 10251
rect 14105 10217 14139 10251
rect 18981 10217 19015 10251
rect 10057 10149 10091 10183
rect 11520 10149 11554 10183
rect 16580 10149 16614 10183
rect 7021 10081 7055 10115
rect 8401 10081 8435 10115
rect 10149 10081 10183 10115
rect 13185 10081 13219 10115
rect 16313 10081 16347 10115
rect 18889 10081 18923 10115
rect 8493 10013 8527 10047
rect 8677 10013 8711 10047
rect 10333 10013 10367 10047
rect 11253 10013 11287 10047
rect 13277 10013 13311 10047
rect 14197 10013 14231 10047
rect 15301 10013 15335 10047
rect 19073 10013 19107 10047
rect 12633 9945 12667 9979
rect 12725 9877 12759 9911
rect 13645 9877 13679 9911
rect 17693 9877 17727 9911
rect 18521 9877 18555 9911
rect 8953 9673 8987 9707
rect 11529 9673 11563 9707
rect 20821 9673 20855 9707
rect 9873 9605 9907 9639
rect 10149 9537 10183 9571
rect 12449 9537 12483 9571
rect 7573 9469 7607 9503
rect 10057 9469 10091 9503
rect 13553 9469 13587 9503
rect 13820 9469 13854 9503
rect 15761 9469 15795 9503
rect 16028 9469 16062 9503
rect 18337 9469 18371 9503
rect 19441 9469 19475 9503
rect 19708 9469 19742 9503
rect 7840 9401 7874 9435
rect 10416 9401 10450 9435
rect 14933 9333 14967 9367
rect 17141 9333 17175 9367
rect 18521 9333 18555 9367
rect 8033 9129 8067 9163
rect 9781 9129 9815 9163
rect 11345 9129 11379 9163
rect 13645 9129 13679 9163
rect 14105 9129 14139 9163
rect 19257 9129 19291 9163
rect 14013 9061 14047 9095
rect 16856 9061 16890 9095
rect 8401 8993 8435 9027
rect 8493 8993 8527 9027
rect 10149 8993 10183 9027
rect 11713 8993 11747 9027
rect 11805 8993 11839 9027
rect 15301 8993 15335 9027
rect 19165 8993 19199 9027
rect 7021 8925 7055 8959
rect 8585 8925 8619 8959
rect 10241 8925 10275 8959
rect 10425 8925 10459 8959
rect 11897 8925 11931 8959
rect 14289 8925 14323 8959
rect 15485 8925 15519 8959
rect 16589 8925 16623 8959
rect 19349 8925 19383 8959
rect 17969 8857 18003 8891
rect 18797 8789 18831 8823
rect 8401 8585 8435 8619
rect 11253 8585 11287 8619
rect 12633 8585 12667 8619
rect 14933 8585 14967 8619
rect 16129 8585 16163 8619
rect 18245 8585 18279 8619
rect 9873 8449 9907 8483
rect 13553 8449 13587 8483
rect 16773 8449 16807 8483
rect 19165 8449 19199 8483
rect 7021 8381 7055 8415
rect 12449 8381 12483 8415
rect 13820 8381 13854 8415
rect 15945 8381 15979 8415
rect 16497 8381 16531 8415
rect 16589 8381 16623 8415
rect 18061 8381 18095 8415
rect 7288 8313 7322 8347
rect 10140 8313 10174 8347
rect 19410 8313 19444 8347
rect 15761 8245 15795 8279
rect 20545 8245 20579 8279
rect 8033 8041 8067 8075
rect 11069 8041 11103 8075
rect 16681 8041 16715 8075
rect 16773 8041 16807 8075
rect 5641 7973 5675 8007
rect 12142 7973 12176 8007
rect 18144 7973 18178 8007
rect 6653 7905 6687 7939
rect 6920 7905 6954 7939
rect 9689 7905 9723 7939
rect 9956 7905 9990 7939
rect 14105 7905 14139 7939
rect 11897 7837 11931 7871
rect 15301 7837 15335 7871
rect 16957 7837 16991 7871
rect 17877 7837 17911 7871
rect 13277 7701 13311 7735
rect 14289 7701 14323 7735
rect 16313 7701 16347 7735
rect 19257 7701 19291 7735
rect 7113 7497 7147 7531
rect 9413 7497 9447 7531
rect 10977 7497 11011 7531
rect 7757 7361 7791 7395
rect 10057 7361 10091 7395
rect 7481 7293 7515 7327
rect 16405 7429 16439 7463
rect 20821 7429 20855 7463
rect 13093 7361 13127 7395
rect 14013 7361 14047 7395
rect 17049 7361 17083 7395
rect 19441 7361 19475 7395
rect 11069 7293 11103 7327
rect 12909 7293 12943 7327
rect 18061 7293 18095 7327
rect 19708 7293 19742 7327
rect 10977 7225 11011 7259
rect 11345 7225 11379 7259
rect 14280 7225 14314 7259
rect 16865 7225 16899 7259
rect 18337 7225 18371 7259
rect 7573 7157 7607 7191
rect 9781 7157 9815 7191
rect 9873 7157 9907 7191
rect 12449 7157 12483 7191
rect 12817 7157 12851 7191
rect 15393 7157 15427 7191
rect 16773 7157 16807 7191
rect 7297 6953 7331 6987
rect 12081 6953 12115 6987
rect 12541 6953 12575 6987
rect 15669 6953 15703 6987
rect 16865 6953 16899 6987
rect 17233 6953 17267 6987
rect 18797 6953 18831 6987
rect 7665 6885 7699 6919
rect 12449 6885 12483 6919
rect 14013 6885 14047 6919
rect 15761 6885 15795 6919
rect 10057 6817 10091 6851
rect 11989 6817 12023 6851
rect 14105 6817 14139 6851
rect 17325 6817 17359 6851
rect 18889 6817 18923 6851
rect 7757 6749 7791 6783
rect 7849 6749 7883 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 12725 6749 12759 6783
rect 14289 6749 14323 6783
rect 15853 6749 15887 6783
rect 17417 6749 17451 6783
rect 19073 6749 19107 6783
rect 9689 6681 9723 6715
rect 13645 6681 13679 6715
rect 11805 6613 11839 6647
rect 15301 6613 15335 6647
rect 18429 6613 18463 6647
rect 8217 6409 8251 6443
rect 10425 6409 10459 6443
rect 13829 6409 13863 6443
rect 17141 6409 17175 6443
rect 11437 6341 11471 6375
rect 5733 6273 5767 6307
rect 6837 6273 6871 6307
rect 15761 6273 15795 6307
rect 9045 6205 9079 6239
rect 11253 6205 11287 6239
rect 12449 6205 12483 6239
rect 12716 6205 12750 6239
rect 14657 6205 14691 6239
rect 16028 6205 16062 6239
rect 18061 6205 18095 6239
rect 18317 6205 18351 6239
rect 20545 6205 20579 6239
rect 7104 6137 7138 6171
rect 9312 6137 9346 6171
rect 14841 6069 14875 6103
rect 19441 6069 19475 6103
rect 20729 6069 20763 6103
rect 7205 5865 7239 5899
rect 14013 5865 14047 5899
rect 15301 5865 15335 5899
rect 15669 5865 15703 5899
rect 6193 5797 6227 5831
rect 7573 5729 7607 5763
rect 9689 5729 9723 5763
rect 10793 5729 10827 5763
rect 11060 5729 11094 5763
rect 15761 5729 15795 5763
rect 16865 5729 16899 5763
rect 18420 5729 18454 5763
rect 5181 5661 5215 5695
rect 7665 5661 7699 5695
rect 7757 5661 7791 5695
rect 14105 5661 14139 5695
rect 14289 5661 14323 5695
rect 15853 5661 15887 5695
rect 17049 5661 17083 5695
rect 18153 5661 18187 5695
rect 9873 5525 9907 5559
rect 12173 5525 12207 5559
rect 13645 5525 13679 5559
rect 19533 5525 19567 5559
rect 8217 5321 8251 5355
rect 10609 5321 10643 5355
rect 12449 5321 12483 5355
rect 15301 5321 15335 5355
rect 17049 5253 17083 5287
rect 18061 5253 18095 5287
rect 6837 5185 6871 5219
rect 9229 5185 9263 5219
rect 13093 5185 13127 5219
rect 15761 5185 15795 5219
rect 15945 5185 15979 5219
rect 18705 5185 18739 5219
rect 20085 5185 20119 5219
rect 20177 5185 20211 5219
rect 12817 5117 12851 5151
rect 14197 5117 14231 5151
rect 15669 5117 15703 5151
rect 16865 5117 16899 5151
rect 18429 5117 18463 5151
rect 5733 5049 5767 5083
rect 7104 5049 7138 5083
rect 9496 5049 9530 5083
rect 12909 5049 12943 5083
rect 18521 5049 18555 5083
rect 14381 4981 14415 5015
rect 19625 4981 19659 5015
rect 19993 4981 20027 5015
rect 7665 4777 7699 4811
rect 8125 4777 8159 4811
rect 9689 4777 9723 4811
rect 11713 4777 11747 4811
rect 11805 4777 11839 4811
rect 6561 4641 6595 4675
rect 8033 4641 8067 4675
rect 10057 4641 10091 4675
rect 12909 4641 12943 4675
rect 13176 4641 13210 4675
rect 15301 4641 15335 4675
rect 15568 4641 15602 4675
rect 17877 4641 17911 4675
rect 19625 4641 19659 4675
rect 8217 4573 8251 4607
rect 10149 4573 10183 4607
rect 10333 4573 10367 4607
rect 11989 4573 12023 4607
rect 17969 4573 18003 4607
rect 18061 4573 18095 4607
rect 19717 4573 19751 4607
rect 19809 4573 19843 4607
rect 6745 4437 6779 4471
rect 11345 4437 11379 4471
rect 14289 4437 14323 4471
rect 16681 4437 16715 4471
rect 17509 4437 17543 4471
rect 19257 4437 19291 4471
rect 8217 4233 8251 4267
rect 16497 4233 16531 4267
rect 6837 4097 6871 4131
rect 9873 4097 9907 4131
rect 14197 4097 14231 4131
rect 10140 4029 10174 4063
rect 12449 4029 12483 4063
rect 13921 4029 13955 4063
rect 14013 4029 14047 4063
rect 15117 4029 15151 4063
rect 19073 4029 19107 4063
rect 7104 3961 7138 3995
rect 15384 3961 15418 3995
rect 19340 3961 19374 3995
rect 5733 3893 5767 3927
rect 11253 3893 11287 3927
rect 12633 3893 12667 3927
rect 13553 3893 13587 3927
rect 18061 3893 18095 3927
rect 20453 3893 20487 3927
rect 7113 3689 7147 3723
rect 8033 3689 8067 3723
rect 8493 3689 8527 3723
rect 15669 3689 15703 3723
rect 16129 3689 16163 3723
rect 10876 3621 10910 3655
rect 19717 3621 19751 3655
rect 5825 3553 5859 3587
rect 6929 3553 6963 3587
rect 8401 3553 8435 3587
rect 13084 3553 13118 3587
rect 16037 3553 16071 3587
rect 17489 3553 17523 3587
rect 19441 3553 19475 3587
rect 8677 3485 8711 3519
rect 10609 3485 10643 3519
rect 12817 3485 12851 3519
rect 16313 3485 16347 3519
rect 17233 3485 17267 3519
rect 4997 3417 5031 3451
rect 6009 3417 6043 3451
rect 11989 3349 12023 3383
rect 14197 3349 14231 3383
rect 18613 3349 18647 3383
rect 7021 3145 7055 3179
rect 9321 3145 9355 3179
rect 10793 3145 10827 3179
rect 15669 3145 15703 3179
rect 18061 3145 18095 3179
rect 19625 3145 19659 3179
rect 7941 3009 7975 3043
rect 11345 3009 11379 3043
rect 13093 3009 13127 3043
rect 14657 3009 14691 3043
rect 16129 3009 16163 3043
rect 16313 3009 16347 3043
rect 18613 3009 18647 3043
rect 20085 3009 20119 3043
rect 20177 3009 20211 3043
rect 5641 2941 5675 2975
rect 6862 2941 6896 2975
rect 18429 2941 18463 2975
rect 4629 2873 4663 2907
rect 8208 2873 8242 2907
rect 12909 2873 12943 2907
rect 14565 2873 14599 2907
rect 16037 2873 16071 2907
rect 18521 2873 18555 2907
rect 19993 2873 20027 2907
rect 5825 2805 5859 2839
rect 11161 2805 11195 2839
rect 11253 2805 11287 2839
rect 12541 2805 12575 2839
rect 13001 2805 13035 2839
rect 14105 2805 14139 2839
rect 14473 2805 14507 2839
rect 8125 2601 8159 2635
rect 10241 2601 10275 2635
rect 13093 2601 13127 2635
rect 16681 2601 16715 2635
rect 8585 2533 8619 2567
rect 7021 2465 7055 2499
rect 8493 2465 8527 2499
rect 11437 2465 11471 2499
rect 13461 2465 13495 2499
rect 13553 2465 13587 2499
rect 15485 2465 15519 2499
rect 17049 2465 17083 2499
rect 19441 2465 19475 2499
rect 5825 2397 5859 2431
rect 8677 2397 8711 2431
rect 10333 2397 10367 2431
rect 10517 2397 10551 2431
rect 13737 2397 13771 2431
rect 16589 2397 16623 2431
rect 17141 2397 17175 2431
rect 17325 2397 17359 2431
rect 19533 2397 19567 2431
rect 19717 2397 19751 2431
rect 9873 2329 9907 2363
rect 7205 2261 7239 2295
rect 11621 2261 11655 2295
rect 15669 2261 15703 2295
rect 16589 2261 16623 2295
rect 19073 2261 19107 2295
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 19058 20584 19064 20596
rect 19019 20556 19064 20584
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 18877 20383 18935 20389
rect 18877 20349 18889 20383
rect 18923 20380 18935 20383
rect 19794 20380 19800 20392
rect 18923 20352 19800 20380
rect 18923 20349 18935 20352
rect 18877 20343 18935 20349
rect 19794 20340 19800 20352
rect 19852 20340 19858 20392
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20349 20039 20383
rect 19981 20343 20039 20349
rect 17954 20272 17960 20324
rect 18012 20312 18018 20324
rect 19996 20312 20024 20343
rect 18012 20284 20024 20312
rect 18012 20272 18018 20284
rect 20162 20244 20168 20256
rect 20123 20216 20168 20244
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 2866 20000 2872 20052
rect 2924 20040 2930 20052
rect 4249 20043 4307 20049
rect 4249 20040 4261 20043
rect 2924 20012 4261 20040
rect 2924 20000 2930 20012
rect 4249 20009 4261 20012
rect 4295 20009 4307 20043
rect 18782 20040 18788 20052
rect 18743 20012 18788 20040
rect 4249 20003 4307 20009
rect 18782 20000 18788 20012
rect 18840 20000 18846 20052
rect 15838 19932 15844 19984
rect 15896 19972 15902 19984
rect 15896 19944 19748 19972
rect 15896 19932 15902 19944
rect 4065 19907 4123 19913
rect 4065 19873 4077 19907
rect 4111 19904 4123 19907
rect 18598 19904 18604 19916
rect 4111 19876 4568 19904
rect 18559 19876 18604 19904
rect 4111 19873 4123 19876
rect 4065 19867 4123 19873
rect 4540 19709 4568 19876
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 19720 19913 19748 19944
rect 19705 19907 19763 19913
rect 19705 19873 19717 19907
rect 19751 19873 19763 19907
rect 19705 19867 19763 19873
rect 17773 19839 17831 19845
rect 17773 19805 17785 19839
rect 17819 19836 17831 19839
rect 20070 19836 20076 19848
rect 17819 19808 20076 19836
rect 17819 19805 17831 19808
rect 17773 19799 17831 19805
rect 20070 19796 20076 19808
rect 20128 19796 20134 19848
rect 19886 19768 19892 19780
rect 19847 19740 19892 19768
rect 19886 19728 19892 19740
rect 19944 19728 19950 19780
rect 4525 19703 4583 19709
rect 4525 19669 4537 19703
rect 4571 19700 4583 19703
rect 4798 19700 4804 19712
rect 4571 19672 4804 19700
rect 4571 19669 4583 19672
rect 4525 19663 4583 19669
rect 4798 19660 4804 19672
rect 4856 19660 4862 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 4798 19456 4804 19508
rect 4856 19496 4862 19508
rect 20714 19496 20720 19508
rect 4856 19468 20720 19496
rect 4856 19456 4862 19468
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 10836 19264 12449 19292
rect 10836 19252 10842 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 13998 19292 14004 19304
rect 13959 19264 14004 19292
rect 12437 19255 12495 19261
rect 13998 19252 14004 19264
rect 14056 19252 14062 19304
rect 17954 19292 17960 19304
rect 14200 19264 17960 19292
rect 12713 19227 12771 19233
rect 12713 19193 12725 19227
rect 12759 19224 12771 19227
rect 14200 19224 14228 19264
rect 17954 19252 17960 19264
rect 18012 19252 18018 19304
rect 18785 19295 18843 19301
rect 18785 19261 18797 19295
rect 18831 19261 18843 19295
rect 18785 19255 18843 19261
rect 12759 19196 14228 19224
rect 14268 19227 14326 19233
rect 12759 19193 12771 19196
rect 12713 19187 12771 19193
rect 14268 19193 14280 19227
rect 14314 19224 14326 19227
rect 14366 19224 14372 19236
rect 14314 19196 14372 19224
rect 14314 19193 14326 19196
rect 14268 19187 14326 19193
rect 14366 19184 14372 19196
rect 14424 19184 14430 19236
rect 18800 19224 18828 19255
rect 19150 19252 19156 19304
rect 19208 19292 19214 19304
rect 19889 19295 19947 19301
rect 19889 19292 19901 19295
rect 19208 19264 19901 19292
rect 19208 19252 19214 19264
rect 19889 19261 19901 19264
rect 19935 19261 19947 19295
rect 19889 19255 19947 19261
rect 20165 19227 20223 19233
rect 20165 19224 20177 19227
rect 18800 19196 20177 19224
rect 20165 19193 20177 19196
rect 20211 19193 20223 19227
rect 20165 19187 20223 19193
rect 14182 19116 14188 19168
rect 14240 19156 14246 19168
rect 15381 19159 15439 19165
rect 15381 19156 15393 19159
rect 14240 19128 15393 19156
rect 14240 19116 14246 19128
rect 15381 19125 15393 19128
rect 15427 19125 15439 19159
rect 18966 19156 18972 19168
rect 18927 19128 18972 19156
rect 15381 19119 15439 19125
rect 18966 19116 18972 19128
rect 19024 19116 19030 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 13998 18912 14004 18964
rect 14056 18952 14062 18964
rect 15194 18952 15200 18964
rect 14056 18924 15200 18952
rect 14056 18912 14062 18924
rect 15194 18912 15200 18924
rect 15252 18912 15258 18964
rect 14093 18887 14151 18893
rect 14093 18853 14105 18887
rect 14139 18884 14151 18887
rect 18598 18884 18604 18896
rect 14139 18856 18604 18884
rect 14139 18853 14151 18856
rect 14093 18847 14151 18853
rect 18598 18844 18604 18856
rect 18656 18844 18662 18896
rect 19794 18884 19800 18896
rect 19755 18856 19800 18884
rect 19794 18844 19800 18856
rect 19852 18844 19858 18896
rect 9766 18776 9772 18828
rect 9824 18816 9830 18828
rect 10321 18819 10379 18825
rect 10321 18816 10333 18819
rect 9824 18788 10333 18816
rect 9824 18776 9830 18788
rect 10321 18785 10333 18788
rect 10367 18785 10379 18819
rect 10321 18779 10379 18785
rect 13817 18819 13875 18825
rect 13817 18785 13829 18819
rect 13863 18816 13875 18819
rect 13906 18816 13912 18828
rect 13863 18788 13912 18816
rect 13863 18785 13875 18788
rect 13817 18779 13875 18785
rect 13906 18776 13912 18788
rect 13964 18776 13970 18828
rect 16574 18776 16580 18828
rect 16632 18816 16638 18828
rect 19521 18819 19579 18825
rect 19521 18816 19533 18819
rect 16632 18788 19533 18816
rect 16632 18776 16638 18788
rect 19521 18785 19533 18788
rect 19567 18785 19579 18819
rect 19521 18779 19579 18785
rect 10597 18751 10655 18757
rect 10597 18717 10609 18751
rect 10643 18748 10655 18751
rect 15838 18748 15844 18760
rect 10643 18720 15844 18748
rect 10643 18717 10655 18720
rect 10597 18711 10655 18717
rect 15838 18708 15844 18720
rect 15896 18708 15902 18760
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 13449 18411 13507 18417
rect 13449 18377 13461 18411
rect 13495 18408 13507 18411
rect 17954 18408 17960 18420
rect 13495 18380 17960 18408
rect 13495 18377 13507 18380
rect 13449 18371 13507 18377
rect 17954 18368 17960 18380
rect 18012 18368 18018 18420
rect 19610 18408 19616 18420
rect 19571 18380 19616 18408
rect 19610 18368 19616 18380
rect 19668 18368 19674 18420
rect 20714 18408 20720 18420
rect 20675 18380 20720 18408
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 9950 18164 9956 18216
rect 10008 18204 10014 18216
rect 10413 18207 10471 18213
rect 10413 18204 10425 18207
rect 10008 18176 10425 18204
rect 10008 18164 10014 18176
rect 10413 18173 10425 18176
rect 10459 18173 10471 18207
rect 13262 18204 13268 18216
rect 13223 18176 13268 18204
rect 10413 18167 10471 18173
rect 13262 18164 13268 18176
rect 13320 18164 13326 18216
rect 19429 18207 19487 18213
rect 19429 18173 19441 18207
rect 19475 18173 19487 18207
rect 20530 18204 20536 18216
rect 20491 18176 20536 18204
rect 19429 18167 19487 18173
rect 10689 18139 10747 18145
rect 10689 18105 10701 18139
rect 10735 18136 10747 18139
rect 19444 18136 19472 18167
rect 20530 18164 20536 18176
rect 20588 18164 20594 18216
rect 10735 18108 19472 18136
rect 10735 18105 10747 18108
rect 10689 18099 10747 18105
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 12986 17688 12992 17740
rect 13044 17728 13050 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 13044 17700 19717 17728
rect 13044 17688 13050 17700
rect 19705 17697 19717 17700
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 19886 17524 19892 17536
rect 19847 17496 19892 17524
rect 19886 17484 19892 17496
rect 19944 17484 19950 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 18966 17320 18972 17332
rect 18927 17292 18972 17320
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 12805 17187 12863 17193
rect 12805 17153 12817 17187
rect 12851 17184 12863 17187
rect 13262 17184 13268 17196
rect 12851 17156 13268 17184
rect 12851 17153 12863 17156
rect 12805 17147 12863 17153
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 20165 17187 20223 17193
rect 20165 17153 20177 17187
rect 20211 17184 20223 17187
rect 20530 17184 20536 17196
rect 20211 17156 20536 17184
rect 20211 17153 20223 17156
rect 20165 17147 20223 17153
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 12529 17119 12587 17125
rect 12529 17085 12541 17119
rect 12575 17116 12587 17119
rect 12618 17116 12624 17128
rect 12575 17088 12624 17116
rect 12575 17085 12587 17088
rect 12529 17079 12587 17085
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 18782 17116 18788 17128
rect 18743 17088 18788 17116
rect 18782 17076 18788 17088
rect 18840 17076 18846 17128
rect 19889 17119 19947 17125
rect 19889 17085 19901 17119
rect 19935 17085 19947 17119
rect 19889 17079 19947 17085
rect 10226 17008 10232 17060
rect 10284 17048 10290 17060
rect 19904 17048 19932 17079
rect 10284 17020 19932 17048
rect 10284 17008 10290 17020
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 18598 16776 18604 16788
rect 18559 16748 18604 16776
rect 18598 16736 18604 16748
rect 18656 16736 18662 16788
rect 12986 16708 12992 16720
rect 12947 16680 12992 16708
rect 12986 16668 12992 16680
rect 13044 16668 13050 16720
rect 16666 16668 16672 16720
rect 16724 16708 16730 16720
rect 16724 16680 18552 16708
rect 16724 16668 16730 16680
rect 12710 16640 12716 16652
rect 12671 16612 12716 16640
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 14734 16600 14740 16652
rect 14792 16640 14798 16652
rect 18417 16643 18475 16649
rect 18417 16640 18429 16643
rect 14792 16612 18429 16640
rect 14792 16600 14798 16612
rect 18417 16609 18429 16612
rect 18463 16609 18475 16643
rect 18524 16640 18552 16680
rect 18782 16668 18788 16720
rect 18840 16708 18846 16720
rect 19797 16711 19855 16717
rect 19797 16708 19809 16711
rect 18840 16680 19809 16708
rect 18840 16668 18846 16680
rect 19797 16677 19809 16680
rect 19843 16677 19855 16711
rect 19797 16671 19855 16677
rect 19521 16643 19579 16649
rect 19521 16640 19533 16643
rect 18524 16612 19533 16640
rect 18417 16603 18475 16609
rect 19521 16609 19533 16612
rect 19567 16609 19579 16643
rect 19521 16603 19579 16609
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 18509 16235 18567 16241
rect 18509 16201 18521 16235
rect 18555 16232 18567 16235
rect 18598 16232 18604 16244
rect 18555 16204 18604 16232
rect 18555 16201 18567 16204
rect 18509 16195 18567 16201
rect 18598 16192 18604 16204
rect 18656 16192 18662 16244
rect 17954 15988 17960 16040
rect 18012 16028 18018 16040
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 18012 16000 18337 16028
rect 18012 15988 18018 16000
rect 18325 15997 18337 16000
rect 18371 15997 18383 16031
rect 18325 15991 18383 15997
rect 19429 16031 19487 16037
rect 19429 15997 19441 16031
rect 19475 15997 19487 16031
rect 20530 16028 20536 16040
rect 20491 16000 20536 16028
rect 19429 15991 19487 15997
rect 18138 15920 18144 15972
rect 18196 15960 18202 15972
rect 19444 15960 19472 15991
rect 20530 15988 20536 16000
rect 20588 15988 20594 16040
rect 18196 15932 19472 15960
rect 18196 15920 18202 15932
rect 19242 15852 19248 15904
rect 19300 15892 19306 15904
rect 19613 15895 19671 15901
rect 19613 15892 19625 15895
rect 19300 15864 19625 15892
rect 19300 15852 19306 15864
rect 19613 15861 19625 15864
rect 19659 15861 19671 15895
rect 19613 15855 19671 15861
rect 20622 15852 20628 15904
rect 20680 15892 20686 15904
rect 20717 15895 20775 15901
rect 20717 15892 20729 15895
rect 20680 15864 20729 15892
rect 20680 15852 20686 15864
rect 20717 15861 20729 15864
rect 20763 15861 20775 15895
rect 20717 15855 20775 15861
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 18782 15688 18788 15700
rect 18743 15660 18788 15688
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 10781 15623 10839 15629
rect 10781 15589 10793 15623
rect 10827 15620 10839 15623
rect 14734 15620 14740 15632
rect 10827 15592 14740 15620
rect 10827 15589 10839 15592
rect 10781 15583 10839 15589
rect 14734 15580 14740 15592
rect 14792 15580 14798 15632
rect 10502 15552 10508 15564
rect 10463 15524 10508 15552
rect 10502 15512 10508 15524
rect 10560 15512 10566 15564
rect 18598 15552 18604 15564
rect 18559 15524 18604 15552
rect 18598 15512 18604 15524
rect 18656 15512 18662 15564
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15552 19763 15555
rect 19978 15552 19984 15564
rect 19751 15524 19984 15552
rect 19751 15521 19763 15524
rect 19705 15515 19763 15521
rect 19978 15512 19984 15524
rect 20036 15512 20042 15564
rect 19886 15348 19892 15360
rect 19847 15320 19892 15348
rect 19886 15308 19892 15320
rect 19944 15308 19950 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 19058 15144 19064 15156
rect 19019 15116 19064 15144
rect 19058 15104 19064 15116
rect 19116 15104 19122 15156
rect 13630 14968 13636 15020
rect 13688 15008 13694 15020
rect 13688 14980 20024 15008
rect 13688 14968 13694 14980
rect 7098 14900 7104 14952
rect 7156 14940 7162 14952
rect 7745 14943 7803 14949
rect 7745 14940 7757 14943
rect 7156 14912 7757 14940
rect 7156 14900 7162 14912
rect 7745 14909 7757 14912
rect 7791 14909 7803 14943
rect 9030 14940 9036 14952
rect 8991 14912 9036 14940
rect 7745 14903 7803 14909
rect 9030 14900 9036 14912
rect 9088 14900 9094 14952
rect 9309 14943 9367 14949
rect 9309 14909 9321 14943
rect 9355 14940 9367 14943
rect 17954 14940 17960 14952
rect 9355 14912 17960 14940
rect 9355 14909 9367 14912
rect 9309 14903 9367 14909
rect 17954 14900 17960 14912
rect 18012 14900 18018 14952
rect 18874 14940 18880 14952
rect 18835 14912 18880 14940
rect 18874 14900 18880 14912
rect 18932 14900 18938 14952
rect 19996 14949 20024 14980
rect 19981 14943 20039 14949
rect 19981 14909 19993 14943
rect 20027 14909 20039 14943
rect 19981 14903 20039 14909
rect 8021 14875 8079 14881
rect 8021 14841 8033 14875
rect 8067 14872 8079 14875
rect 18598 14872 18604 14884
rect 8067 14844 18604 14872
rect 8067 14841 8079 14844
rect 8021 14835 8079 14841
rect 18598 14832 18604 14844
rect 18656 14832 18662 14884
rect 18690 14832 18696 14884
rect 18748 14872 18754 14884
rect 20257 14875 20315 14881
rect 20257 14872 20269 14875
rect 18748 14844 20269 14872
rect 18748 14832 18754 14844
rect 20257 14841 20269 14844
rect 20303 14841 20315 14875
rect 20257 14835 20315 14841
rect 16945 14807 17003 14813
rect 16945 14773 16957 14807
rect 16991 14804 17003 14807
rect 19058 14804 19064 14816
rect 16991 14776 19064 14804
rect 16991 14773 17003 14776
rect 16945 14767 17003 14773
rect 19058 14764 19064 14776
rect 19116 14764 19122 14816
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 8297 14535 8355 14541
rect 8297 14501 8309 14535
rect 8343 14532 8355 14535
rect 18138 14532 18144 14544
rect 8343 14504 18144 14532
rect 8343 14501 8355 14504
rect 8297 14495 8355 14501
rect 18138 14492 18144 14504
rect 18196 14492 18202 14544
rect 18874 14492 18880 14544
rect 18932 14532 18938 14544
rect 19797 14535 19855 14541
rect 19797 14532 19809 14535
rect 18932 14504 19809 14532
rect 18932 14492 18938 14504
rect 19797 14501 19809 14504
rect 19843 14501 19855 14535
rect 19797 14495 19855 14501
rect 7190 14424 7196 14476
rect 7248 14464 7254 14476
rect 8021 14467 8079 14473
rect 8021 14464 8033 14467
rect 7248 14436 8033 14464
rect 7248 14424 7254 14436
rect 8021 14433 8033 14436
rect 8067 14433 8079 14467
rect 17310 14464 17316 14476
rect 17271 14436 17316 14464
rect 8021 14427 8079 14433
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 18417 14467 18475 14473
rect 18417 14433 18429 14467
rect 18463 14464 18475 14467
rect 18690 14464 18696 14476
rect 18463 14436 18696 14464
rect 18463 14433 18475 14436
rect 18417 14427 18475 14433
rect 18690 14424 18696 14436
rect 18748 14424 18754 14476
rect 19521 14467 19579 14473
rect 19521 14433 19533 14467
rect 19567 14433 19579 14467
rect 19521 14427 19579 14433
rect 12526 14396 12532 14408
rect 12487 14368 12532 14396
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 16301 14399 16359 14405
rect 16301 14365 16313 14399
rect 16347 14396 16359 14399
rect 17862 14396 17868 14408
rect 16347 14368 17868 14396
rect 16347 14365 16359 14368
rect 16301 14359 16359 14365
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 7650 14288 7656 14340
rect 7708 14328 7714 14340
rect 19536 14328 19564 14427
rect 7708 14300 19564 14328
rect 7708 14288 7714 14300
rect 17497 14263 17555 14269
rect 17497 14229 17509 14263
rect 17543 14260 17555 14263
rect 17770 14260 17776 14272
rect 17543 14232 17776 14260
rect 17543 14229 17555 14232
rect 17497 14223 17555 14229
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 18598 14260 18604 14272
rect 18559 14232 18604 14260
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 12437 14059 12495 14065
rect 12437 14025 12449 14059
rect 12483 14056 12495 14059
rect 12710 14056 12716 14068
rect 12483 14028 12716 14056
rect 12483 14025 12495 14028
rect 12437 14019 12495 14025
rect 12710 14016 12716 14028
rect 12768 14016 12774 14068
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 16574 14056 16580 14068
rect 15611 14028 16580 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 10962 13948 10968 14000
rect 11020 13988 11026 14000
rect 11020 13960 19840 13988
rect 11020 13948 11026 13960
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 16209 13923 16267 13929
rect 13044 13892 13089 13920
rect 13044 13880 13050 13892
rect 16209 13889 16221 13923
rect 16255 13920 16267 13923
rect 16482 13920 16488 13932
rect 16255 13892 16488 13920
rect 16255 13889 16267 13892
rect 16209 13883 16267 13889
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 17310 13880 17316 13932
rect 17368 13920 17374 13932
rect 18693 13923 18751 13929
rect 18693 13920 18705 13923
rect 17368 13892 18705 13920
rect 17368 13880 17374 13892
rect 18693 13889 18705 13892
rect 18739 13889 18751 13923
rect 18693 13883 18751 13889
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12584 13824 12817 13852
rect 12584 13812 12590 13824
rect 12805 13821 12817 13824
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 14642 13812 14648 13864
rect 14700 13852 14706 13864
rect 16025 13855 16083 13861
rect 16025 13852 16037 13855
rect 14700 13824 16037 13852
rect 14700 13812 14706 13824
rect 16025 13821 16037 13824
rect 16071 13821 16083 13855
rect 18506 13852 18512 13864
rect 18467 13824 18512 13852
rect 16025 13815 16083 13821
rect 18506 13812 18512 13824
rect 18564 13812 18570 13864
rect 19812 13861 19840 13960
rect 19978 13920 19984 13932
rect 19939 13892 19984 13920
rect 19978 13880 19984 13892
rect 20036 13880 20042 13932
rect 19797 13855 19855 13861
rect 19797 13821 19809 13855
rect 19843 13821 19855 13855
rect 19797 13815 19855 13821
rect 12342 13676 12348 13728
rect 12400 13716 12406 13728
rect 12897 13719 12955 13725
rect 12897 13716 12909 13719
rect 12400 13688 12909 13716
rect 12400 13676 12406 13688
rect 12897 13685 12909 13688
rect 12943 13685 12955 13719
rect 12897 13679 12955 13685
rect 14553 13719 14611 13725
rect 14553 13685 14565 13719
rect 14599 13716 14611 13719
rect 15562 13716 15568 13728
rect 14599 13688 15568 13716
rect 14599 13685 14611 13688
rect 14553 13679 14611 13685
rect 15562 13676 15568 13688
rect 15620 13676 15626 13728
rect 15930 13716 15936 13728
rect 15891 13688 15936 13716
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 12713 13515 12771 13521
rect 12713 13481 12725 13515
rect 12759 13512 12771 13515
rect 12986 13512 12992 13524
rect 12759 13484 12992 13512
rect 12759 13481 12771 13484
rect 12713 13475 12771 13481
rect 12986 13472 12992 13484
rect 13044 13472 13050 13524
rect 14185 13515 14243 13521
rect 14185 13481 14197 13515
rect 14231 13512 14243 13515
rect 15930 13512 15936 13524
rect 14231 13484 15936 13512
rect 14231 13481 14243 13484
rect 14185 13475 14243 13481
rect 15930 13472 15936 13484
rect 15988 13472 15994 13524
rect 17862 13472 17868 13524
rect 17920 13512 17926 13524
rect 17957 13515 18015 13521
rect 17957 13512 17969 13515
rect 17920 13484 17969 13512
rect 17920 13472 17926 13484
rect 17957 13481 17969 13484
rect 18003 13481 18015 13515
rect 17957 13475 18015 13481
rect 19150 13472 19156 13524
rect 19208 13512 19214 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 19208 13484 19257 13512
rect 19208 13472 19214 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 11600 13379 11658 13385
rect 11600 13345 11612 13379
rect 11646 13376 11658 13379
rect 11974 13376 11980 13388
rect 11646 13348 11980 13376
rect 11646 13345 11658 13348
rect 11600 13339 11658 13345
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 15194 13336 15200 13388
rect 15252 13376 15258 13388
rect 15289 13379 15347 13385
rect 15289 13376 15301 13379
rect 15252 13348 15301 13376
rect 15252 13336 15258 13348
rect 15289 13345 15301 13348
rect 15335 13345 15347 13379
rect 15289 13339 15347 13345
rect 15378 13336 15384 13388
rect 15436 13376 15442 13388
rect 15545 13379 15603 13385
rect 15545 13376 15557 13379
rect 15436 13348 15557 13376
rect 15436 13336 15442 13348
rect 15545 13345 15557 13348
rect 15591 13345 15603 13379
rect 15545 13339 15603 13345
rect 19334 13336 19340 13388
rect 19392 13376 19398 13388
rect 19613 13379 19671 13385
rect 19613 13376 19625 13379
rect 19392 13348 19625 13376
rect 19392 13336 19398 13348
rect 19613 13345 19625 13348
rect 19659 13345 19671 13379
rect 19613 13339 19671 13345
rect 10134 13268 10140 13320
rect 10192 13308 10198 13320
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 10192 13280 11345 13308
rect 10192 13268 10198 13280
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 18046 13308 18052 13320
rect 18007 13280 18052 13308
rect 11333 13271 11391 13277
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 18138 13268 18144 13320
rect 18196 13308 18202 13320
rect 18196 13280 18241 13308
rect 18196 13268 18202 13280
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19484 13280 19717 13308
rect 19484 13268 19490 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 19794 13268 19800 13320
rect 19852 13308 19858 13320
rect 19852 13280 19897 13308
rect 19852 13268 19858 13280
rect 17589 13243 17647 13249
rect 17589 13209 17601 13243
rect 17635 13240 17647 13243
rect 18506 13240 18512 13252
rect 17635 13212 18512 13240
rect 17635 13209 17647 13212
rect 17589 13203 17647 13209
rect 18506 13200 18512 13212
rect 18564 13200 18570 13252
rect 16482 13132 16488 13184
rect 16540 13172 16546 13184
rect 16669 13175 16727 13181
rect 16669 13172 16681 13175
rect 16540 13144 16681 13172
rect 16540 13132 16546 13144
rect 16669 13141 16681 13144
rect 16715 13141 16727 13175
rect 16669 13135 16727 13141
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 15194 12928 15200 12980
rect 15252 12968 15258 12980
rect 15473 12971 15531 12977
rect 15473 12968 15485 12971
rect 15252 12940 15485 12968
rect 15252 12928 15258 12940
rect 15473 12937 15485 12940
rect 15519 12937 15531 12971
rect 15473 12931 15531 12937
rect 9214 12792 9220 12844
rect 9272 12832 9278 12844
rect 10134 12832 10140 12844
rect 9272 12804 10140 12832
rect 9272 12792 9278 12804
rect 10134 12792 10140 12804
rect 10192 12792 10198 12844
rect 15488 12832 15516 12931
rect 15749 12835 15807 12841
rect 15749 12832 15761 12835
rect 15488 12804 15761 12832
rect 15749 12801 15761 12804
rect 15795 12801 15807 12835
rect 20530 12832 20536 12844
rect 20491 12804 20536 12832
rect 15749 12795 15807 12801
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12764 12863 12767
rect 12894 12764 12900 12776
rect 12851 12736 12900 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 15654 12764 15660 12776
rect 15615 12736 15660 12764
rect 15654 12724 15660 12736
rect 15712 12724 15718 12776
rect 15764 12764 15792 12795
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 16016 12767 16074 12773
rect 15764 12736 15976 12764
rect 10404 12699 10462 12705
rect 10404 12665 10416 12699
rect 10450 12696 10462 12699
rect 10594 12696 10600 12708
rect 10450 12668 10600 12696
rect 10450 12665 10462 12668
rect 10404 12659 10462 12665
rect 10594 12656 10600 12668
rect 10652 12656 10658 12708
rect 12986 12656 12992 12708
rect 13044 12705 13050 12708
rect 13044 12699 13108 12705
rect 13044 12665 13062 12699
rect 13096 12665 13108 12699
rect 13044 12659 13108 12665
rect 13044 12656 13050 12659
rect 11517 12631 11575 12637
rect 11517 12597 11529 12631
rect 11563 12628 11575 12631
rect 11974 12628 11980 12640
rect 11563 12600 11980 12628
rect 11563 12597 11575 12600
rect 11517 12591 11575 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 14182 12628 14188 12640
rect 14143 12600 14188 12628
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 15948 12628 15976 12736
rect 16016 12733 16028 12767
rect 16062 12764 16074 12767
rect 16482 12764 16488 12776
rect 16062 12736 16488 12764
rect 16062 12733 16074 12736
rect 16016 12727 16074 12733
rect 16482 12724 16488 12736
rect 16540 12724 16546 12776
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12764 18107 12767
rect 19058 12764 19064 12776
rect 18095 12736 19064 12764
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 18064 12696 18092 12727
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 20254 12764 20260 12776
rect 20215 12736 20260 12764
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 16500 12668 18092 12696
rect 16500 12640 16528 12668
rect 18138 12656 18144 12708
rect 18196 12696 18202 12708
rect 18294 12699 18352 12705
rect 18294 12696 18306 12699
rect 18196 12668 18306 12696
rect 18196 12656 18202 12668
rect 18294 12665 18306 12668
rect 18340 12665 18352 12699
rect 18294 12659 18352 12665
rect 16482 12628 16488 12640
rect 15948 12600 16488 12628
rect 16482 12588 16488 12600
rect 16540 12588 16546 12640
rect 17129 12631 17187 12637
rect 17129 12597 17141 12631
rect 17175 12628 17187 12631
rect 17310 12628 17316 12640
rect 17175 12600 17316 12628
rect 17175 12597 17187 12600
rect 17129 12591 17187 12597
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 18690 12588 18696 12640
rect 18748 12628 18754 12640
rect 19429 12631 19487 12637
rect 19429 12628 19441 12631
rect 18748 12600 19441 12628
rect 18748 12588 18754 12600
rect 19429 12597 19441 12600
rect 19475 12597 19487 12631
rect 19429 12591 19487 12597
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 9861 12427 9919 12433
rect 9861 12393 9873 12427
rect 9907 12424 9919 12427
rect 10502 12424 10508 12436
rect 9907 12396 10508 12424
rect 9907 12393 9919 12396
rect 9861 12387 9919 12393
rect 10502 12384 10508 12396
rect 10560 12384 10566 12436
rect 11425 12427 11483 12433
rect 11425 12393 11437 12427
rect 11471 12424 11483 12427
rect 12342 12424 12348 12436
rect 11471 12396 12348 12424
rect 11471 12393 11483 12396
rect 11425 12387 11483 12393
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 15841 12427 15899 12433
rect 15841 12393 15853 12427
rect 15887 12424 15899 12427
rect 17862 12424 17868 12436
rect 15887 12396 17868 12424
rect 15887 12393 15899 12396
rect 15841 12387 15899 12393
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 18138 12424 18144 12436
rect 18099 12396 18144 12424
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 11885 12359 11943 12365
rect 11885 12325 11897 12359
rect 11931 12356 11943 12359
rect 15102 12356 15108 12368
rect 11931 12328 15108 12356
rect 11931 12325 11943 12328
rect 11885 12319 11943 12325
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 17402 12356 17408 12368
rect 15672 12328 17408 12356
rect 8573 12291 8631 12297
rect 8573 12257 8585 12291
rect 8619 12288 8631 12291
rect 10229 12291 10287 12297
rect 10229 12288 10241 12291
rect 8619 12260 10241 12288
rect 8619 12257 8631 12260
rect 8573 12251 8631 12257
rect 10229 12257 10241 12260
rect 10275 12257 10287 12291
rect 10229 12251 10287 12257
rect 11793 12291 11851 12297
rect 11793 12257 11805 12291
rect 11839 12257 11851 12291
rect 11793 12251 11851 12257
rect 10318 12220 10324 12232
rect 10279 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10505 12223 10563 12229
rect 10505 12189 10517 12223
rect 10551 12220 10563 12223
rect 10594 12220 10600 12232
rect 10551 12192 10600 12220
rect 10551 12189 10563 12192
rect 10505 12183 10563 12189
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 11808 12220 11836 12251
rect 12894 12248 12900 12300
rect 12952 12288 12958 12300
rect 12989 12291 13047 12297
rect 12989 12288 13001 12291
rect 12952 12260 13001 12288
rect 12952 12248 12958 12260
rect 12989 12257 13001 12260
rect 13035 12257 13047 12291
rect 12989 12251 13047 12257
rect 13256 12291 13314 12297
rect 13256 12257 13268 12291
rect 13302 12288 13314 12291
rect 13814 12288 13820 12300
rect 13302 12260 13820 12288
rect 13302 12257 13314 12260
rect 13256 12251 13314 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 15672 12297 15700 12328
rect 17402 12316 17408 12328
rect 17460 12316 17466 12368
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 16482 12248 16488 12300
rect 16540 12288 16546 12300
rect 16761 12291 16819 12297
rect 16761 12288 16773 12291
rect 16540 12260 16773 12288
rect 16540 12248 16546 12260
rect 16761 12257 16773 12260
rect 16807 12257 16819 12291
rect 16761 12251 16819 12257
rect 17028 12291 17086 12297
rect 17028 12257 17040 12291
rect 17074 12288 17086 12291
rect 17310 12288 17316 12300
rect 17074 12260 17316 12288
rect 17074 12257 17086 12260
rect 17028 12251 17086 12257
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 18874 12248 18880 12300
rect 18932 12288 18938 12300
rect 19613 12291 19671 12297
rect 19613 12288 19625 12291
rect 18932 12260 19625 12288
rect 18932 12248 18938 12260
rect 19613 12257 19625 12260
rect 19659 12257 19671 12291
rect 19613 12251 19671 12257
rect 19702 12248 19708 12300
rect 19760 12288 19766 12300
rect 19760 12260 19805 12288
rect 19760 12248 19766 12260
rect 11882 12220 11888 12232
rect 11808 12192 11888 12220
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 11974 12180 11980 12232
rect 12032 12220 12038 12232
rect 19889 12223 19947 12229
rect 12032 12192 12077 12220
rect 12032 12180 12038 12192
rect 19889 12189 19901 12223
rect 19935 12220 19947 12223
rect 20622 12220 20628 12232
rect 19935 12192 20628 12220
rect 19935 12189 19947 12192
rect 19889 12183 19947 12189
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 9582 12044 9588 12096
rect 9640 12084 9646 12096
rect 14274 12084 14280 12096
rect 9640 12056 14280 12084
rect 9640 12044 9646 12056
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 14369 12087 14427 12093
rect 14369 12053 14381 12087
rect 14415 12084 14427 12087
rect 15378 12084 15384 12096
rect 14415 12056 15384 12084
rect 14415 12053 14427 12056
rect 14369 12047 14427 12053
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 19245 12087 19303 12093
rect 19245 12053 19257 12087
rect 19291 12084 19303 12087
rect 19518 12084 19524 12096
rect 19291 12056 19524 12084
rect 19291 12053 19303 12056
rect 19245 12047 19303 12053
rect 19518 12044 19524 12056
rect 19576 12044 19582 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 10594 11880 10600 11892
rect 10555 11852 10600 11880
rect 10594 11840 10600 11852
rect 10652 11840 10658 11892
rect 13081 11883 13139 11889
rect 13081 11849 13093 11883
rect 13127 11880 13139 11883
rect 13906 11880 13912 11892
rect 13127 11852 13912 11880
rect 13127 11849 13139 11852
rect 13081 11843 13139 11849
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 14642 11880 14648 11892
rect 14603 11852 14648 11880
rect 14642 11840 14648 11852
rect 14700 11840 14706 11892
rect 16209 11883 16267 11889
rect 16209 11849 16221 11883
rect 16255 11880 16267 11883
rect 16666 11880 16672 11892
rect 16255 11852 16672 11880
rect 16255 11849 16267 11852
rect 16209 11843 16267 11849
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 1210 11704 1216 11756
rect 1268 11744 1274 11756
rect 13725 11747 13783 11753
rect 1268 11716 9352 11744
rect 1268 11704 1274 11716
rect 9214 11676 9220 11688
rect 9175 11648 9220 11676
rect 9214 11636 9220 11648
rect 9272 11636 9278 11688
rect 9324 11676 9352 11716
rect 13725 11713 13737 11747
rect 13771 11744 13783 11747
rect 13814 11744 13820 11756
rect 13771 11716 13820 11744
rect 13771 11713 13783 11716
rect 13725 11707 13783 11713
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 15102 11744 15108 11756
rect 14700 11716 15108 11744
rect 14700 11704 14706 11716
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11744 15347 11747
rect 15378 11744 15384 11756
rect 15335 11716 15384 11744
rect 15335 11713 15347 11716
rect 15289 11707 15347 11713
rect 15378 11704 15384 11716
rect 15436 11704 15442 11756
rect 15470 11704 15476 11756
rect 15528 11744 15534 11756
rect 16761 11747 16819 11753
rect 16761 11744 16773 11747
rect 15528 11716 16773 11744
rect 15528 11704 15534 11716
rect 16761 11713 16773 11716
rect 16807 11713 16819 11747
rect 16761 11707 16819 11713
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11744 18107 11747
rect 19334 11744 19340 11756
rect 18095 11716 19340 11744
rect 18095 11713 18107 11716
rect 18049 11707 18107 11713
rect 19334 11704 19340 11716
rect 19392 11704 19398 11756
rect 19518 11744 19524 11756
rect 19479 11716 19524 11744
rect 19518 11704 19524 11716
rect 19576 11704 19582 11756
rect 19705 11747 19763 11753
rect 19705 11713 19717 11747
rect 19751 11744 19763 11747
rect 20806 11744 20812 11756
rect 19751 11716 20812 11744
rect 19751 11713 19763 11716
rect 19705 11707 19763 11713
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 15013 11679 15071 11685
rect 15013 11676 15025 11679
rect 9324 11648 15025 11676
rect 15013 11645 15025 11648
rect 15059 11645 15071 11679
rect 15013 11639 15071 11645
rect 15562 11636 15568 11688
rect 15620 11676 15626 11688
rect 16577 11679 16635 11685
rect 16577 11676 16589 11679
rect 15620 11648 16589 11676
rect 15620 11636 15626 11648
rect 16577 11645 16589 11648
rect 16623 11645 16635 11679
rect 16577 11639 16635 11645
rect 9484 11611 9542 11617
rect 9484 11577 9496 11611
rect 9530 11608 9542 11611
rect 9858 11608 9864 11620
rect 9530 11580 9864 11608
rect 9530 11577 9542 11580
rect 9484 11571 9542 11577
rect 9858 11568 9864 11580
rect 9916 11568 9922 11620
rect 12618 11568 12624 11620
rect 12676 11608 12682 11620
rect 19429 11611 19487 11617
rect 12676 11580 19196 11608
rect 12676 11568 12682 11580
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 12710 11540 12716 11552
rect 8352 11512 12716 11540
rect 8352 11500 8358 11512
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 13446 11540 13452 11552
rect 13407 11512 13452 11540
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 13538 11500 13544 11552
rect 13596 11540 13602 11552
rect 16666 11540 16672 11552
rect 13596 11512 13641 11540
rect 16627 11512 16672 11540
rect 13596 11500 13602 11512
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 16850 11500 16856 11552
rect 16908 11540 16914 11552
rect 19061 11543 19119 11549
rect 19061 11540 19073 11543
rect 16908 11512 19073 11540
rect 16908 11500 16914 11512
rect 19061 11509 19073 11512
rect 19107 11509 19119 11543
rect 19168 11540 19196 11580
rect 19429 11577 19441 11611
rect 19475 11608 19487 11611
rect 20625 11611 20683 11617
rect 20625 11608 20637 11611
rect 19475 11580 20637 11608
rect 19475 11577 19487 11580
rect 19429 11571 19487 11577
rect 20625 11577 20637 11580
rect 20671 11577 20683 11611
rect 20625 11571 20683 11577
rect 20162 11540 20168 11552
rect 19168 11512 20168 11540
rect 19061 11503 19119 11509
rect 20162 11500 20168 11512
rect 20220 11500 20226 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 9769 11339 9827 11345
rect 9769 11305 9781 11339
rect 9815 11336 9827 11339
rect 10318 11336 10324 11348
rect 9815 11308 10324 11336
rect 9815 11305 9827 11308
rect 9769 11299 9827 11305
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 11974 11296 11980 11348
rect 12032 11336 12038 11348
rect 12032 11308 13400 11336
rect 12032 11296 12038 11308
rect 4062 11228 4068 11280
rect 4120 11268 4126 11280
rect 12618 11268 12624 11280
rect 4120 11240 12624 11268
rect 4120 11228 4126 11240
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 12710 11228 12716 11280
rect 12768 11268 12774 11280
rect 13081 11271 13139 11277
rect 13081 11268 13093 11271
rect 12768 11240 13093 11268
rect 12768 11228 12774 11240
rect 13081 11237 13093 11240
rect 13127 11237 13139 11271
rect 13081 11231 13139 11237
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 10137 11203 10195 11209
rect 10137 11200 10149 11203
rect 9732 11172 10149 11200
rect 9732 11160 9738 11172
rect 10137 11169 10149 11172
rect 10183 11169 10195 11203
rect 10137 11163 10195 11169
rect 10229 11203 10287 11209
rect 10229 11169 10241 11203
rect 10275 11200 10287 11203
rect 10410 11200 10416 11212
rect 10275 11172 10416 11200
rect 10275 11169 10287 11172
rect 10229 11163 10287 11169
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 11974 11209 11980 11212
rect 11969 11200 11980 11209
rect 11935 11172 11980 11200
rect 11969 11163 11980 11172
rect 11974 11160 11980 11163
rect 12032 11160 12038 11212
rect 13372 11200 13400 11308
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 15289 11339 15347 11345
rect 15289 11336 15301 11339
rect 13504 11308 15301 11336
rect 13504 11296 13510 11308
rect 15289 11305 15301 11308
rect 15335 11305 15347 11339
rect 15289 11299 15347 11305
rect 15654 11296 15660 11348
rect 15712 11336 15718 11348
rect 16114 11336 16120 11348
rect 15712 11308 16120 11336
rect 15712 11296 15718 11308
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 16761 11339 16819 11345
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 18046 11336 18052 11348
rect 16807 11308 18052 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 19794 11336 19800 11348
rect 19755 11308 19800 11336
rect 19794 11296 19800 11308
rect 19852 11296 19858 11348
rect 14274 11228 14280 11280
rect 14332 11268 14338 11280
rect 16577 11271 16635 11277
rect 16577 11268 16589 11271
rect 14332 11240 16589 11268
rect 14332 11228 14338 11240
rect 16577 11237 16589 11240
rect 16623 11268 16635 11271
rect 17129 11271 17187 11277
rect 17129 11268 17141 11271
rect 16623 11240 17141 11268
rect 16623 11237 16635 11240
rect 16577 11231 16635 11237
rect 17129 11237 17141 11240
rect 17175 11237 17187 11271
rect 17129 11231 17187 11237
rect 14645 11203 14703 11209
rect 14645 11200 14657 11203
rect 13372 11172 14657 11200
rect 14645 11169 14657 11172
rect 14691 11200 14703 11203
rect 16301 11203 16359 11209
rect 16301 11200 16313 11203
rect 14691 11172 16313 11200
rect 14691 11169 14703 11172
rect 14645 11163 14703 11169
rect 16301 11169 16313 11172
rect 16347 11169 16359 11203
rect 17218 11200 17224 11212
rect 17179 11172 17224 11200
rect 16301 11163 16359 11169
rect 17218 11160 17224 11172
rect 17276 11160 17282 11212
rect 18138 11160 18144 11212
rect 18196 11200 18202 11212
rect 18690 11209 18696 11212
rect 18673 11203 18696 11209
rect 18673 11200 18685 11203
rect 18196 11172 18685 11200
rect 18196 11160 18202 11172
rect 18673 11169 18685 11172
rect 18748 11200 18754 11212
rect 18748 11172 18821 11200
rect 18673 11163 18696 11169
rect 18690 11160 18696 11163
rect 18748 11160 18754 11172
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11101 10379 11135
rect 17310 11132 17316 11144
rect 17271 11104 17316 11132
rect 10321 11095 10379 11101
rect 9858 11024 9864 11076
rect 9916 11064 9922 11076
rect 10336 11064 10364 11095
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 18417 11135 18475 11141
rect 18417 11101 18429 11135
rect 18463 11101 18475 11135
rect 18417 11095 18475 11101
rect 9916 11036 10364 11064
rect 11793 11067 11851 11073
rect 9916 11024 9922 11036
rect 11793 11033 11805 11067
rect 11839 11064 11851 11067
rect 12158 11064 12164 11076
rect 11839 11036 12164 11064
rect 11839 11033 11851 11036
rect 11793 11027 11851 11033
rect 12158 11024 12164 11036
rect 12216 11024 12222 11076
rect 11882 10956 11888 11008
rect 11940 10996 11946 11008
rect 15286 10996 15292 11008
rect 11940 10968 15292 10996
rect 11940 10956 11946 10968
rect 15286 10956 15292 10968
rect 15344 10956 15350 11008
rect 16298 10956 16304 11008
rect 16356 10996 16362 11008
rect 18432 10996 18460 11095
rect 19058 10996 19064 11008
rect 16356 10968 19064 10996
rect 16356 10956 16362 10968
rect 19058 10956 19064 10968
rect 19116 10956 19122 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 9858 10792 9864 10804
rect 9819 10764 9864 10792
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 10778 10792 10784 10804
rect 10739 10764 10784 10792
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 10870 10752 10876 10804
rect 10928 10792 10934 10804
rect 13814 10792 13820 10804
rect 10928 10764 13676 10792
rect 13775 10764 13820 10792
rect 10928 10752 10934 10764
rect 11425 10659 11483 10665
rect 11425 10625 11437 10659
rect 11471 10656 11483 10659
rect 11698 10656 11704 10668
rect 11471 10628 11704 10656
rect 11471 10625 11483 10628
rect 11425 10619 11483 10625
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 9122 10588 9128 10600
rect 8527 10560 9128 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 11790 10588 11796 10600
rect 9324 10560 11796 10588
rect 8748 10523 8806 10529
rect 8748 10489 8760 10523
rect 8794 10520 8806 10523
rect 8938 10520 8944 10532
rect 8794 10492 8944 10520
rect 8794 10489 8806 10492
rect 8748 10483 8806 10489
rect 8938 10480 8944 10492
rect 8996 10480 9002 10532
rect 5074 10412 5080 10464
rect 5132 10452 5138 10464
rect 9324 10452 9352 10560
rect 11790 10548 11796 10560
rect 11848 10548 11854 10600
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10588 12495 10591
rect 12483 10560 12940 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 12912 10532 12940 10560
rect 11149 10523 11207 10529
rect 11149 10489 11161 10523
rect 11195 10520 11207 10523
rect 11195 10492 12480 10520
rect 11195 10489 11207 10492
rect 11149 10483 11207 10489
rect 12452 10464 12480 10492
rect 12618 10480 12624 10532
rect 12676 10529 12682 10532
rect 12676 10523 12740 10529
rect 12676 10489 12694 10523
rect 12728 10489 12740 10523
rect 12676 10483 12740 10489
rect 12676 10480 12682 10483
rect 12894 10480 12900 10532
rect 12952 10480 12958 10532
rect 13648 10520 13676 10764
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 15470 10792 15476 10804
rect 14108 10764 15056 10792
rect 15431 10764 15476 10792
rect 14108 10665 14136 10764
rect 15028 10724 15056 10764
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 16393 10795 16451 10801
rect 16393 10761 16405 10795
rect 16439 10792 16451 10795
rect 19426 10792 19432 10804
rect 16439 10764 19432 10792
rect 16439 10761 16451 10764
rect 16393 10755 16451 10761
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 20622 10752 20628 10804
rect 20680 10792 20686 10804
rect 20809 10795 20867 10801
rect 20809 10792 20821 10795
rect 20680 10764 20821 10792
rect 20680 10752 20686 10764
rect 20809 10761 20821 10764
rect 20855 10761 20867 10795
rect 20809 10755 20867 10761
rect 16298 10724 16304 10736
rect 15028 10696 16304 10724
rect 16298 10684 16304 10696
rect 16356 10684 16362 10736
rect 14093 10659 14151 10665
rect 14093 10625 14105 10659
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 18138 10656 18144 10668
rect 17083 10628 18144 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 18138 10616 18144 10628
rect 18196 10616 18202 10668
rect 19058 10616 19064 10668
rect 19116 10656 19122 10668
rect 19429 10659 19487 10665
rect 19429 10656 19441 10659
rect 19116 10628 19441 10656
rect 19116 10616 19122 10628
rect 19429 10625 19441 10628
rect 19475 10625 19487 10659
rect 19429 10619 19487 10625
rect 14182 10548 14188 10600
rect 14240 10588 14246 10600
rect 14349 10591 14407 10597
rect 14349 10588 14361 10591
rect 14240 10560 14361 10588
rect 14240 10548 14246 10560
rect 14349 10557 14361 10560
rect 14395 10557 14407 10591
rect 14349 10551 14407 10557
rect 18325 10591 18383 10597
rect 18325 10557 18337 10591
rect 18371 10588 18383 10591
rect 18598 10588 18604 10600
rect 18371 10560 18604 10588
rect 18371 10557 18383 10560
rect 18325 10551 18383 10557
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 16761 10523 16819 10529
rect 16761 10520 16773 10523
rect 13648 10492 16773 10520
rect 16761 10489 16773 10492
rect 16807 10489 16819 10523
rect 16761 10483 16819 10489
rect 19696 10523 19754 10529
rect 19696 10489 19708 10523
rect 19742 10520 19754 10523
rect 19794 10520 19800 10532
rect 19742 10492 19800 10520
rect 19742 10489 19754 10492
rect 19696 10483 19754 10489
rect 19794 10480 19800 10492
rect 19852 10480 19858 10532
rect 11238 10452 11244 10464
rect 5132 10424 9352 10452
rect 11199 10424 11244 10452
rect 5132 10412 5138 10424
rect 11238 10412 11244 10424
rect 11296 10412 11302 10464
rect 12434 10412 12440 10464
rect 12492 10412 12498 10464
rect 16853 10455 16911 10461
rect 16853 10421 16865 10455
rect 16899 10452 16911 10455
rect 16942 10452 16948 10464
rect 16899 10424 16948 10452
rect 16899 10421 16911 10424
rect 16853 10415 16911 10421
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 18509 10455 18567 10461
rect 18509 10421 18521 10455
rect 18555 10452 18567 10455
rect 20346 10452 20352 10464
rect 18555 10424 20352 10452
rect 18555 10421 18567 10424
rect 18509 10415 18567 10421
rect 20346 10412 20352 10424
rect 20404 10412 20410 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 8021 10251 8079 10257
rect 8021 10217 8033 10251
rect 8067 10248 8079 10251
rect 9030 10248 9036 10260
rect 8067 10220 9036 10248
rect 8067 10217 8079 10220
rect 8021 10211 8079 10217
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9677 10251 9735 10257
rect 9677 10217 9689 10251
rect 9723 10248 9735 10251
rect 10226 10248 10232 10260
rect 9723 10220 10232 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 10226 10208 10232 10220
rect 10284 10208 10290 10260
rect 11882 10248 11888 10260
rect 11256 10220 11888 10248
rect 10045 10183 10103 10189
rect 10045 10149 10057 10183
rect 10091 10180 10103 10183
rect 11256 10180 11284 10220
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 13081 10251 13139 10257
rect 13081 10217 13093 10251
rect 13127 10248 13139 10251
rect 13998 10248 14004 10260
rect 13127 10220 13299 10248
rect 13959 10220 14004 10248
rect 13127 10217 13139 10220
rect 13081 10211 13139 10217
rect 13271 10192 13299 10220
rect 13998 10208 14004 10220
rect 14056 10208 14062 10260
rect 14093 10251 14151 10257
rect 14093 10217 14105 10251
rect 14139 10248 14151 10251
rect 17218 10248 17224 10260
rect 14139 10220 17224 10248
rect 14139 10217 14151 10220
rect 14093 10211 14151 10217
rect 17218 10208 17224 10220
rect 17276 10208 17282 10260
rect 18966 10248 18972 10260
rect 18927 10220 18972 10248
rect 18966 10208 18972 10220
rect 19024 10208 19030 10260
rect 10091 10152 11284 10180
rect 11508 10183 11566 10189
rect 10091 10149 10103 10152
rect 10045 10143 10103 10149
rect 11508 10149 11520 10183
rect 11554 10180 11566 10183
rect 11698 10180 11704 10192
rect 11554 10152 11704 10180
rect 11554 10149 11566 10152
rect 11508 10143 11566 10149
rect 11698 10140 11704 10152
rect 11756 10140 11762 10192
rect 13262 10140 13268 10192
rect 13320 10140 13326 10192
rect 16568 10183 16626 10189
rect 13556 10152 16436 10180
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10112 7067 10115
rect 8389 10115 8447 10121
rect 8389 10112 8401 10115
rect 7055 10084 8401 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 8389 10081 8401 10084
rect 8435 10081 8447 10115
rect 8389 10075 8447 10081
rect 10137 10115 10195 10121
rect 10137 10081 10149 10115
rect 10183 10112 10195 10115
rect 11790 10112 11796 10124
rect 10183 10084 11796 10112
rect 10183 10081 10195 10084
rect 10137 10075 10195 10081
rect 11790 10072 11796 10084
rect 11848 10072 11854 10124
rect 13173 10115 13231 10121
rect 13173 10081 13185 10115
rect 13219 10112 13231 10115
rect 13556 10112 13584 10152
rect 16298 10112 16304 10124
rect 13219 10084 13584 10112
rect 16259 10084 16304 10112
rect 13219 10081 13231 10084
rect 13173 10075 13231 10081
rect 1762 10004 1768 10056
rect 1820 10044 1826 10056
rect 8478 10044 8484 10056
rect 1820 10016 7788 10044
rect 8439 10016 8484 10044
rect 1820 10004 1826 10016
rect 7760 9976 7788 10016
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 8665 10047 8723 10053
rect 8665 10013 8677 10047
rect 8711 10044 8723 10047
rect 8938 10044 8944 10056
rect 8711 10016 8944 10044
rect 8711 10013 8723 10016
rect 8665 10007 8723 10013
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 10226 10044 10232 10056
rect 9048 10016 10232 10044
rect 9048 9976 9076 10016
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10044 10379 10047
rect 11054 10044 11060 10056
rect 10367 10016 11060 10044
rect 10367 10013 10379 10016
rect 10321 10007 10379 10013
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 11241 10047 11299 10053
rect 11241 10013 11253 10047
rect 11287 10013 11299 10047
rect 13188 10044 13216 10075
rect 16298 10072 16304 10084
rect 16356 10072 16362 10124
rect 16408 10112 16436 10152
rect 16568 10149 16580 10183
rect 16614 10180 16626 10183
rect 20806 10180 20812 10192
rect 16614 10152 20812 10180
rect 16614 10149 16626 10152
rect 16568 10143 16626 10149
rect 20806 10140 20812 10152
rect 20864 10140 20870 10192
rect 17310 10112 17316 10124
rect 16408 10084 17316 10112
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 18874 10112 18880 10124
rect 18835 10084 18880 10112
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 11241 10007 11299 10013
rect 12268 10016 13216 10044
rect 13265 10047 13323 10053
rect 7760 9948 9076 9976
rect 9214 9936 9220 9988
rect 9272 9976 9278 9988
rect 11256 9976 11284 10007
rect 9272 9948 11284 9976
rect 9272 9936 9278 9948
rect 10410 9868 10416 9920
rect 10468 9908 10474 9920
rect 12268 9908 12296 10016
rect 13265 10013 13277 10047
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 12618 9976 12624 9988
rect 12531 9948 12624 9976
rect 12618 9936 12624 9948
rect 12676 9976 12682 9988
rect 13280 9976 13308 10007
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 15289 10047 15347 10053
rect 14240 10016 14285 10044
rect 14240 10004 14246 10016
rect 15289 10013 15301 10047
rect 15335 10044 15347 10047
rect 16206 10044 16212 10056
rect 15335 10016 16212 10044
rect 15335 10013 15347 10016
rect 15289 10007 15347 10013
rect 16206 10004 16212 10016
rect 16264 10004 16270 10056
rect 19061 10047 19119 10053
rect 19061 10013 19073 10047
rect 19107 10013 19119 10047
rect 19061 10007 19119 10013
rect 19076 9976 19104 10007
rect 12676 9948 13308 9976
rect 17696 9948 19104 9976
rect 12676 9936 12682 9948
rect 17696 9920 17724 9948
rect 10468 9880 12296 9908
rect 12713 9911 12771 9917
rect 10468 9868 10474 9880
rect 12713 9877 12725 9911
rect 12759 9908 12771 9911
rect 13538 9908 13544 9920
rect 12759 9880 13544 9908
rect 12759 9877 12771 9880
rect 12713 9871 12771 9877
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 13633 9911 13691 9917
rect 13633 9877 13645 9911
rect 13679 9908 13691 9911
rect 16666 9908 16672 9920
rect 13679 9880 16672 9908
rect 13679 9877 13691 9880
rect 13633 9871 13691 9877
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 17678 9908 17684 9920
rect 17639 9880 17684 9908
rect 17678 9868 17684 9880
rect 17736 9868 17742 9920
rect 17770 9868 17776 9920
rect 17828 9908 17834 9920
rect 18509 9911 18567 9917
rect 18509 9908 18521 9911
rect 17828 9880 18521 9908
rect 17828 9868 17834 9880
rect 18509 9877 18521 9880
rect 18555 9877 18567 9911
rect 18509 9871 18567 9877
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 8938 9704 8944 9716
rect 8899 9676 8944 9704
rect 8938 9664 8944 9676
rect 8996 9664 9002 9716
rect 11517 9707 11575 9713
rect 11517 9673 11529 9707
rect 11563 9704 11575 9707
rect 11698 9704 11704 9716
rect 11563 9676 11704 9704
rect 11563 9673 11575 9676
rect 11517 9667 11575 9673
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 20806 9704 20812 9716
rect 20767 9676 20812 9704
rect 20806 9664 20812 9676
rect 20864 9664 20870 9716
rect 9214 9596 9220 9648
rect 9272 9636 9278 9648
rect 9861 9639 9919 9645
rect 9861 9636 9873 9639
rect 9272 9608 9873 9636
rect 9272 9596 9278 9608
rect 9861 9605 9873 9608
rect 9907 9636 9919 9639
rect 9907 9608 10180 9636
rect 9907 9605 9919 9608
rect 9861 9599 9919 9605
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9500 7619 9503
rect 9232 9500 9260 9596
rect 10152 9577 10180 9608
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9537 10195 9571
rect 12434 9568 12440 9580
rect 12395 9540 12440 9568
rect 10137 9531 10195 9537
rect 12434 9528 12440 9540
rect 12492 9528 12498 9580
rect 7607 9472 9260 9500
rect 10045 9503 10103 9509
rect 7607 9469 7619 9472
rect 7561 9463 7619 9469
rect 10045 9469 10057 9503
rect 10091 9469 10103 9503
rect 12158 9500 12164 9512
rect 10045 9463 10103 9469
rect 10244 9472 12164 9500
rect 7828 9435 7886 9441
rect 7828 9401 7840 9435
rect 7874 9432 7886 9435
rect 8570 9432 8576 9444
rect 7874 9404 8576 9432
rect 7874 9401 7886 9404
rect 7828 9395 7886 9401
rect 8570 9392 8576 9404
rect 8628 9392 8634 9444
rect 10060 9432 10088 9463
rect 10244 9432 10272 9472
rect 12158 9460 12164 9472
rect 12216 9460 12222 9512
rect 13538 9500 13544 9512
rect 13499 9472 13544 9500
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 13808 9503 13866 9509
rect 13808 9469 13820 9503
rect 13854 9500 13866 9503
rect 15470 9500 15476 9512
rect 13854 9472 15476 9500
rect 13854 9469 13866 9472
rect 13808 9463 13866 9469
rect 15470 9460 15476 9472
rect 15528 9460 15534 9512
rect 15749 9503 15807 9509
rect 15749 9469 15761 9503
rect 15795 9469 15807 9503
rect 15749 9463 15807 9469
rect 16016 9503 16074 9509
rect 16016 9469 16028 9503
rect 16062 9500 16074 9503
rect 17678 9500 17684 9512
rect 16062 9472 17684 9500
rect 16062 9469 16074 9472
rect 16016 9463 16074 9469
rect 10060 9404 10272 9432
rect 10404 9435 10462 9441
rect 10404 9401 10416 9435
rect 10450 9432 10462 9435
rect 11146 9432 11152 9444
rect 10450 9404 11152 9432
rect 10450 9401 10462 9404
rect 10404 9395 10462 9401
rect 11146 9392 11152 9404
rect 11204 9392 11210 9444
rect 15764 9432 15792 9463
rect 17678 9460 17684 9472
rect 17736 9460 17742 9512
rect 18325 9503 18383 9509
rect 18325 9469 18337 9503
rect 18371 9500 18383 9503
rect 18782 9500 18788 9512
rect 18371 9472 18788 9500
rect 18371 9469 18383 9472
rect 18325 9463 18383 9469
rect 18782 9460 18788 9472
rect 18840 9460 18846 9512
rect 19426 9500 19432 9512
rect 19387 9472 19432 9500
rect 19426 9460 19432 9472
rect 19484 9460 19490 9512
rect 19696 9503 19754 9509
rect 19696 9469 19708 9503
rect 19742 9500 19754 9503
rect 20622 9500 20628 9512
rect 19742 9472 20628 9500
rect 19742 9469 19754 9472
rect 19696 9463 19754 9469
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 16298 9432 16304 9444
rect 15764 9404 16304 9432
rect 16298 9392 16304 9404
rect 16356 9392 16362 9444
rect 16666 9392 16672 9444
rect 16724 9432 16730 9444
rect 16724 9404 18552 9432
rect 16724 9392 16730 9404
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 11974 9364 11980 9376
rect 11112 9336 11980 9364
rect 11112 9324 11118 9336
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 12250 9324 12256 9376
rect 12308 9364 12314 9376
rect 12618 9364 12624 9376
rect 12308 9336 12624 9364
rect 12308 9324 12314 9336
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 14274 9324 14280 9376
rect 14332 9364 14338 9376
rect 14921 9367 14979 9373
rect 14921 9364 14933 9367
rect 14332 9336 14933 9364
rect 14332 9324 14338 9336
rect 14921 9333 14933 9336
rect 14967 9333 14979 9367
rect 17126 9364 17132 9376
rect 17087 9336 17132 9364
rect 14921 9327 14979 9333
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 18524 9373 18552 9404
rect 18509 9367 18567 9373
rect 18509 9333 18521 9367
rect 18555 9333 18567 9367
rect 18509 9327 18567 9333
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 8021 9163 8079 9169
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 8478 9160 8484 9172
rect 8067 9132 8484 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 9766 9160 9772 9172
rect 9727 9132 9772 9160
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 11238 9120 11244 9172
rect 11296 9160 11302 9172
rect 11333 9163 11391 9169
rect 11333 9160 11345 9163
rect 11296 9132 11345 9160
rect 11296 9120 11302 9132
rect 11333 9129 11345 9132
rect 11379 9129 11391 9163
rect 11333 9123 11391 9129
rect 11790 9120 11796 9172
rect 11848 9160 11854 9172
rect 13633 9163 13691 9169
rect 13633 9160 13645 9163
rect 11848 9132 13645 9160
rect 11848 9120 11854 9132
rect 13633 9129 13645 9132
rect 13679 9129 13691 9163
rect 13633 9123 13691 9129
rect 14093 9163 14151 9169
rect 14093 9129 14105 9163
rect 14139 9160 14151 9163
rect 16942 9160 16948 9172
rect 14139 9132 16948 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 16942 9120 16948 9132
rect 17000 9160 17006 9172
rect 19242 9160 19248 9172
rect 17000 9132 17264 9160
rect 19203 9132 19248 9160
rect 17000 9120 17006 9132
rect 8496 9064 11836 9092
rect 6546 8984 6552 9036
rect 6604 9024 6610 9036
rect 8496 9033 8524 9064
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 6604 8996 8401 9024
rect 6604 8984 6610 8996
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 8389 8987 8447 8993
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 8993 8539 9027
rect 10134 9024 10140 9036
rect 10095 8996 10140 9024
rect 8481 8987 8539 8993
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 11808 9033 11836 9064
rect 12066 9052 12072 9104
rect 12124 9092 12130 9104
rect 14001 9095 14059 9101
rect 14001 9092 14013 9095
rect 12124 9064 14013 9092
rect 12124 9052 12130 9064
rect 14001 9061 14013 9064
rect 14047 9061 14059 9095
rect 14001 9055 14059 9061
rect 16844 9095 16902 9101
rect 16844 9061 16856 9095
rect 16890 9092 16902 9095
rect 17126 9092 17132 9104
rect 16890 9064 17132 9092
rect 16890 9061 16902 9064
rect 16844 9055 16902 9061
rect 17126 9052 17132 9064
rect 17184 9052 17190 9104
rect 17236 9092 17264 9132
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 17236 9064 19288 9092
rect 19260 9036 19288 9064
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 10336 8996 11713 9024
rect 7006 8956 7012 8968
rect 6967 8928 7012 8956
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 10226 8956 10232 8968
rect 8628 8928 8673 8956
rect 10187 8928 10232 8956
rect 8628 8916 8634 8928
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 7282 8848 7288 8900
rect 7340 8888 7346 8900
rect 10336 8888 10364 8996
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 11701 8987 11759 8993
rect 11793 9027 11851 9033
rect 11793 8993 11805 9027
rect 11839 9024 11851 9027
rect 13446 9024 13452 9036
rect 11839 8996 13452 9024
rect 11839 8993 11851 8996
rect 11793 8987 11851 8993
rect 13446 8984 13452 8996
rect 13504 8984 13510 9036
rect 15286 9024 15292 9036
rect 15247 8996 15292 9024
rect 15286 8984 15292 8996
rect 15344 8984 15350 9036
rect 16390 8984 16396 9036
rect 16448 9024 16454 9036
rect 18874 9024 18880 9036
rect 16448 8996 18880 9024
rect 16448 8984 16454 8996
rect 18874 8984 18880 8996
rect 18932 9024 18938 9036
rect 19153 9027 19211 9033
rect 19153 9024 19165 9027
rect 18932 8996 19165 9024
rect 18932 8984 18938 8996
rect 19153 8993 19165 8996
rect 19199 8993 19211 9027
rect 19153 8987 19211 8993
rect 19242 8984 19248 9036
rect 19300 8984 19306 9036
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8956 10471 8959
rect 11054 8956 11060 8968
rect 10459 8928 11060 8956
rect 10459 8925 10471 8928
rect 10413 8919 10471 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8925 11943 8959
rect 11885 8919 11943 8925
rect 7340 8860 10364 8888
rect 7340 8848 7346 8860
rect 11146 8848 11152 8900
rect 11204 8888 11210 8900
rect 11900 8888 11928 8919
rect 11974 8916 11980 8968
rect 12032 8956 12038 8968
rect 13722 8956 13728 8968
rect 12032 8928 13728 8956
rect 12032 8916 12038 8928
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 14274 8956 14280 8968
rect 14235 8928 14280 8956
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 15473 8959 15531 8965
rect 15473 8925 15485 8959
rect 15519 8925 15531 8959
rect 15473 8919 15531 8925
rect 11204 8860 11928 8888
rect 11204 8848 11210 8860
rect 12802 8848 12808 8900
rect 12860 8888 12866 8900
rect 15488 8888 15516 8919
rect 15746 8916 15752 8968
rect 15804 8956 15810 8968
rect 16482 8956 16488 8968
rect 15804 8928 16488 8956
rect 15804 8916 15810 8928
rect 16482 8916 16488 8928
rect 16540 8956 16546 8968
rect 16577 8959 16635 8965
rect 16577 8956 16589 8959
rect 16540 8928 16589 8956
rect 16540 8916 16546 8928
rect 16577 8925 16589 8928
rect 16623 8925 16635 8959
rect 19058 8956 19064 8968
rect 16577 8919 16635 8925
rect 17880 8928 19064 8956
rect 12860 8860 15516 8888
rect 12860 8848 12866 8860
rect 4338 8780 4344 8832
rect 4396 8820 4402 8832
rect 12066 8820 12072 8832
rect 4396 8792 12072 8820
rect 4396 8780 4402 8792
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 17880 8820 17908 8928
rect 19058 8916 19064 8928
rect 19116 8916 19122 8968
rect 19337 8959 19395 8965
rect 19337 8925 19349 8959
rect 19383 8925 19395 8959
rect 19337 8919 19395 8925
rect 17957 8891 18015 8897
rect 17957 8857 17969 8891
rect 18003 8888 18015 8891
rect 18138 8888 18144 8900
rect 18003 8860 18144 8888
rect 18003 8857 18015 8860
rect 17957 8851 18015 8857
rect 18138 8848 18144 8860
rect 18196 8888 18202 8900
rect 19352 8888 19380 8919
rect 18196 8860 19380 8888
rect 18196 8848 18202 8860
rect 12676 8792 17908 8820
rect 18785 8823 18843 8829
rect 12676 8780 12682 8792
rect 18785 8789 18797 8823
rect 18831 8820 18843 8823
rect 18874 8820 18880 8832
rect 18831 8792 18880 8820
rect 18831 8789 18843 8792
rect 18785 8783 18843 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 7282 8616 7288 8628
rect 2372 8588 7288 8616
rect 2372 8576 2378 8588
rect 7282 8576 7288 8588
rect 7340 8576 7346 8628
rect 8389 8619 8447 8625
rect 8389 8585 8401 8619
rect 8435 8616 8447 8619
rect 8570 8616 8576 8628
rect 8435 8588 8576 8616
rect 8435 8585 8447 8588
rect 8389 8579 8447 8585
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 11204 8588 11253 8616
rect 11204 8576 11210 8588
rect 11241 8585 11253 8588
rect 11287 8585 11299 8619
rect 12618 8616 12624 8628
rect 12579 8588 12624 8616
rect 11241 8579 11299 8585
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 13722 8576 13728 8628
rect 13780 8616 13786 8628
rect 14921 8619 14979 8625
rect 14921 8616 14933 8619
rect 13780 8588 14933 8616
rect 13780 8576 13786 8588
rect 14921 8585 14933 8588
rect 14967 8585 14979 8619
rect 14921 8579 14979 8585
rect 15286 8576 15292 8628
rect 15344 8616 15350 8628
rect 16117 8619 16175 8625
rect 16117 8616 16129 8619
rect 15344 8588 16129 8616
rect 15344 8576 15350 8588
rect 16117 8585 16129 8588
rect 16163 8585 16175 8619
rect 16117 8579 16175 8585
rect 16758 8576 16764 8628
rect 16816 8616 16822 8628
rect 18233 8619 18291 8625
rect 18233 8616 18245 8619
rect 16816 8588 18245 8616
rect 16816 8576 16822 8588
rect 18233 8585 18245 8588
rect 18279 8585 18291 8619
rect 19426 8616 19432 8628
rect 18233 8579 18291 8585
rect 19168 8588 19432 8616
rect 16482 8508 16488 8560
rect 16540 8548 16546 8560
rect 19168 8548 19196 8588
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 16540 8520 19196 8548
rect 16540 8508 16546 8520
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 9272 8452 9873 8480
rect 9272 8440 9278 8452
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 13538 8480 13544 8492
rect 13499 8452 13544 8480
rect 9861 8443 9919 8449
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 16761 8483 16819 8489
rect 16761 8449 16773 8483
rect 16807 8480 16819 8483
rect 17126 8480 17132 8492
rect 16807 8452 17132 8480
rect 16807 8449 16819 8452
rect 16761 8443 16819 8449
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 19168 8489 19196 8520
rect 19153 8483 19211 8489
rect 19153 8449 19165 8483
rect 19199 8449 19211 8483
rect 19153 8443 19211 8449
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 9232 8412 9260 8440
rect 7055 8384 9260 8412
rect 12437 8415 12495 8421
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 12437 8381 12449 8415
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 13808 8415 13866 8421
rect 13808 8381 13820 8415
rect 13854 8412 13866 8415
rect 14274 8412 14280 8424
rect 13854 8384 14280 8412
rect 13854 8381 13866 8384
rect 13808 8375 13866 8381
rect 7024 8344 7052 8375
rect 6840 8316 7052 8344
rect 7276 8347 7334 8353
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 6840 8276 6868 8316
rect 7276 8313 7288 8347
rect 7322 8344 7334 8347
rect 7742 8344 7748 8356
rect 7322 8316 7748 8344
rect 7322 8313 7334 8316
rect 7276 8307 7334 8313
rect 7742 8304 7748 8316
rect 7800 8304 7806 8356
rect 10128 8347 10186 8353
rect 10128 8313 10140 8347
rect 10174 8344 10186 8347
rect 11054 8344 11060 8356
rect 10174 8316 11060 8344
rect 10174 8313 10186 8316
rect 10128 8307 10186 8313
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 12452 8344 12480 8375
rect 14274 8372 14280 8384
rect 14332 8372 14338 8424
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8412 15991 8415
rect 16114 8412 16120 8424
rect 15979 8384 16120 8412
rect 15979 8381 15991 8384
rect 15933 8375 15991 8381
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 16206 8372 16212 8424
rect 16264 8412 16270 8424
rect 16485 8415 16543 8421
rect 16485 8412 16497 8415
rect 16264 8384 16497 8412
rect 16264 8372 16270 8384
rect 16485 8381 16497 8384
rect 16531 8381 16543 8415
rect 16485 8375 16543 8381
rect 16577 8415 16635 8421
rect 16577 8381 16589 8415
rect 16623 8412 16635 8415
rect 17770 8412 17776 8424
rect 16623 8384 17776 8412
rect 16623 8381 16635 8384
rect 16577 8375 16635 8381
rect 17770 8372 17776 8384
rect 17828 8372 17834 8424
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8412 18107 8415
rect 18690 8412 18696 8424
rect 18095 8384 18696 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18690 8372 18696 8384
rect 18748 8372 18754 8424
rect 18598 8344 18604 8356
rect 12452 8316 18604 8344
rect 18598 8304 18604 8316
rect 18656 8304 18662 8356
rect 19334 8304 19340 8356
rect 19392 8353 19398 8356
rect 19392 8347 19456 8353
rect 19392 8313 19410 8347
rect 19444 8313 19456 8347
rect 19392 8307 19456 8313
rect 19392 8304 19398 8307
rect 6696 8248 6868 8276
rect 6696 8236 6702 8248
rect 13538 8236 13544 8288
rect 13596 8276 13602 8288
rect 15746 8276 15752 8288
rect 13596 8248 15752 8276
rect 13596 8236 13602 8248
rect 15746 8236 15752 8248
rect 15804 8236 15810 8288
rect 20530 8276 20536 8288
rect 20491 8248 20536 8276
rect 20530 8236 20536 8248
rect 20588 8236 20594 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 7800 8044 8033 8072
rect 7800 8032 7806 8044
rect 8021 8041 8033 8044
rect 8067 8041 8079 8075
rect 11054 8072 11060 8084
rect 11015 8044 11060 8072
rect 8021 8035 8079 8041
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 16390 8072 16396 8084
rect 11900 8044 16396 8072
rect 5629 8007 5687 8013
rect 5629 7973 5641 8007
rect 5675 8004 5687 8007
rect 10134 8004 10140 8016
rect 5675 7976 10140 8004
rect 5675 7973 5687 7976
rect 5629 7967 5687 7973
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 10318 7964 10324 8016
rect 10376 8004 10382 8016
rect 11900 8004 11928 8044
rect 16390 8032 16396 8044
rect 16448 8072 16454 8084
rect 16669 8075 16727 8081
rect 16669 8072 16681 8075
rect 16448 8044 16681 8072
rect 16448 8032 16454 8044
rect 16669 8041 16681 8044
rect 16715 8041 16727 8075
rect 16669 8035 16727 8041
rect 16761 8075 16819 8081
rect 16761 8041 16773 8075
rect 16807 8072 16819 8075
rect 18046 8072 18052 8084
rect 16807 8044 18052 8072
rect 16807 8041 16819 8044
rect 16761 8035 16819 8041
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 10376 7976 11928 8004
rect 10376 7964 10382 7976
rect 11974 7964 11980 8016
rect 12032 8004 12038 8016
rect 12130 8007 12188 8013
rect 12130 8004 12142 8007
rect 12032 7976 12142 8004
rect 12032 7964 12038 7976
rect 12130 7973 12142 7976
rect 12176 7973 12188 8007
rect 12130 7967 12188 7973
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 16850 8004 16856 8016
rect 12768 7976 16856 8004
rect 12768 7964 12774 7976
rect 16850 7964 16856 7976
rect 16908 7964 16914 8016
rect 18138 8013 18144 8016
rect 18132 8004 18144 8013
rect 18099 7976 18144 8004
rect 18132 7967 18144 7976
rect 18138 7964 18144 7967
rect 18196 7964 18202 8016
rect 6638 7936 6644 7948
rect 6599 7908 6644 7936
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 6908 7939 6966 7945
rect 6908 7905 6920 7939
rect 6954 7936 6966 7939
rect 7466 7936 7472 7948
rect 6954 7908 7472 7936
rect 6954 7905 6966 7908
rect 6908 7899 6966 7905
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 9214 7896 9220 7948
rect 9272 7936 9278 7948
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 9272 7908 9689 7936
rect 9272 7896 9278 7908
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 9944 7939 10002 7945
rect 9944 7905 9956 7939
rect 9990 7936 10002 7939
rect 10410 7936 10416 7948
rect 9990 7908 10416 7936
rect 9990 7905 10002 7908
rect 9944 7899 10002 7905
rect 10410 7896 10416 7908
rect 10468 7896 10474 7948
rect 14093 7939 14151 7945
rect 14093 7905 14105 7939
rect 14139 7936 14151 7939
rect 20530 7936 20536 7948
rect 14139 7908 16528 7936
rect 14139 7905 14151 7908
rect 14093 7899 14151 7905
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7837 11943 7871
rect 11885 7831 11943 7837
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7868 15347 7871
rect 15838 7868 15844 7880
rect 15335 7840 15844 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 11900 7732 11928 7831
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 12894 7732 12900 7744
rect 11900 7704 12900 7732
rect 12894 7692 12900 7704
rect 12952 7692 12958 7744
rect 13262 7732 13268 7744
rect 13223 7704 13268 7732
rect 13262 7692 13268 7704
rect 13320 7692 13326 7744
rect 14277 7735 14335 7741
rect 14277 7701 14289 7735
rect 14323 7732 14335 7735
rect 16114 7732 16120 7744
rect 14323 7704 16120 7732
rect 14323 7701 14335 7704
rect 14277 7695 14335 7701
rect 16114 7692 16120 7704
rect 16172 7692 16178 7744
rect 16298 7732 16304 7744
rect 16259 7704 16304 7732
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 16500 7732 16528 7908
rect 16960 7908 20536 7936
rect 16960 7877 16988 7908
rect 20530 7896 20536 7908
rect 20588 7896 20594 7948
rect 16945 7871 17003 7877
rect 16945 7837 16957 7871
rect 16991 7837 17003 7871
rect 16945 7831 17003 7837
rect 17865 7871 17923 7877
rect 17865 7837 17877 7871
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 16574 7760 16580 7812
rect 16632 7800 16638 7812
rect 17770 7800 17776 7812
rect 16632 7772 17776 7800
rect 16632 7760 16638 7772
rect 17770 7760 17776 7772
rect 17828 7800 17834 7812
rect 17880 7800 17908 7831
rect 17828 7772 17908 7800
rect 17828 7760 17834 7772
rect 18138 7732 18144 7744
rect 16500 7704 18144 7732
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 19245 7735 19303 7741
rect 19245 7701 19257 7735
rect 19291 7732 19303 7735
rect 19334 7732 19340 7744
rect 19291 7704 19340 7732
rect 19291 7701 19303 7704
rect 19245 7695 19303 7701
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 7098 7528 7104 7540
rect 7059 7500 7104 7528
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 9306 7488 9312 7540
rect 9364 7528 9370 7540
rect 9401 7531 9459 7537
rect 9401 7528 9413 7531
rect 9364 7500 9413 7528
rect 9364 7488 9370 7500
rect 9401 7497 9413 7500
rect 9447 7497 9459 7531
rect 9401 7491 9459 7497
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 10226 7528 10232 7540
rect 9640 7500 10232 7528
rect 9640 7488 9646 7500
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 10965 7531 11023 7537
rect 10965 7497 10977 7531
rect 11011 7528 11023 7531
rect 18690 7528 18696 7540
rect 11011 7500 18696 7528
rect 11011 7497 11023 7500
rect 10965 7491 11023 7497
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 20162 7488 20168 7540
rect 20220 7528 20226 7540
rect 20220 7500 20392 7528
rect 20220 7488 20226 7500
rect 16393 7463 16451 7469
rect 16393 7429 16405 7463
rect 16439 7460 16451 7463
rect 20364 7460 20392 7500
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 22094 7528 22100 7540
rect 20772 7500 22100 7528
rect 20772 7488 20778 7500
rect 22094 7488 22100 7500
rect 22152 7488 22158 7540
rect 20809 7463 20867 7469
rect 20809 7460 20821 7463
rect 16439 7432 18092 7460
rect 20364 7432 20821 7460
rect 16439 7429 16451 7432
rect 16393 7423 16451 7429
rect 5810 7352 5816 7404
rect 5868 7392 5874 7404
rect 7742 7392 7748 7404
rect 5868 7364 7604 7392
rect 7703 7364 7748 7392
rect 5868 7352 5874 7364
rect 7006 7284 7012 7336
rect 7064 7324 7070 7336
rect 7469 7327 7527 7333
rect 7469 7324 7481 7327
rect 7064 7296 7481 7324
rect 7064 7284 7070 7296
rect 7469 7293 7481 7296
rect 7515 7293 7527 7327
rect 7576 7324 7604 7364
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 10045 7395 10103 7401
rect 10045 7361 10057 7395
rect 10091 7392 10103 7395
rect 10410 7392 10416 7404
rect 10091 7364 10416 7392
rect 10091 7361 10103 7364
rect 10045 7355 10103 7361
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13262 7392 13268 7404
rect 13127 7364 13268 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 13596 7364 14013 7392
rect 13596 7352 13602 7364
rect 14001 7361 14013 7364
rect 14047 7361 14059 7395
rect 17034 7392 17040 7404
rect 16995 7364 17040 7392
rect 14001 7355 14059 7361
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 10778 7324 10784 7336
rect 7576 7296 10784 7324
rect 7469 7287 7527 7293
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 11057 7327 11115 7333
rect 11057 7293 11069 7327
rect 11103 7324 11115 7327
rect 12710 7324 12716 7336
rect 11103 7296 12716 7324
rect 11103 7293 11115 7296
rect 11057 7287 11115 7293
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 12897 7327 12955 7333
rect 12897 7293 12909 7327
rect 12943 7324 12955 7327
rect 16206 7324 16212 7336
rect 12943 7296 16212 7324
rect 12943 7293 12955 7296
rect 12897 7287 12955 7293
rect 7374 7216 7380 7268
rect 7432 7256 7438 7268
rect 10965 7259 11023 7265
rect 10965 7256 10977 7259
rect 7432 7228 10977 7256
rect 7432 7216 7438 7228
rect 10965 7225 10977 7228
rect 11011 7225 11023 7259
rect 10965 7219 11023 7225
rect 11146 7216 11152 7268
rect 11204 7256 11210 7268
rect 11333 7259 11391 7265
rect 11333 7256 11345 7259
rect 11204 7228 11345 7256
rect 11204 7216 11210 7228
rect 11333 7225 11345 7228
rect 11379 7225 11391 7259
rect 11333 7219 11391 7225
rect 11974 7216 11980 7268
rect 12032 7256 12038 7268
rect 12912 7256 12940 7287
rect 16206 7284 16212 7296
rect 16264 7324 16270 7336
rect 17954 7324 17960 7336
rect 16264 7296 17960 7324
rect 16264 7284 16270 7296
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 18064 7333 18092 7432
rect 20809 7429 20821 7432
rect 20855 7429 20867 7463
rect 20809 7423 20867 7429
rect 19426 7392 19432 7404
rect 19387 7364 19432 7392
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 19696 7327 19754 7333
rect 19696 7293 19708 7327
rect 19742 7324 19754 7327
rect 20530 7324 20536 7336
rect 19742 7296 20536 7324
rect 19742 7293 19754 7296
rect 19696 7287 19754 7293
rect 20530 7284 20536 7296
rect 20588 7284 20594 7336
rect 12032 7228 12940 7256
rect 14268 7259 14326 7265
rect 12032 7216 12038 7228
rect 14268 7225 14280 7259
rect 14314 7256 14326 7259
rect 14366 7256 14372 7268
rect 14314 7228 14372 7256
rect 14314 7225 14326 7228
rect 14268 7219 14326 7225
rect 14366 7216 14372 7228
rect 14424 7216 14430 7268
rect 16574 7216 16580 7268
rect 16632 7256 16638 7268
rect 16853 7259 16911 7265
rect 16853 7256 16865 7259
rect 16632 7228 16865 7256
rect 16632 7216 16638 7228
rect 16853 7225 16865 7228
rect 16899 7225 16911 7259
rect 16853 7219 16911 7225
rect 18325 7259 18383 7265
rect 18325 7225 18337 7259
rect 18371 7225 18383 7259
rect 18325 7219 18383 7225
rect 7558 7188 7564 7200
rect 7519 7160 7564 7188
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 9766 7188 9772 7200
rect 9727 7160 9772 7188
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 12437 7191 12495 7197
rect 9916 7160 9961 7188
rect 9916 7148 9922 7160
rect 12437 7157 12449 7191
rect 12483 7188 12495 7191
rect 12526 7188 12532 7200
rect 12483 7160 12532 7188
rect 12483 7157 12495 7160
rect 12437 7151 12495 7157
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 12805 7191 12863 7197
rect 12805 7157 12817 7191
rect 12851 7188 12863 7191
rect 14090 7188 14096 7200
rect 12851 7160 14096 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 15378 7188 15384 7200
rect 15339 7160 15384 7188
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 15930 7148 15936 7200
rect 15988 7188 15994 7200
rect 16761 7191 16819 7197
rect 16761 7188 16773 7191
rect 15988 7160 16773 7188
rect 15988 7148 15994 7160
rect 16761 7157 16773 7160
rect 16807 7157 16819 7191
rect 16761 7151 16819 7157
rect 17402 7148 17408 7200
rect 17460 7188 17466 7200
rect 18340 7188 18368 7219
rect 17460 7160 18368 7188
rect 17460 7148 17466 7160
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 7285 6987 7343 6993
rect 7285 6953 7297 6987
rect 7331 6984 7343 6987
rect 7558 6984 7564 6996
rect 7331 6956 7564 6984
rect 7331 6953 7343 6956
rect 7285 6947 7343 6953
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 12069 6987 12127 6993
rect 12069 6953 12081 6987
rect 12115 6984 12127 6987
rect 12250 6984 12256 6996
rect 12115 6956 12256 6984
rect 12115 6953 12127 6956
rect 12069 6947 12127 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12526 6984 12532 6996
rect 12487 6956 12532 6984
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 15657 6987 15715 6993
rect 15657 6953 15669 6987
rect 15703 6984 15715 6987
rect 16853 6987 16911 6993
rect 16853 6984 16865 6987
rect 15703 6956 16865 6984
rect 15703 6953 15715 6956
rect 15657 6947 15715 6953
rect 16853 6953 16865 6956
rect 16899 6953 16911 6987
rect 17218 6984 17224 6996
rect 17179 6956 17224 6984
rect 16853 6947 16911 6953
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 18785 6987 18843 6993
rect 18785 6953 18797 6987
rect 18831 6984 18843 6987
rect 19150 6984 19156 6996
rect 18831 6956 19156 6984
rect 18831 6953 18843 6956
rect 18785 6947 18843 6953
rect 19150 6944 19156 6956
rect 19208 6944 19214 6996
rect 7098 6876 7104 6928
rect 7156 6916 7162 6928
rect 7653 6919 7711 6925
rect 7653 6916 7665 6919
rect 7156 6888 7665 6916
rect 7156 6876 7162 6888
rect 7653 6885 7665 6888
rect 7699 6885 7711 6919
rect 7653 6879 7711 6885
rect 12434 6876 12440 6928
rect 12492 6916 12498 6928
rect 13998 6916 14004 6928
rect 12492 6888 12537 6916
rect 13959 6888 14004 6916
rect 12492 6876 12498 6888
rect 13998 6876 14004 6888
rect 14056 6876 14062 6928
rect 15470 6876 15476 6928
rect 15528 6916 15534 6928
rect 15749 6919 15807 6925
rect 15749 6916 15761 6919
rect 15528 6888 15761 6916
rect 15528 6876 15534 6888
rect 15749 6885 15761 6888
rect 15795 6885 15807 6919
rect 15749 6879 15807 6885
rect 16298 6876 16304 6928
rect 16356 6916 16362 6928
rect 20070 6916 20076 6928
rect 16356 6888 20076 6916
rect 16356 6876 16362 6888
rect 20070 6876 20076 6888
rect 20128 6876 20134 6928
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 10042 6848 10048 6860
rect 7524 6820 7880 6848
rect 10003 6820 10048 6848
rect 7524 6808 7530 6820
rect 7852 6789 7880 6820
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 11977 6851 12035 6857
rect 11977 6817 11989 6851
rect 12023 6848 12035 6851
rect 12158 6848 12164 6860
rect 12023 6820 12164 6848
rect 12023 6817 12035 6820
rect 11977 6811 12035 6817
rect 12158 6808 12164 6820
rect 12216 6808 12222 6860
rect 14093 6851 14151 6857
rect 14093 6817 14105 6851
rect 14139 6848 14151 6851
rect 17310 6848 17316 6860
rect 14139 6820 17080 6848
rect 17271 6820 17316 6848
rect 14139 6817 14151 6820
rect 14093 6811 14151 6817
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6780 7895 6783
rect 8202 6780 8208 6792
rect 7883 6752 8208 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 7760 6712 7788 6743
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 9858 6780 9864 6792
rect 8312 6752 9864 6780
rect 8312 6712 8340 6752
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10318 6780 10324 6792
rect 10279 6752 10324 6780
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 12710 6780 12716 6792
rect 11112 6752 12716 6780
rect 11112 6740 11118 6752
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 7760 6684 8340 6712
rect 9677 6715 9735 6721
rect 9677 6681 9689 6715
rect 9723 6712 9735 6715
rect 9950 6712 9956 6724
rect 9723 6684 9956 6712
rect 9723 6681 9735 6684
rect 9677 6675 9735 6681
rect 9950 6672 9956 6684
rect 10008 6672 10014 6724
rect 13630 6712 13636 6724
rect 10060 6684 13492 6712
rect 13591 6684 13636 6712
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 10060 6644 10088 6684
rect 5776 6616 10088 6644
rect 5776 6604 5782 6616
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 11790 6644 11796 6656
rect 10836 6616 11796 6644
rect 10836 6604 10842 6616
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 13464 6644 13492 6684
rect 13630 6672 13636 6684
rect 13688 6672 13694 6724
rect 14292 6712 14320 6743
rect 15378 6740 15384 6792
rect 15436 6780 15442 6792
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15436 6752 15853 6780
rect 15436 6740 15442 6752
rect 15841 6749 15853 6752
rect 15887 6780 15899 6783
rect 16022 6780 16028 6792
rect 15887 6752 16028 6780
rect 15887 6749 15899 6752
rect 15841 6743 15899 6749
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 17052 6780 17080 6820
rect 17310 6808 17316 6820
rect 17368 6808 17374 6860
rect 18874 6808 18880 6860
rect 18932 6848 18938 6860
rect 18932 6820 18977 6848
rect 18932 6808 18938 6820
rect 17402 6780 17408 6792
rect 17052 6752 17264 6780
rect 17363 6752 17408 6780
rect 17126 6712 17132 6724
rect 14292 6684 17132 6712
rect 17126 6672 17132 6684
rect 17184 6672 17190 6724
rect 17236 6712 17264 6752
rect 17402 6740 17408 6752
rect 17460 6740 17466 6792
rect 19061 6783 19119 6789
rect 19061 6749 19073 6783
rect 19107 6780 19119 6783
rect 19334 6780 19340 6792
rect 19107 6752 19340 6780
rect 19107 6749 19119 6752
rect 19061 6743 19119 6749
rect 19334 6740 19340 6752
rect 19392 6740 19398 6792
rect 19610 6712 19616 6724
rect 17236 6684 19616 6712
rect 19610 6672 19616 6684
rect 19668 6672 19674 6724
rect 15194 6644 15200 6656
rect 13464 6616 15200 6644
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 15289 6647 15347 6653
rect 15289 6613 15301 6647
rect 15335 6644 15347 6647
rect 16574 6644 16580 6656
rect 15335 6616 16580 6644
rect 15335 6613 15347 6616
rect 15289 6607 15347 6613
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 16850 6604 16856 6656
rect 16908 6644 16914 6656
rect 18417 6647 18475 6653
rect 18417 6644 18429 6647
rect 16908 6616 18429 6644
rect 16908 6604 16914 6616
rect 18417 6613 18429 6616
rect 18463 6613 18475 6647
rect 18417 6607 18475 6613
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 8202 6440 8208 6452
rect 8163 6412 8208 6440
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 10410 6440 10416 6452
rect 10371 6412 10416 6440
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 12618 6440 12624 6452
rect 11256 6412 12624 6440
rect 5718 6304 5724 6316
rect 5679 6276 5724 6304
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6696 6276 6837 6304
rect 6696 6264 6702 6276
rect 6825 6273 6837 6276
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6236 9091 6239
rect 10778 6236 10784 6248
rect 9079 6208 10784 6236
rect 9079 6205 9091 6208
rect 9033 6199 9091 6205
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 11256 6245 11284 6412
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 13817 6443 13875 6449
rect 13817 6440 13829 6443
rect 12768 6412 13829 6440
rect 12768 6400 12774 6412
rect 13817 6409 13829 6412
rect 13863 6409 13875 6443
rect 13817 6403 13875 6409
rect 13906 6400 13912 6452
rect 13964 6440 13970 6452
rect 16942 6440 16948 6452
rect 13964 6412 16948 6440
rect 13964 6400 13970 6412
rect 16942 6400 16948 6412
rect 17000 6400 17006 6452
rect 17034 6400 17040 6452
rect 17092 6440 17098 6452
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 17092 6412 17141 6440
rect 17092 6400 17098 6412
rect 17129 6409 17141 6412
rect 17175 6440 17187 6443
rect 17678 6440 17684 6452
rect 17175 6412 17684 6440
rect 17175 6409 17187 6412
rect 17129 6403 17187 6409
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 11425 6375 11483 6381
rect 11425 6341 11437 6375
rect 11471 6372 11483 6375
rect 12158 6372 12164 6384
rect 11471 6344 12164 6372
rect 11471 6341 11483 6344
rect 11425 6335 11483 6341
rect 12158 6332 12164 6344
rect 12216 6332 12222 6384
rect 15746 6304 15752 6316
rect 15707 6276 15752 6304
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 17678 6264 17684 6316
rect 17736 6304 17742 6316
rect 17736 6276 18184 6304
rect 17736 6264 17742 6276
rect 11241 6239 11299 6245
rect 11241 6205 11253 6239
rect 11287 6205 11299 6239
rect 11241 6199 11299 6205
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 12704 6239 12762 6245
rect 12483 6208 12517 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 12704 6205 12716 6239
rect 12750 6236 12762 6239
rect 13262 6236 13268 6248
rect 12750 6208 13268 6236
rect 12750 6205 12762 6208
rect 12704 6199 12762 6205
rect 7092 6171 7150 6177
rect 7092 6137 7104 6171
rect 7138 6168 7150 6171
rect 7742 6168 7748 6180
rect 7138 6140 7748 6168
rect 7138 6137 7150 6140
rect 7092 6131 7150 6137
rect 7742 6128 7748 6140
rect 7800 6128 7806 6180
rect 9300 6171 9358 6177
rect 9300 6137 9312 6171
rect 9346 6168 9358 6171
rect 10318 6168 10324 6180
rect 9346 6140 10324 6168
rect 9346 6137 9358 6140
rect 9300 6131 9358 6137
rect 10318 6128 10324 6140
rect 10376 6128 10382 6180
rect 11790 6128 11796 6180
rect 11848 6168 11854 6180
rect 12452 6168 12480 6199
rect 13262 6196 13268 6208
rect 13320 6196 13326 6248
rect 16022 6245 16028 6248
rect 14645 6239 14703 6245
rect 14645 6205 14657 6239
rect 14691 6205 14703 6239
rect 16016 6236 16028 6245
rect 15983 6208 16028 6236
rect 14645 6199 14703 6205
rect 16016 6199 16028 6208
rect 12894 6168 12900 6180
rect 11848 6140 12900 6168
rect 11848 6128 11854 6140
rect 12894 6128 12900 6140
rect 12952 6128 12958 6180
rect 14660 6168 14688 6199
rect 16022 6196 16028 6199
rect 16080 6196 16086 6248
rect 17034 6196 17040 6248
rect 17092 6236 17098 6248
rect 17218 6236 17224 6248
rect 17092 6208 17224 6236
rect 17092 6196 17098 6208
rect 17218 6196 17224 6208
rect 17276 6196 17282 6248
rect 17770 6196 17776 6248
rect 17828 6236 17834 6248
rect 18046 6236 18052 6248
rect 17828 6208 18052 6236
rect 17828 6196 17834 6208
rect 18046 6196 18052 6208
rect 18104 6196 18110 6248
rect 18156 6236 18184 6276
rect 18305 6239 18363 6245
rect 18305 6236 18317 6239
rect 18156 6208 18317 6236
rect 18305 6205 18317 6208
rect 18351 6205 18363 6239
rect 18305 6199 18363 6205
rect 20438 6196 20444 6248
rect 20496 6236 20502 6248
rect 20533 6239 20591 6245
rect 20533 6236 20545 6239
rect 20496 6208 20545 6236
rect 20496 6196 20502 6208
rect 20533 6205 20545 6208
rect 20579 6205 20591 6239
rect 20533 6199 20591 6205
rect 14660 6140 16436 6168
rect 12618 6060 12624 6112
rect 12676 6100 12682 6112
rect 13906 6100 13912 6112
rect 12676 6072 13912 6100
rect 12676 6060 12682 6072
rect 13906 6060 13912 6072
rect 13964 6060 13970 6112
rect 14829 6103 14887 6109
rect 14829 6069 14841 6103
rect 14875 6100 14887 6103
rect 15562 6100 15568 6112
rect 14875 6072 15568 6100
rect 14875 6069 14887 6072
rect 14829 6063 14887 6069
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 16408 6100 16436 6140
rect 16482 6128 16488 6180
rect 16540 6168 16546 6180
rect 17402 6168 17408 6180
rect 16540 6140 17408 6168
rect 16540 6128 16546 6140
rect 17402 6128 17408 6140
rect 17460 6128 17466 6180
rect 18782 6100 18788 6112
rect 16408 6072 18788 6100
rect 18782 6060 18788 6072
rect 18840 6060 18846 6112
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 19429 6103 19487 6109
rect 19429 6100 19441 6103
rect 19392 6072 19441 6100
rect 19392 6060 19398 6072
rect 19429 6069 19441 6072
rect 19475 6069 19487 6103
rect 19429 6063 19487 6069
rect 19702 6060 19708 6112
rect 19760 6100 19766 6112
rect 20717 6103 20775 6109
rect 20717 6100 20729 6103
rect 19760 6072 20729 6100
rect 19760 6060 19766 6072
rect 20717 6069 20729 6072
rect 20763 6069 20775 6103
rect 20717 6063 20775 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 7190 5896 7196 5908
rect 7151 5868 7196 5896
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 10042 5896 10048 5908
rect 8128 5868 10048 5896
rect 6181 5831 6239 5837
rect 6181 5797 6193 5831
rect 6227 5828 6239 5831
rect 8128 5828 8156 5868
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 10410 5856 10416 5908
rect 10468 5896 10474 5908
rect 14001 5899 14059 5905
rect 14001 5896 14013 5899
rect 10468 5868 14013 5896
rect 10468 5856 10474 5868
rect 14001 5865 14013 5868
rect 14047 5865 14059 5899
rect 14001 5859 14059 5865
rect 15289 5899 15347 5905
rect 15289 5865 15301 5899
rect 15335 5865 15347 5899
rect 15654 5896 15660 5908
rect 15567 5868 15660 5896
rect 15289 5859 15347 5865
rect 6227 5800 8156 5828
rect 6227 5797 6239 5800
rect 6181 5791 6239 5797
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7561 5763 7619 5769
rect 7561 5760 7573 5763
rect 6972 5732 7573 5760
rect 6972 5720 6978 5732
rect 7561 5729 7573 5732
rect 7607 5729 7619 5763
rect 7561 5723 7619 5729
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 10594 5760 10600 5772
rect 9723 5732 10600 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 10778 5760 10784 5772
rect 10739 5732 10784 5760
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 11054 5769 11060 5772
rect 11048 5760 11060 5769
rect 11015 5732 11060 5760
rect 11048 5723 11060 5732
rect 11054 5720 11060 5723
rect 11112 5720 11118 5772
rect 15304 5760 15332 5859
rect 15654 5856 15660 5868
rect 15712 5896 15718 5908
rect 18782 5896 18788 5908
rect 15712 5868 18788 5896
rect 15712 5856 15718 5868
rect 18782 5856 18788 5868
rect 18840 5856 18846 5908
rect 15470 5760 15476 5772
rect 15304 5732 15476 5760
rect 15470 5720 15476 5732
rect 15528 5720 15534 5772
rect 15749 5763 15807 5769
rect 15749 5729 15761 5763
rect 15795 5760 15807 5763
rect 16206 5760 16212 5772
rect 15795 5732 16212 5760
rect 15795 5729 15807 5732
rect 15749 5723 15807 5729
rect 16206 5720 16212 5732
rect 16264 5720 16270 5772
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 18408 5763 18466 5769
rect 16908 5732 16953 5760
rect 16908 5720 16914 5732
rect 18408 5729 18420 5763
rect 18454 5760 18466 5763
rect 19334 5760 19340 5772
rect 18454 5732 19340 5760
rect 18454 5729 18466 5732
rect 18408 5723 18466 5729
rect 19334 5720 19340 5732
rect 19392 5720 19398 5772
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5692 5227 5695
rect 6086 5692 6092 5704
rect 5215 5664 6092 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 7650 5692 7656 5704
rect 7611 5664 7656 5692
rect 7650 5652 7656 5664
rect 7708 5652 7714 5704
rect 7742 5652 7748 5704
rect 7800 5692 7806 5704
rect 14093 5695 14151 5701
rect 7800 5664 7845 5692
rect 7800 5652 7806 5664
rect 14093 5661 14105 5695
rect 14139 5692 14151 5695
rect 14182 5692 14188 5704
rect 14139 5664 14188 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5692 14335 5695
rect 14366 5692 14372 5704
rect 14323 5664 14372 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 14366 5652 14372 5664
rect 14424 5692 14430 5704
rect 15841 5695 15899 5701
rect 14424 5664 15415 5692
rect 14424 5652 14430 5664
rect 15387 5624 15415 5664
rect 15841 5661 15853 5695
rect 15887 5692 15899 5695
rect 16482 5692 16488 5704
rect 15887 5664 16488 5692
rect 15887 5661 15899 5664
rect 15841 5655 15899 5661
rect 15856 5624 15884 5655
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 17037 5695 17095 5701
rect 17037 5661 17049 5695
rect 17083 5661 17095 5695
rect 17037 5655 17095 5661
rect 15387 5596 15884 5624
rect 16666 5584 16672 5636
rect 16724 5624 16730 5636
rect 17052 5624 17080 5655
rect 18046 5652 18052 5704
rect 18104 5692 18110 5704
rect 18141 5695 18199 5701
rect 18141 5692 18153 5695
rect 18104 5664 18153 5692
rect 18104 5652 18110 5664
rect 18141 5661 18153 5664
rect 18187 5661 18199 5695
rect 18141 5655 18199 5661
rect 16724 5596 17080 5624
rect 16724 5584 16730 5596
rect 9858 5556 9864 5568
rect 9819 5528 9864 5556
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 11790 5516 11796 5568
rect 11848 5556 11854 5568
rect 12161 5559 12219 5565
rect 12161 5556 12173 5559
rect 11848 5528 12173 5556
rect 11848 5516 11854 5528
rect 12161 5525 12173 5528
rect 12207 5525 12219 5559
rect 12161 5519 12219 5525
rect 13633 5559 13691 5565
rect 13633 5525 13645 5559
rect 13679 5556 13691 5559
rect 14918 5556 14924 5568
rect 13679 5528 14924 5556
rect 13679 5525 13691 5528
rect 13633 5519 13691 5525
rect 14918 5516 14924 5528
rect 14976 5516 14982 5568
rect 19426 5516 19432 5568
rect 19484 5556 19490 5568
rect 19521 5559 19579 5565
rect 19521 5556 19533 5559
rect 19484 5528 19533 5556
rect 19484 5516 19490 5528
rect 19521 5525 19533 5528
rect 19567 5525 19579 5559
rect 19521 5519 19579 5525
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 7742 5312 7748 5364
rect 7800 5352 7806 5364
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 7800 5324 8217 5352
rect 7800 5312 7806 5324
rect 8205 5321 8217 5324
rect 8251 5321 8263 5355
rect 8205 5315 8263 5321
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 10597 5355 10655 5361
rect 10597 5352 10609 5355
rect 10376 5324 10609 5352
rect 10376 5312 10382 5324
rect 10597 5321 10609 5324
rect 10643 5321 10655 5355
rect 10597 5315 10655 5321
rect 10686 5312 10692 5364
rect 10744 5352 10750 5364
rect 11790 5352 11796 5364
rect 10744 5324 11796 5352
rect 10744 5312 10750 5324
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 15289 5355 15347 5361
rect 12492 5324 12537 5352
rect 12492 5312 12498 5324
rect 15289 5321 15301 5355
rect 15335 5352 15347 5355
rect 15930 5352 15936 5364
rect 15335 5324 15936 5352
rect 15335 5321 15347 5324
rect 15289 5315 15347 5321
rect 15930 5312 15936 5324
rect 15988 5312 15994 5364
rect 14550 5244 14556 5296
rect 14608 5284 14614 5296
rect 17037 5287 17095 5293
rect 17037 5284 17049 5287
rect 14608 5256 17049 5284
rect 14608 5244 14614 5256
rect 17037 5253 17049 5256
rect 17083 5253 17095 5287
rect 17037 5247 17095 5253
rect 18049 5287 18107 5293
rect 18049 5253 18061 5287
rect 18095 5284 18107 5287
rect 19886 5284 19892 5296
rect 18095 5256 19892 5284
rect 18095 5253 18107 5256
rect 18049 5247 18107 5253
rect 19886 5244 19892 5256
rect 19944 5244 19950 5296
rect 6638 5176 6644 5228
rect 6696 5216 6702 5228
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6696 5188 6837 5216
rect 6696 5176 6702 5188
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 9214 5216 9220 5228
rect 9175 5188 9220 5216
rect 6825 5179 6883 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5216 13139 5219
rect 13262 5216 13268 5228
rect 13127 5188 13268 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 14918 5176 14924 5228
rect 14976 5216 14982 5228
rect 15749 5219 15807 5225
rect 15749 5216 15761 5219
rect 14976 5188 15761 5216
rect 14976 5176 14982 5188
rect 15749 5185 15761 5188
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5216 15991 5219
rect 16022 5216 16028 5228
rect 15979 5188 16028 5216
rect 15979 5185 15991 5188
rect 15933 5179 15991 5185
rect 16022 5176 16028 5188
rect 16080 5176 16086 5228
rect 18693 5219 18751 5225
rect 18693 5185 18705 5219
rect 18739 5216 18751 5219
rect 19334 5216 19340 5228
rect 18739 5188 19340 5216
rect 18739 5185 18751 5188
rect 18693 5179 18751 5185
rect 19334 5176 19340 5188
rect 19392 5216 19398 5228
rect 19794 5216 19800 5228
rect 19392 5188 19800 5216
rect 19392 5176 19398 5188
rect 19794 5176 19800 5188
rect 19852 5176 19858 5228
rect 20070 5216 20076 5228
rect 20031 5188 20076 5216
rect 20070 5176 20076 5188
rect 20128 5176 20134 5228
rect 20162 5176 20168 5228
rect 20220 5216 20226 5228
rect 20220 5188 20265 5216
rect 20220 5176 20226 5188
rect 12805 5151 12863 5157
rect 12805 5148 12817 5151
rect 9324 5120 12817 5148
rect 5721 5083 5779 5089
rect 5721 5049 5733 5083
rect 5767 5080 5779 5083
rect 6914 5080 6920 5092
rect 5767 5052 6920 5080
rect 5767 5049 5779 5052
rect 5721 5043 5779 5049
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 7092 5083 7150 5089
rect 7092 5049 7104 5083
rect 7138 5080 7150 5083
rect 8202 5080 8208 5092
rect 7138 5052 8208 5080
rect 7138 5049 7150 5052
rect 7092 5043 7150 5049
rect 8202 5040 8208 5052
rect 8260 5040 8266 5092
rect 6086 4972 6092 5024
rect 6144 5012 6150 5024
rect 9324 5012 9352 5120
rect 12805 5117 12817 5120
rect 12851 5117 12863 5151
rect 12805 5111 12863 5117
rect 14185 5151 14243 5157
rect 14185 5117 14197 5151
rect 14231 5148 14243 5151
rect 14458 5148 14464 5160
rect 14231 5120 14464 5148
rect 14231 5117 14243 5120
rect 14185 5111 14243 5117
rect 14458 5108 14464 5120
rect 14516 5108 14522 5160
rect 14642 5108 14648 5160
rect 14700 5148 14706 5160
rect 14700 5120 15148 5148
rect 14700 5108 14706 5120
rect 9484 5083 9542 5089
rect 9484 5049 9496 5083
rect 9530 5080 9542 5083
rect 10686 5080 10692 5092
rect 9530 5052 10692 5080
rect 9530 5049 9542 5052
rect 9484 5043 9542 5049
rect 10686 5040 10692 5052
rect 10744 5040 10750 5092
rect 11054 5040 11060 5092
rect 11112 5080 11118 5092
rect 12897 5083 12955 5089
rect 12897 5080 12909 5083
rect 11112 5052 12909 5080
rect 11112 5040 11118 5052
rect 12897 5049 12909 5052
rect 12943 5049 12955 5083
rect 15120 5080 15148 5120
rect 15194 5108 15200 5160
rect 15252 5148 15258 5160
rect 15657 5151 15715 5157
rect 15657 5148 15669 5151
rect 15252 5120 15669 5148
rect 15252 5108 15258 5120
rect 15657 5117 15669 5120
rect 15703 5117 15715 5151
rect 15657 5111 15715 5117
rect 16853 5151 16911 5157
rect 16853 5117 16865 5151
rect 16899 5148 16911 5151
rect 17586 5148 17592 5160
rect 16899 5120 17592 5148
rect 16899 5117 16911 5120
rect 16853 5111 16911 5117
rect 17586 5108 17592 5120
rect 17644 5108 17650 5160
rect 18417 5151 18475 5157
rect 18417 5117 18429 5151
rect 18463 5148 18475 5151
rect 19242 5148 19248 5160
rect 18463 5120 19248 5148
rect 18463 5117 18475 5120
rect 18417 5111 18475 5117
rect 19242 5108 19248 5120
rect 19300 5108 19306 5160
rect 18509 5083 18567 5089
rect 18509 5080 18521 5083
rect 15120 5052 18521 5080
rect 12897 5043 12955 5049
rect 18509 5049 18521 5052
rect 18555 5080 18567 5083
rect 19150 5080 19156 5092
rect 18555 5052 19156 5080
rect 18555 5049 18567 5052
rect 18509 5043 18567 5049
rect 19150 5040 19156 5052
rect 19208 5040 19214 5092
rect 6144 4984 9352 5012
rect 6144 4972 6150 4984
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 14090 5012 14096 5024
rect 11756 4984 14096 5012
rect 11756 4972 11762 4984
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 14369 5015 14427 5021
rect 14369 4981 14381 5015
rect 14415 5012 14427 5015
rect 14734 5012 14740 5024
rect 14415 4984 14740 5012
rect 14415 4981 14427 4984
rect 14369 4975 14427 4981
rect 14734 4972 14740 4984
rect 14792 4972 14798 5024
rect 19426 4972 19432 5024
rect 19484 5012 19490 5024
rect 19613 5015 19671 5021
rect 19613 5012 19625 5015
rect 19484 4984 19625 5012
rect 19484 4972 19490 4984
rect 19613 4981 19625 4984
rect 19659 4981 19671 5015
rect 19978 5012 19984 5024
rect 19939 4984 19984 5012
rect 19613 4975 19671 4981
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 7650 4808 7656 4820
rect 7611 4780 7656 4808
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 8113 4811 8171 4817
rect 8113 4777 8125 4811
rect 8159 4808 8171 4811
rect 8386 4808 8392 4820
rect 8159 4780 8392 4808
rect 8159 4777 8171 4780
rect 8113 4771 8171 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 9677 4811 9735 4817
rect 9677 4777 9689 4811
rect 9723 4808 9735 4811
rect 10134 4808 10140 4820
rect 9723 4780 10140 4808
rect 9723 4777 9735 4780
rect 9677 4771 9735 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 11698 4808 11704 4820
rect 11659 4780 11704 4808
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 11793 4811 11851 4817
rect 11793 4777 11805 4811
rect 11839 4808 11851 4811
rect 11974 4808 11980 4820
rect 11839 4780 11980 4808
rect 11839 4777 11851 4780
rect 11793 4771 11851 4777
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 17954 4808 17960 4820
rect 13096 4780 17960 4808
rect 13096 4740 13124 4780
rect 17954 4768 17960 4780
rect 18012 4768 18018 4820
rect 15746 4740 15752 4752
rect 6564 4712 13124 4740
rect 15304 4712 15752 4740
rect 6564 4681 6592 4712
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4641 6607 4675
rect 6549 4635 6607 4641
rect 7650 4632 7656 4684
rect 7708 4672 7714 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7708 4644 8033 4672
rect 7708 4632 7714 4644
rect 8021 4641 8033 4644
rect 8067 4641 8079 4675
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 8021 4635 8079 4641
rect 8128 4644 10057 4672
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 8128 4604 8156 4644
rect 10045 4641 10057 4644
rect 10091 4641 10103 4675
rect 10045 4635 10103 4641
rect 12897 4675 12955 4681
rect 12897 4641 12909 4675
rect 12943 4672 12955 4675
rect 12986 4672 12992 4684
rect 12943 4644 12992 4672
rect 12943 4641 12955 4644
rect 12897 4635 12955 4641
rect 12986 4632 12992 4644
rect 13044 4632 13050 4684
rect 13164 4675 13222 4681
rect 13164 4641 13176 4675
rect 13210 4672 13222 4675
rect 13210 4644 15148 4672
rect 13210 4641 13222 4644
rect 13164 4635 13222 4641
rect 4856 4576 8156 4604
rect 4856 4564 4862 4576
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 8260 4576 8305 4604
rect 8260 4564 8266 4576
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 8444 4576 10149 4604
rect 8444 4564 8450 4576
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4604 10379 4607
rect 10686 4604 10692 4616
rect 10367 4576 10692 4604
rect 10367 4573 10379 4576
rect 10321 4567 10379 4573
rect 10152 4536 10180 4567
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 11974 4604 11980 4616
rect 11935 4576 11980 4604
rect 11974 4564 11980 4576
rect 12032 4564 12038 4616
rect 11698 4536 11704 4548
rect 10152 4508 11704 4536
rect 11698 4496 11704 4508
rect 11756 4496 11762 4548
rect 6730 4468 6736 4480
rect 6691 4440 6736 4468
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 8478 4428 8484 4480
rect 8536 4468 8542 4480
rect 11333 4471 11391 4477
rect 11333 4468 11345 4471
rect 8536 4440 11345 4468
rect 8536 4428 8542 4440
rect 11333 4437 11345 4440
rect 11379 4437 11391 4471
rect 14274 4468 14280 4480
rect 14235 4440 14280 4468
rect 11333 4431 11391 4437
rect 14274 4428 14280 4440
rect 14332 4428 14338 4480
rect 15120 4468 15148 4644
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 15304 4681 15332 4712
rect 15746 4700 15752 4712
rect 15804 4700 15810 4752
rect 15289 4675 15347 4681
rect 15289 4672 15301 4675
rect 15252 4644 15301 4672
rect 15252 4632 15258 4644
rect 15289 4641 15301 4644
rect 15335 4641 15347 4675
rect 15289 4635 15347 4641
rect 15556 4675 15614 4681
rect 15556 4641 15568 4675
rect 15602 4672 15614 4675
rect 17862 4672 17868 4684
rect 15602 4644 16528 4672
rect 17823 4644 17868 4672
rect 15602 4641 15614 4644
rect 15556 4635 15614 4641
rect 16500 4548 16528 4644
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 19058 4632 19064 4684
rect 19116 4672 19122 4684
rect 19613 4675 19671 4681
rect 19613 4672 19625 4675
rect 19116 4644 19625 4672
rect 19116 4632 19122 4644
rect 19613 4641 19625 4644
rect 19659 4641 19671 4675
rect 19613 4635 19671 4641
rect 17954 4604 17960 4616
rect 17915 4576 17960 4604
rect 17954 4564 17960 4576
rect 18012 4564 18018 4616
rect 18049 4607 18107 4613
rect 18049 4573 18061 4607
rect 18095 4573 18107 4607
rect 18049 4567 18107 4573
rect 16482 4496 16488 4548
rect 16540 4536 16546 4548
rect 18064 4536 18092 4567
rect 18966 4564 18972 4616
rect 19024 4604 19030 4616
rect 19705 4607 19763 4613
rect 19705 4604 19717 4607
rect 19024 4576 19717 4604
rect 19024 4564 19030 4576
rect 19705 4573 19717 4576
rect 19751 4573 19763 4607
rect 19705 4567 19763 4573
rect 19794 4564 19800 4616
rect 19852 4604 19858 4616
rect 19852 4576 19897 4604
rect 19852 4564 19858 4576
rect 16540 4508 18092 4536
rect 16540 4496 16546 4508
rect 16298 4468 16304 4480
rect 15120 4440 16304 4468
rect 16298 4428 16304 4440
rect 16356 4468 16362 4480
rect 16669 4471 16727 4477
rect 16669 4468 16681 4471
rect 16356 4440 16681 4468
rect 16356 4428 16362 4440
rect 16669 4437 16681 4440
rect 16715 4437 16727 4471
rect 17494 4468 17500 4480
rect 17455 4440 17500 4468
rect 16669 4431 16727 4437
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 19245 4471 19303 4477
rect 19245 4437 19257 4471
rect 19291 4468 19303 4471
rect 20070 4468 20076 4480
rect 19291 4440 20076 4468
rect 19291 4437 19303 4440
rect 19245 4431 19303 4437
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 8202 4264 8208 4276
rect 8163 4236 8208 4264
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 16482 4264 16488 4276
rect 9692 4236 16344 4264
rect 16443 4236 16488 4264
rect 9692 4196 9720 4236
rect 16316 4196 16344 4236
rect 16482 4224 16488 4236
rect 16540 4224 16546 4276
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 20162 4264 20168 4276
rect 19392 4236 20168 4264
rect 19392 4224 19398 4236
rect 20162 4224 20168 4236
rect 20220 4224 20226 4276
rect 18046 4196 18052 4208
rect 8220 4168 9720 4196
rect 14200 4168 15148 4196
rect 16316 4168 18052 4196
rect 8220 4140 8248 4168
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 6696 4100 6837 4128
rect 6696 4088 6702 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 8202 4088 8208 4140
rect 8260 4088 8266 4140
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 14200 4137 14228 4168
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 9272 4100 9873 4128
rect 9272 4088 9278 4100
rect 9861 4097 9873 4100
rect 9907 4097 9919 4131
rect 14185 4131 14243 4137
rect 9861 4091 9919 4097
rect 10888 4100 13952 4128
rect 9766 4060 9772 4072
rect 6932 4032 9772 4060
rect 2866 3952 2872 4004
rect 2924 3992 2930 4004
rect 6932 3992 6960 4032
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 10128 4063 10186 4069
rect 10128 4029 10140 4063
rect 10174 4060 10186 4063
rect 10502 4060 10508 4072
rect 10174 4032 10508 4060
rect 10174 4029 10186 4032
rect 10128 4023 10186 4029
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 10594 4020 10600 4072
rect 10652 4060 10658 4072
rect 10888 4060 10916 4100
rect 10652 4032 10916 4060
rect 12437 4063 12495 4069
rect 10652 4020 10658 4032
rect 12437 4029 12449 4063
rect 12483 4060 12495 4063
rect 12802 4060 12808 4072
rect 12483 4032 12808 4060
rect 12483 4029 12495 4032
rect 12437 4023 12495 4029
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 13924 4069 13952 4100
rect 14185 4097 14197 4131
rect 14231 4097 14243 4131
rect 15120 4128 15148 4168
rect 18046 4156 18052 4168
rect 18104 4156 18110 4208
rect 15120 4100 15240 4128
rect 14185 4091 14243 4097
rect 13909 4063 13967 4069
rect 13909 4029 13921 4063
rect 13955 4029 13967 4063
rect 13909 4023 13967 4029
rect 14001 4063 14059 4069
rect 14001 4029 14013 4063
rect 14047 4060 14059 4063
rect 14090 4060 14096 4072
rect 14047 4032 14096 4060
rect 14047 4029 14059 4032
rect 14001 4023 14059 4029
rect 14090 4020 14096 4032
rect 14148 4020 14154 4072
rect 15102 4060 15108 4072
rect 15063 4032 15108 4060
rect 15102 4020 15108 4032
rect 15160 4020 15166 4072
rect 2924 3964 6960 3992
rect 7092 3995 7150 4001
rect 2924 3952 2930 3964
rect 7092 3961 7104 3995
rect 7138 3992 7150 3995
rect 8570 3992 8576 4004
rect 7138 3964 8576 3992
rect 7138 3961 7150 3964
rect 7092 3955 7150 3961
rect 8570 3952 8576 3964
rect 8628 3952 8634 4004
rect 15212 3992 15240 4100
rect 16114 4088 16120 4140
rect 16172 4128 16178 4140
rect 17218 4128 17224 4140
rect 16172 4100 17224 4128
rect 16172 4088 16178 4100
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 15746 4020 15752 4072
rect 15804 4060 15810 4072
rect 16390 4060 16396 4072
rect 15804 4032 16396 4060
rect 15804 4020 15810 4032
rect 16390 4020 16396 4032
rect 16448 4060 16454 4072
rect 19061 4063 19119 4069
rect 19061 4060 19073 4063
rect 16448 4032 19073 4060
rect 16448 4020 16454 4032
rect 19061 4029 19073 4032
rect 19107 4029 19119 4063
rect 19061 4023 19119 4029
rect 19168 4032 19656 4060
rect 15378 4001 15384 4004
rect 15372 3992 15384 4001
rect 8680 3964 14504 3992
rect 15212 3964 15384 3992
rect 5718 3924 5724 3936
rect 5679 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 7190 3884 7196 3936
rect 7248 3924 7254 3936
rect 8680 3924 8708 3964
rect 7248 3896 8708 3924
rect 7248 3884 7254 3896
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 10226 3924 10232 3936
rect 8812 3896 10232 3924
rect 8812 3884 8818 3896
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 11238 3924 11244 3936
rect 11199 3896 11244 3924
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12621 3927 12679 3933
rect 12621 3924 12633 3927
rect 12492 3896 12633 3924
rect 12492 3884 12498 3896
rect 12621 3893 12633 3896
rect 12667 3893 12679 3927
rect 13538 3924 13544 3936
rect 13499 3896 13544 3924
rect 12621 3887 12679 3893
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 14476 3924 14504 3964
rect 15372 3955 15384 3964
rect 15378 3952 15384 3955
rect 15436 3952 15442 4004
rect 15470 3952 15476 4004
rect 15528 3992 15534 4004
rect 16758 3992 16764 4004
rect 15528 3964 16764 3992
rect 15528 3952 15534 3964
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 17126 3952 17132 4004
rect 17184 3992 17190 4004
rect 19168 3992 19196 4032
rect 19334 4001 19340 4004
rect 17184 3964 19196 3992
rect 17184 3952 17190 3964
rect 19328 3955 19340 4001
rect 19392 3992 19398 4004
rect 19628 3992 19656 4032
rect 19392 3964 19428 3992
rect 19628 3964 20484 3992
rect 19334 3952 19340 3955
rect 19392 3952 19398 3964
rect 17586 3924 17592 3936
rect 14476 3896 17592 3924
rect 17586 3884 17592 3896
rect 17644 3884 17650 3936
rect 18049 3927 18107 3933
rect 18049 3893 18061 3927
rect 18095 3924 18107 3927
rect 19978 3924 19984 3936
rect 18095 3896 19984 3924
rect 18095 3893 18107 3896
rect 18049 3887 18107 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 20456 3933 20484 3964
rect 20441 3927 20499 3933
rect 20441 3893 20453 3927
rect 20487 3893 20499 3927
rect 20441 3887 20499 3893
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 6454 3720 6460 3732
rect 5684 3692 6460 3720
rect 5684 3680 5690 3692
rect 6454 3680 6460 3692
rect 6512 3680 6518 3732
rect 7101 3723 7159 3729
rect 7101 3689 7113 3723
rect 7147 3720 7159 3723
rect 7190 3720 7196 3732
rect 7147 3692 7196 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 7558 3680 7564 3732
rect 7616 3720 7622 3732
rect 8021 3723 8079 3729
rect 8021 3720 8033 3723
rect 7616 3692 8033 3720
rect 7616 3680 7622 3692
rect 8021 3689 8033 3692
rect 8067 3689 8079 3723
rect 8478 3720 8484 3732
rect 8439 3692 8484 3720
rect 8021 3683 8079 3689
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 9674 3720 9680 3732
rect 8588 3692 9680 3720
rect 5994 3612 6000 3664
rect 6052 3652 6058 3664
rect 8588 3652 8616 3692
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 13354 3680 13360 3732
rect 13412 3720 13418 3732
rect 15470 3720 15476 3732
rect 13412 3692 15476 3720
rect 13412 3680 13418 3692
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 15657 3723 15715 3729
rect 15657 3689 15669 3723
rect 15703 3720 15715 3723
rect 15746 3720 15752 3732
rect 15703 3692 15752 3720
rect 15703 3689 15715 3692
rect 15657 3683 15715 3689
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 16117 3723 16175 3729
rect 16117 3689 16129 3723
rect 16163 3720 16175 3723
rect 17494 3720 17500 3732
rect 16163 3692 17500 3720
rect 16163 3689 16175 3692
rect 16117 3683 16175 3689
rect 17494 3680 17500 3692
rect 17552 3680 17558 3732
rect 17586 3680 17592 3732
rect 17644 3720 17650 3732
rect 19978 3720 19984 3732
rect 17644 3692 19984 3720
rect 17644 3680 17650 3692
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 6052 3624 8616 3652
rect 6052 3612 6058 3624
rect 9214 3612 9220 3664
rect 9272 3652 9278 3664
rect 10594 3652 10600 3664
rect 9272 3624 10600 3652
rect 9272 3612 9278 3624
rect 10594 3612 10600 3624
rect 10652 3612 10658 3664
rect 10864 3655 10922 3661
rect 10864 3621 10876 3655
rect 10910 3652 10922 3655
rect 11238 3652 11244 3664
rect 10910 3624 11244 3652
rect 10910 3621 10922 3624
rect 10864 3615 10922 3621
rect 11238 3612 11244 3624
rect 11296 3612 11302 3664
rect 16758 3652 16764 3664
rect 12636 3624 16764 3652
rect 5810 3584 5816 3596
rect 5771 3556 5816 3584
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 8202 3584 8208 3596
rect 6963 3556 8208 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 8386 3584 8392 3596
rect 8347 3556 8392 3584
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 8570 3544 8576 3596
rect 8628 3544 8634 3596
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 8904 3556 11652 3584
rect 8904 3544 8910 3556
rect 8588 3516 8616 3544
rect 8665 3519 8723 3525
rect 8665 3516 8677 3519
rect 8588 3488 8677 3516
rect 8665 3485 8677 3488
rect 8711 3516 8723 3519
rect 9306 3516 9312 3528
rect 8711 3488 9312 3516
rect 8711 3485 8723 3488
rect 8665 3479 8723 3485
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 10594 3516 10600 3528
rect 10555 3488 10600 3516
rect 10594 3476 10600 3488
rect 10652 3476 10658 3528
rect 11624 3516 11652 3556
rect 11624 3488 12388 3516
rect 3326 3408 3332 3460
rect 3384 3448 3390 3460
rect 4798 3448 4804 3460
rect 3384 3420 4804 3448
rect 3384 3408 3390 3420
rect 4798 3408 4804 3420
rect 4856 3408 4862 3460
rect 4982 3448 4988 3460
rect 4943 3420 4988 3448
rect 4982 3408 4988 3420
rect 5040 3408 5046 3460
rect 5997 3451 6055 3457
rect 5997 3417 6009 3451
rect 6043 3448 6055 3451
rect 12250 3448 12256 3460
rect 6043 3420 10640 3448
rect 6043 3417 6055 3420
rect 5997 3411 6055 3417
rect 5534 3340 5540 3392
rect 5592 3380 5598 3392
rect 8754 3380 8760 3392
rect 5592 3352 8760 3380
rect 5592 3340 5598 3352
rect 8754 3340 8760 3352
rect 8812 3340 8818 3392
rect 10612 3380 10640 3420
rect 11900 3420 12256 3448
rect 11900 3380 11928 3420
rect 12250 3408 12256 3420
rect 12308 3408 12314 3460
rect 10612 3352 11928 3380
rect 11974 3340 11980 3392
rect 12032 3380 12038 3392
rect 12360 3380 12388 3488
rect 12636 3380 12664 3624
rect 16758 3612 16764 3624
rect 16816 3612 16822 3664
rect 16942 3612 16948 3664
rect 17000 3652 17006 3664
rect 19705 3655 19763 3661
rect 19705 3652 19717 3655
rect 17000 3624 19717 3652
rect 17000 3612 17006 3624
rect 19705 3621 19717 3624
rect 19751 3621 19763 3655
rect 19705 3615 19763 3621
rect 13072 3587 13130 3593
rect 13072 3553 13084 3587
rect 13118 3584 13130 3587
rect 14274 3584 14280 3596
rect 13118 3556 14280 3584
rect 13118 3553 13130 3556
rect 13072 3547 13130 3553
rect 14274 3544 14280 3556
rect 14332 3544 14338 3596
rect 15654 3544 15660 3596
rect 15712 3584 15718 3596
rect 16025 3587 16083 3593
rect 16025 3584 16037 3587
rect 15712 3556 16037 3584
rect 15712 3544 15718 3556
rect 16025 3553 16037 3556
rect 16071 3553 16083 3587
rect 16025 3547 16083 3553
rect 17126 3544 17132 3596
rect 17184 3584 17190 3596
rect 17477 3587 17535 3593
rect 17477 3584 17489 3587
rect 17184 3556 17489 3584
rect 17184 3544 17190 3556
rect 17477 3553 17489 3556
rect 17523 3553 17535 3587
rect 19426 3584 19432 3596
rect 19387 3556 19432 3584
rect 17477 3547 17535 3553
rect 19426 3544 19432 3556
rect 19484 3544 19490 3596
rect 20346 3544 20352 3596
rect 20404 3584 20410 3596
rect 21542 3584 21548 3596
rect 20404 3556 21548 3584
rect 20404 3544 20410 3556
rect 21542 3544 21548 3556
rect 21600 3544 21606 3596
rect 12802 3516 12808 3528
rect 12763 3488 12808 3516
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 16298 3516 16304 3528
rect 16259 3488 16304 3516
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 16390 3476 16396 3528
rect 16448 3516 16454 3528
rect 17221 3519 17279 3525
rect 17221 3516 17233 3519
rect 16448 3488 17233 3516
rect 16448 3476 16454 3488
rect 17221 3485 17233 3488
rect 17267 3485 17279 3519
rect 17221 3479 17279 3485
rect 14090 3408 14096 3460
rect 14148 3448 14154 3460
rect 19702 3448 19708 3460
rect 14148 3420 15792 3448
rect 14148 3408 14154 3420
rect 12032 3352 12077 3380
rect 12360 3352 12664 3380
rect 12032 3340 12038 3352
rect 12986 3340 12992 3392
rect 13044 3380 13050 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 13044 3352 14197 3380
rect 13044 3340 13050 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 15764 3380 15792 3420
rect 18156 3420 19708 3448
rect 18156 3380 18184 3420
rect 19702 3408 19708 3420
rect 19760 3408 19766 3460
rect 18598 3380 18604 3392
rect 15764 3352 18184 3380
rect 18559 3352 18604 3380
rect 14185 3343 14243 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 7006 3176 7012 3188
rect 6967 3148 7012 3176
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 9306 3176 9312 3188
rect 7116 3148 8892 3176
rect 9267 3148 9312 3176
rect 3878 3068 3884 3120
rect 3936 3108 3942 3120
rect 7116 3108 7144 3148
rect 3936 3080 7144 3108
rect 8864 3108 8892 3148
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 10781 3179 10839 3185
rect 10781 3145 10793 3179
rect 10827 3176 10839 3179
rect 10962 3176 10968 3188
rect 10827 3148 10968 3176
rect 10827 3145 10839 3148
rect 10781 3139 10839 3145
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 12526 3136 12532 3188
rect 12584 3176 12590 3188
rect 15194 3176 15200 3188
rect 12584 3148 15200 3176
rect 12584 3136 12590 3148
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 15654 3176 15660 3188
rect 15615 3148 15660 3176
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 15746 3136 15752 3188
rect 15804 3176 15810 3188
rect 15804 3148 16252 3176
rect 15804 3136 15810 3148
rect 8864 3080 8984 3108
rect 3936 3068 3942 3080
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 7929 3043 7987 3049
rect 7929 3040 7941 3043
rect 6788 3012 7941 3040
rect 6788 3000 6794 3012
rect 7929 3009 7941 3012
rect 7975 3009 7987 3043
rect 8956 3040 8984 3080
rect 10502 3068 10508 3120
rect 10560 3108 10566 3120
rect 10560 3080 11468 3108
rect 10560 3068 10566 3080
rect 11054 3040 11060 3052
rect 8956 3012 11060 3040
rect 7929 3003 7987 3009
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 11333 3043 11391 3049
rect 11333 3040 11345 3043
rect 11296 3012 11345 3040
rect 11296 3000 11302 3012
rect 11333 3009 11345 3012
rect 11379 3009 11391 3043
rect 11440 3040 11468 3080
rect 11882 3068 11888 3120
rect 11940 3108 11946 3120
rect 11940 3080 13216 3108
rect 11940 3068 11946 3080
rect 12986 3040 12992 3052
rect 11440 3012 12992 3040
rect 11333 3003 11391 3009
rect 12986 3000 12992 3012
rect 13044 3040 13050 3052
rect 13081 3043 13139 3049
rect 13081 3040 13093 3043
rect 13044 3012 13093 3040
rect 13044 3000 13050 3012
rect 13081 3009 13093 3012
rect 13127 3009 13139 3043
rect 13188 3040 13216 3080
rect 13538 3068 13544 3120
rect 13596 3108 13602 3120
rect 16224 3108 16252 3148
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 18012 3148 18061 3176
rect 18012 3136 18018 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 19610 3176 19616 3188
rect 19571 3148 19616 3176
rect 18049 3139 18107 3145
rect 19610 3136 19616 3148
rect 19668 3136 19674 3188
rect 13596 3080 16160 3108
rect 16224 3080 18920 3108
rect 13596 3068 13602 3080
rect 13630 3040 13636 3052
rect 13188 3012 13636 3040
rect 13081 3003 13139 3009
rect 13630 3000 13636 3012
rect 13688 3000 13694 3052
rect 13722 3000 13728 3052
rect 13780 3040 13786 3052
rect 14274 3040 14280 3052
rect 13780 3012 14280 3040
rect 13780 3000 13786 3012
rect 14274 3000 14280 3012
rect 14332 3040 14338 3052
rect 16132 3049 16160 3080
rect 14645 3043 14703 3049
rect 14645 3040 14657 3043
rect 14332 3012 14657 3040
rect 14332 3000 14338 3012
rect 14645 3009 14657 3012
rect 14691 3009 14703 3043
rect 16117 3043 16175 3049
rect 14645 3003 14703 3009
rect 15856 3012 16059 3040
rect 5629 2975 5687 2981
rect 5629 2941 5641 2975
rect 5675 2972 5687 2975
rect 6850 2975 6908 2981
rect 5675 2944 6776 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 4617 2907 4675 2913
rect 4617 2873 4629 2907
rect 4663 2904 4675 2907
rect 6748 2904 6776 2944
rect 6850 2941 6862 2975
rect 6896 2972 6908 2975
rect 7374 2972 7380 2984
rect 6896 2944 7380 2972
rect 6896 2941 6908 2944
rect 6850 2935 6908 2941
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 15856 2972 15884 3012
rect 7668 2944 15884 2972
rect 7668 2904 7696 2944
rect 15930 2932 15936 2984
rect 15988 2932 15994 2984
rect 16031 2972 16059 3012
rect 16117 3009 16129 3043
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3040 16359 3043
rect 16482 3040 16488 3052
rect 16347 3012 16488 3040
rect 16347 3009 16359 3012
rect 16301 3003 16359 3009
rect 16482 3000 16488 3012
rect 16540 3000 16546 3052
rect 17402 3000 17408 3052
rect 17460 3040 17466 3052
rect 18598 3040 18604 3052
rect 17460 3012 18604 3040
rect 17460 3000 17466 3012
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 18046 2972 18052 2984
rect 16031 2944 18052 2972
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18417 2975 18475 2981
rect 18417 2941 18429 2975
rect 18463 2972 18475 2975
rect 18782 2972 18788 2984
rect 18463 2944 18788 2972
rect 18463 2941 18475 2944
rect 18417 2935 18475 2941
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 18892 2972 18920 3080
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 19702 3108 19708 3120
rect 19484 3080 19708 3108
rect 19484 3068 19490 3080
rect 19702 3068 19708 3080
rect 19760 3068 19766 3120
rect 20070 3040 20076 3052
rect 20031 3012 20076 3040
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 20162 3000 20168 3052
rect 20220 3040 20226 3052
rect 20220 3012 20265 3040
rect 20220 3000 20226 3012
rect 20254 2972 20260 2984
rect 18892 2944 20260 2972
rect 20254 2932 20260 2944
rect 20312 2932 20318 2984
rect 4663 2876 6592 2904
rect 6748 2876 7696 2904
rect 8196 2907 8254 2913
rect 4663 2873 4675 2876
rect 4617 2867 4675 2873
rect 198 2796 204 2848
rect 256 2836 262 2848
rect 5534 2836 5540 2848
rect 256 2808 5540 2836
rect 256 2796 262 2808
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 5810 2836 5816 2848
rect 5771 2808 5816 2836
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 6564 2836 6592 2876
rect 8196 2873 8208 2907
rect 8242 2904 8254 2907
rect 8662 2904 8668 2916
rect 8242 2876 8668 2904
rect 8242 2873 8254 2876
rect 8196 2867 8254 2873
rect 8662 2864 8668 2876
rect 8720 2904 8726 2916
rect 11974 2904 11980 2916
rect 8720 2876 11980 2904
rect 8720 2864 8726 2876
rect 11974 2864 11980 2876
rect 12032 2864 12038 2916
rect 12897 2907 12955 2913
rect 12897 2873 12909 2907
rect 12943 2904 12955 2907
rect 14553 2907 14611 2913
rect 12943 2876 13952 2904
rect 12943 2873 12955 2876
rect 12897 2867 12955 2873
rect 10226 2836 10232 2848
rect 6564 2808 10232 2836
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 11146 2836 11152 2848
rect 11107 2808 11152 2836
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 11241 2839 11299 2845
rect 11241 2805 11253 2839
rect 11287 2836 11299 2839
rect 12529 2839 12587 2845
rect 12529 2836 12541 2839
rect 11287 2808 12541 2836
rect 11287 2805 11299 2808
rect 11241 2799 11299 2805
rect 12529 2805 12541 2808
rect 12575 2805 12587 2839
rect 12529 2799 12587 2805
rect 12986 2796 12992 2848
rect 13044 2836 13050 2848
rect 13924 2836 13952 2876
rect 14553 2873 14565 2907
rect 14599 2904 14611 2907
rect 14642 2904 14648 2916
rect 14599 2876 14648 2904
rect 14599 2873 14611 2876
rect 14553 2867 14611 2873
rect 14642 2864 14648 2876
rect 14700 2864 14706 2916
rect 15948 2904 15976 2932
rect 16025 2907 16083 2913
rect 16025 2904 16037 2907
rect 15948 2876 16037 2904
rect 16025 2873 16037 2876
rect 16071 2873 16083 2907
rect 16025 2867 16083 2873
rect 18138 2864 18144 2916
rect 18196 2904 18202 2916
rect 18509 2907 18567 2913
rect 18509 2904 18521 2907
rect 18196 2876 18521 2904
rect 18196 2864 18202 2876
rect 18509 2873 18521 2876
rect 18555 2873 18567 2907
rect 18509 2867 18567 2873
rect 19886 2864 19892 2916
rect 19944 2904 19950 2916
rect 19981 2907 20039 2913
rect 19981 2904 19993 2907
rect 19944 2876 19993 2904
rect 19944 2864 19950 2876
rect 19981 2873 19993 2876
rect 20027 2873 20039 2907
rect 19981 2867 20039 2873
rect 14093 2839 14151 2845
rect 14093 2836 14105 2839
rect 13044 2808 13089 2836
rect 13924 2808 14105 2836
rect 13044 2796 13050 2808
rect 14093 2805 14105 2808
rect 14139 2805 14151 2839
rect 14458 2836 14464 2848
rect 14419 2808 14464 2836
rect 14093 2799 14151 2805
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 16206 2836 16212 2848
rect 15252 2808 16212 2836
rect 15252 2796 15258 2808
rect 16206 2796 16212 2808
rect 16264 2796 16270 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 8113 2635 8171 2641
rect 8113 2601 8125 2635
rect 8159 2632 8171 2635
rect 8386 2632 8392 2644
rect 8159 2604 8392 2632
rect 8159 2601 8171 2604
rect 8113 2595 8171 2601
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 10226 2632 10232 2644
rect 10187 2604 10232 2632
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 12986 2592 12992 2644
rect 13044 2632 13050 2644
rect 13081 2635 13139 2641
rect 13081 2632 13093 2635
rect 13044 2604 13093 2632
rect 13044 2592 13050 2604
rect 13081 2601 13093 2604
rect 13127 2601 13139 2635
rect 13081 2595 13139 2601
rect 16669 2635 16727 2641
rect 16669 2601 16681 2635
rect 16715 2632 16727 2635
rect 17862 2632 17868 2644
rect 16715 2604 17868 2632
rect 16715 2601 16727 2604
rect 16669 2595 16727 2601
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 8202 2524 8208 2576
rect 8260 2564 8266 2576
rect 8573 2567 8631 2573
rect 8573 2564 8585 2567
rect 8260 2536 8585 2564
rect 8260 2524 8266 2536
rect 8573 2533 8585 2536
rect 8619 2533 8631 2567
rect 8573 2527 8631 2533
rect 11698 2524 11704 2576
rect 11756 2564 11762 2576
rect 11756 2536 13584 2564
rect 11756 2524 11762 2536
rect 7006 2496 7012 2508
rect 6967 2468 7012 2496
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2465 8539 2499
rect 8481 2459 8539 2465
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 8496 2428 8524 2459
rect 11238 2456 11244 2508
rect 11296 2496 11302 2508
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 11296 2468 11437 2496
rect 11296 2456 11302 2468
rect 11425 2465 11437 2468
rect 11471 2465 11483 2499
rect 13446 2496 13452 2508
rect 13407 2468 13452 2496
rect 11425 2459 11483 2465
rect 13446 2456 13452 2468
rect 13504 2456 13510 2508
rect 13556 2505 13584 2536
rect 15378 2524 15384 2576
rect 15436 2564 15442 2576
rect 17402 2564 17408 2576
rect 15436 2536 17408 2564
rect 15436 2524 15442 2536
rect 17402 2524 17408 2536
rect 17460 2524 17466 2576
rect 13541 2499 13599 2505
rect 13541 2465 13553 2499
rect 13587 2496 13599 2499
rect 15473 2499 15531 2505
rect 13587 2468 15424 2496
rect 13587 2465 13599 2468
rect 13541 2459 13599 2465
rect 8662 2428 8668 2440
rect 5859 2400 8524 2428
rect 8623 2400 8668 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 8812 2400 10333 2428
rect 8812 2388 8818 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10502 2428 10508 2440
rect 10463 2400 10508 2428
rect 10321 2391 10379 2397
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 13722 2428 13728 2440
rect 13683 2400 13728 2428
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 15396 2428 15424 2468
rect 15473 2465 15485 2499
rect 15519 2496 15531 2499
rect 16666 2496 16672 2508
rect 15519 2468 16672 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 17034 2496 17040 2508
rect 16995 2468 17040 2496
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 16577 2431 16635 2437
rect 16577 2428 16589 2431
rect 15396 2400 16589 2428
rect 16577 2397 16589 2400
rect 16623 2397 16635 2431
rect 17126 2428 17132 2440
rect 17087 2400 17132 2428
rect 16577 2391 16635 2397
rect 17126 2388 17132 2400
rect 17184 2388 17190 2440
rect 17313 2431 17371 2437
rect 17313 2397 17325 2431
rect 17359 2428 17371 2431
rect 17420 2428 17448 2524
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 18966 2496 18972 2508
rect 18012 2468 18972 2496
rect 18012 2456 18018 2468
rect 18966 2456 18972 2468
rect 19024 2496 19030 2508
rect 19242 2496 19248 2508
rect 19024 2468 19248 2496
rect 19024 2456 19030 2468
rect 19242 2456 19248 2468
rect 19300 2456 19306 2508
rect 19429 2499 19487 2505
rect 19429 2496 19441 2499
rect 19352 2468 19441 2496
rect 17359 2400 17448 2428
rect 17359 2397 17371 2400
rect 17313 2391 17371 2397
rect 5718 2320 5724 2372
rect 5776 2360 5782 2372
rect 9861 2363 9919 2369
rect 5776 2332 7328 2360
rect 5776 2320 5782 2332
rect 7190 2292 7196 2304
rect 7151 2264 7196 2292
rect 7190 2252 7196 2264
rect 7248 2252 7254 2304
rect 7300 2292 7328 2332
rect 9861 2329 9873 2363
rect 9907 2360 9919 2363
rect 11146 2360 11152 2372
rect 9907 2332 11152 2360
rect 9907 2329 9919 2332
rect 9861 2323 9919 2329
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 19352 2360 19380 2468
rect 19429 2465 19441 2468
rect 19475 2465 19487 2499
rect 19429 2459 19487 2465
rect 19518 2428 19524 2440
rect 19479 2400 19524 2428
rect 19518 2388 19524 2400
rect 19576 2388 19582 2440
rect 19705 2431 19763 2437
rect 19705 2397 19717 2431
rect 19751 2428 19763 2431
rect 20162 2428 20168 2440
rect 19751 2400 20168 2428
rect 19751 2397 19763 2400
rect 19705 2391 19763 2397
rect 20162 2388 20168 2400
rect 20220 2388 20226 2440
rect 11256 2332 19380 2360
rect 11256 2292 11284 2332
rect 7300 2264 11284 2292
rect 11609 2295 11667 2301
rect 11609 2261 11621 2295
rect 11655 2292 11667 2295
rect 11698 2292 11704 2304
rect 11655 2264 11704 2292
rect 11655 2261 11667 2264
rect 11609 2255 11667 2261
rect 11698 2252 11704 2264
rect 11756 2252 11762 2304
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 13596 2264 15669 2292
rect 13596 2252 13602 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 16577 2295 16635 2301
rect 16577 2261 16589 2295
rect 16623 2292 16635 2295
rect 17954 2292 17960 2304
rect 16623 2264 17960 2292
rect 16623 2261 16635 2264
rect 16577 2255 16635 2261
rect 17954 2252 17960 2264
rect 18012 2252 18018 2304
rect 19058 2292 19064 2304
rect 19019 2264 19064 2292
rect 19058 2252 19064 2264
rect 19116 2252 19122 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 7190 2048 7196 2100
rect 7248 2088 7254 2100
rect 20438 2088 20444 2100
rect 7248 2060 20444 2088
rect 7248 2048 7254 2060
rect 20438 2048 20444 2060
rect 20496 2048 20502 2100
rect 9766 1980 9772 2032
rect 9824 2020 9830 2032
rect 19518 2020 19524 2032
rect 9824 1992 19524 2020
rect 9824 1980 9830 1992
rect 19518 1980 19524 1992
rect 19576 1980 19582 2032
rect 7006 1912 7012 1964
rect 7064 1952 7070 1964
rect 7064 1924 13400 1952
rect 7064 1912 7070 1924
rect 13372 1748 13400 1924
rect 13998 1912 14004 1964
rect 14056 1952 14062 1964
rect 19058 1952 19064 1964
rect 14056 1924 19064 1952
rect 14056 1912 14062 1924
rect 19058 1912 19064 1924
rect 19116 1912 19122 1964
rect 17126 1844 17132 1896
rect 17184 1884 17190 1896
rect 17310 1884 17316 1896
rect 17184 1856 17316 1884
rect 17184 1844 17190 1856
rect 17310 1844 17316 1856
rect 17368 1844 17374 1896
rect 13446 1776 13452 1828
rect 13504 1816 13510 1828
rect 18966 1816 18972 1828
rect 13504 1788 18972 1816
rect 13504 1776 13510 1788
rect 18966 1776 18972 1788
rect 19024 1776 19030 1828
rect 18690 1748 18696 1760
rect 13372 1720 18696 1748
rect 18690 1708 18696 1720
rect 18748 1708 18754 1760
rect 9858 1640 9864 1692
rect 9916 1680 9922 1692
rect 18322 1680 18328 1692
rect 9916 1652 18328 1680
rect 9916 1640 9922 1652
rect 18322 1640 18328 1652
rect 18380 1640 18386 1692
rect 12158 1096 12164 1148
rect 12216 1136 12222 1148
rect 17770 1136 17776 1148
rect 12216 1108 17776 1136
rect 12216 1096 12222 1108
rect 17770 1096 17776 1108
rect 17828 1096 17834 1148
rect 19426 552 19432 604
rect 19484 592 19490 604
rect 19702 592 19708 604
rect 19484 564 19708 592
rect 19484 552 19490 564
rect 19702 552 19708 564
rect 19760 552 19766 604
<< via1 >>
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 19064 20587 19116 20596
rect 19064 20553 19073 20587
rect 19073 20553 19107 20587
rect 19107 20553 19116 20587
rect 19064 20544 19116 20553
rect 19800 20340 19852 20392
rect 17960 20272 18012 20324
rect 20168 20247 20220 20256
rect 20168 20213 20177 20247
rect 20177 20213 20211 20247
rect 20211 20213 20220 20247
rect 20168 20204 20220 20213
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 2872 20000 2924 20052
rect 18788 20043 18840 20052
rect 18788 20009 18797 20043
rect 18797 20009 18831 20043
rect 18831 20009 18840 20043
rect 18788 20000 18840 20009
rect 15844 19932 15896 19984
rect 18604 19907 18656 19916
rect 18604 19873 18613 19907
rect 18613 19873 18647 19907
rect 18647 19873 18656 19907
rect 18604 19864 18656 19873
rect 20076 19796 20128 19848
rect 19892 19771 19944 19780
rect 19892 19737 19901 19771
rect 19901 19737 19935 19771
rect 19935 19737 19944 19771
rect 19892 19728 19944 19737
rect 4804 19660 4856 19712
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 4804 19456 4856 19508
rect 20720 19456 20772 19508
rect 10784 19252 10836 19304
rect 14004 19295 14056 19304
rect 14004 19261 14013 19295
rect 14013 19261 14047 19295
rect 14047 19261 14056 19295
rect 14004 19252 14056 19261
rect 17960 19252 18012 19304
rect 14372 19184 14424 19236
rect 19156 19252 19208 19304
rect 14188 19116 14240 19168
rect 18972 19159 19024 19168
rect 18972 19125 18981 19159
rect 18981 19125 19015 19159
rect 19015 19125 19024 19159
rect 18972 19116 19024 19125
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 14004 18912 14056 18964
rect 15200 18912 15252 18964
rect 18604 18844 18656 18896
rect 19800 18887 19852 18896
rect 19800 18853 19809 18887
rect 19809 18853 19843 18887
rect 19843 18853 19852 18887
rect 19800 18844 19852 18853
rect 9772 18776 9824 18828
rect 13912 18776 13964 18828
rect 16580 18776 16632 18828
rect 15844 18708 15896 18760
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 17960 18368 18012 18420
rect 19616 18411 19668 18420
rect 19616 18377 19625 18411
rect 19625 18377 19659 18411
rect 19659 18377 19668 18411
rect 19616 18368 19668 18377
rect 20720 18411 20772 18420
rect 20720 18377 20729 18411
rect 20729 18377 20763 18411
rect 20763 18377 20772 18411
rect 20720 18368 20772 18377
rect 9956 18164 10008 18216
rect 13268 18207 13320 18216
rect 13268 18173 13277 18207
rect 13277 18173 13311 18207
rect 13311 18173 13320 18207
rect 13268 18164 13320 18173
rect 20536 18207 20588 18216
rect 20536 18173 20545 18207
rect 20545 18173 20579 18207
rect 20579 18173 20588 18207
rect 20536 18164 20588 18173
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 12992 17688 13044 17740
rect 19892 17527 19944 17536
rect 19892 17493 19901 17527
rect 19901 17493 19935 17527
rect 19935 17493 19944 17527
rect 19892 17484 19944 17493
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 18972 17323 19024 17332
rect 18972 17289 18981 17323
rect 18981 17289 19015 17323
rect 19015 17289 19024 17323
rect 18972 17280 19024 17289
rect 13268 17144 13320 17196
rect 20536 17144 20588 17196
rect 12624 17076 12676 17128
rect 18788 17119 18840 17128
rect 18788 17085 18797 17119
rect 18797 17085 18831 17119
rect 18831 17085 18840 17119
rect 18788 17076 18840 17085
rect 10232 17008 10284 17060
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 18604 16779 18656 16788
rect 18604 16745 18613 16779
rect 18613 16745 18647 16779
rect 18647 16745 18656 16779
rect 18604 16736 18656 16745
rect 12992 16711 13044 16720
rect 12992 16677 13001 16711
rect 13001 16677 13035 16711
rect 13035 16677 13044 16711
rect 12992 16668 13044 16677
rect 16672 16668 16724 16720
rect 12716 16643 12768 16652
rect 12716 16609 12725 16643
rect 12725 16609 12759 16643
rect 12759 16609 12768 16643
rect 12716 16600 12768 16609
rect 14740 16600 14792 16652
rect 18788 16668 18840 16720
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 18604 16192 18656 16244
rect 17960 15988 18012 16040
rect 20536 16031 20588 16040
rect 18144 15920 18196 15972
rect 20536 15997 20545 16031
rect 20545 15997 20579 16031
rect 20579 15997 20588 16031
rect 20536 15988 20588 15997
rect 19248 15852 19300 15904
rect 20628 15852 20680 15904
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 18788 15691 18840 15700
rect 18788 15657 18797 15691
rect 18797 15657 18831 15691
rect 18831 15657 18840 15691
rect 18788 15648 18840 15657
rect 14740 15580 14792 15632
rect 10508 15555 10560 15564
rect 10508 15521 10517 15555
rect 10517 15521 10551 15555
rect 10551 15521 10560 15555
rect 10508 15512 10560 15521
rect 18604 15555 18656 15564
rect 18604 15521 18613 15555
rect 18613 15521 18647 15555
rect 18647 15521 18656 15555
rect 18604 15512 18656 15521
rect 19984 15512 20036 15564
rect 19892 15351 19944 15360
rect 19892 15317 19901 15351
rect 19901 15317 19935 15351
rect 19935 15317 19944 15351
rect 19892 15308 19944 15317
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 19064 15147 19116 15156
rect 19064 15113 19073 15147
rect 19073 15113 19107 15147
rect 19107 15113 19116 15147
rect 19064 15104 19116 15113
rect 13636 14968 13688 15020
rect 7104 14900 7156 14952
rect 9036 14943 9088 14952
rect 9036 14909 9045 14943
rect 9045 14909 9079 14943
rect 9079 14909 9088 14943
rect 9036 14900 9088 14909
rect 17960 14900 18012 14952
rect 18880 14943 18932 14952
rect 18880 14909 18889 14943
rect 18889 14909 18923 14943
rect 18923 14909 18932 14943
rect 18880 14900 18932 14909
rect 18604 14832 18656 14884
rect 18696 14832 18748 14884
rect 19064 14764 19116 14816
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 18144 14492 18196 14544
rect 18880 14492 18932 14544
rect 7196 14424 7248 14476
rect 17316 14467 17368 14476
rect 17316 14433 17325 14467
rect 17325 14433 17359 14467
rect 17359 14433 17368 14467
rect 17316 14424 17368 14433
rect 18696 14424 18748 14476
rect 12532 14399 12584 14408
rect 12532 14365 12541 14399
rect 12541 14365 12575 14399
rect 12575 14365 12584 14399
rect 12532 14356 12584 14365
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 17868 14356 17920 14408
rect 7656 14288 7708 14340
rect 17776 14220 17828 14272
rect 18604 14263 18656 14272
rect 18604 14229 18613 14263
rect 18613 14229 18647 14263
rect 18647 14229 18656 14263
rect 18604 14220 18656 14229
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 12716 14016 12768 14068
rect 16580 14016 16632 14068
rect 10968 13948 11020 14000
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 16488 13880 16540 13932
rect 17316 13880 17368 13932
rect 12532 13812 12584 13864
rect 14648 13812 14700 13864
rect 18512 13855 18564 13864
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 19984 13923 20036 13932
rect 19984 13889 19993 13923
rect 19993 13889 20027 13923
rect 20027 13889 20036 13923
rect 19984 13880 20036 13889
rect 12348 13676 12400 13728
rect 15568 13676 15620 13728
rect 15936 13719 15988 13728
rect 15936 13685 15945 13719
rect 15945 13685 15979 13719
rect 15979 13685 15988 13719
rect 15936 13676 15988 13685
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 12992 13472 13044 13524
rect 15936 13472 15988 13524
rect 17868 13472 17920 13524
rect 19156 13472 19208 13524
rect 11980 13336 12032 13388
rect 15200 13336 15252 13388
rect 15384 13336 15436 13388
rect 19340 13336 19392 13388
rect 10140 13268 10192 13320
rect 18052 13311 18104 13320
rect 18052 13277 18061 13311
rect 18061 13277 18095 13311
rect 18095 13277 18104 13311
rect 18052 13268 18104 13277
rect 18144 13311 18196 13320
rect 18144 13277 18153 13311
rect 18153 13277 18187 13311
rect 18187 13277 18196 13311
rect 18144 13268 18196 13277
rect 19432 13268 19484 13320
rect 19800 13311 19852 13320
rect 19800 13277 19809 13311
rect 19809 13277 19843 13311
rect 19843 13277 19852 13311
rect 19800 13268 19852 13277
rect 18512 13200 18564 13252
rect 16488 13132 16540 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 15200 12928 15252 12980
rect 9220 12792 9272 12844
rect 10140 12835 10192 12844
rect 10140 12801 10149 12835
rect 10149 12801 10183 12835
rect 10183 12801 10192 12835
rect 10140 12792 10192 12801
rect 20536 12835 20588 12844
rect 12900 12724 12952 12776
rect 15660 12767 15712 12776
rect 15660 12733 15669 12767
rect 15669 12733 15703 12767
rect 15703 12733 15712 12767
rect 15660 12724 15712 12733
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 10600 12656 10652 12708
rect 12992 12656 13044 12708
rect 11980 12588 12032 12640
rect 14188 12631 14240 12640
rect 14188 12597 14197 12631
rect 14197 12597 14231 12631
rect 14231 12597 14240 12631
rect 14188 12588 14240 12597
rect 16488 12724 16540 12776
rect 19064 12724 19116 12776
rect 20260 12767 20312 12776
rect 20260 12733 20269 12767
rect 20269 12733 20303 12767
rect 20303 12733 20312 12767
rect 20260 12724 20312 12733
rect 18144 12656 18196 12708
rect 16488 12588 16540 12640
rect 17316 12588 17368 12640
rect 18696 12588 18748 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 10508 12384 10560 12436
rect 12348 12384 12400 12436
rect 17868 12384 17920 12436
rect 18144 12427 18196 12436
rect 18144 12393 18153 12427
rect 18153 12393 18187 12427
rect 18187 12393 18196 12427
rect 18144 12384 18196 12393
rect 15108 12316 15160 12368
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 10600 12180 10652 12232
rect 12900 12248 12952 12300
rect 13820 12248 13872 12300
rect 17408 12316 17460 12368
rect 16488 12248 16540 12300
rect 17316 12248 17368 12300
rect 18880 12248 18932 12300
rect 19708 12291 19760 12300
rect 19708 12257 19717 12291
rect 19717 12257 19751 12291
rect 19751 12257 19760 12291
rect 19708 12248 19760 12257
rect 11888 12180 11940 12232
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 20628 12180 20680 12232
rect 9588 12044 9640 12096
rect 14280 12044 14332 12096
rect 15384 12044 15436 12096
rect 19524 12044 19576 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 10600 11883 10652 11892
rect 10600 11849 10609 11883
rect 10609 11849 10643 11883
rect 10643 11849 10652 11883
rect 10600 11840 10652 11849
rect 13912 11840 13964 11892
rect 14648 11883 14700 11892
rect 14648 11849 14657 11883
rect 14657 11849 14691 11883
rect 14691 11849 14700 11883
rect 14648 11840 14700 11849
rect 16672 11840 16724 11892
rect 1216 11704 1268 11756
rect 9220 11679 9272 11688
rect 9220 11645 9229 11679
rect 9229 11645 9263 11679
rect 9263 11645 9272 11679
rect 9220 11636 9272 11645
rect 13820 11704 13872 11756
rect 14648 11704 14700 11756
rect 15108 11747 15160 11756
rect 15108 11713 15117 11747
rect 15117 11713 15151 11747
rect 15151 11713 15160 11747
rect 15108 11704 15160 11713
rect 15384 11704 15436 11756
rect 15476 11704 15528 11756
rect 19340 11704 19392 11756
rect 19524 11747 19576 11756
rect 19524 11713 19533 11747
rect 19533 11713 19567 11747
rect 19567 11713 19576 11747
rect 19524 11704 19576 11713
rect 20812 11704 20864 11756
rect 15568 11636 15620 11688
rect 9864 11568 9916 11620
rect 12624 11568 12676 11620
rect 8300 11500 8352 11552
rect 12716 11500 12768 11552
rect 13452 11543 13504 11552
rect 13452 11509 13461 11543
rect 13461 11509 13495 11543
rect 13495 11509 13504 11543
rect 13452 11500 13504 11509
rect 13544 11543 13596 11552
rect 13544 11509 13553 11543
rect 13553 11509 13587 11543
rect 13587 11509 13596 11543
rect 16672 11543 16724 11552
rect 13544 11500 13596 11509
rect 16672 11509 16681 11543
rect 16681 11509 16715 11543
rect 16715 11509 16724 11543
rect 16672 11500 16724 11509
rect 16856 11500 16908 11552
rect 20168 11500 20220 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 10324 11296 10376 11348
rect 11980 11296 12032 11348
rect 4068 11228 4120 11280
rect 12624 11228 12676 11280
rect 12716 11228 12768 11280
rect 9680 11160 9732 11212
rect 10416 11160 10468 11212
rect 11980 11203 12032 11212
rect 11980 11169 11981 11203
rect 11981 11169 12015 11203
rect 12015 11169 12032 11203
rect 11980 11160 12032 11169
rect 13452 11296 13504 11348
rect 15660 11296 15712 11348
rect 16120 11339 16172 11348
rect 16120 11305 16129 11339
rect 16129 11305 16163 11339
rect 16163 11305 16172 11339
rect 16120 11296 16172 11305
rect 18052 11296 18104 11348
rect 19800 11339 19852 11348
rect 19800 11305 19809 11339
rect 19809 11305 19843 11339
rect 19843 11305 19852 11339
rect 19800 11296 19852 11305
rect 14280 11228 14332 11280
rect 17224 11203 17276 11212
rect 17224 11169 17233 11203
rect 17233 11169 17267 11203
rect 17267 11169 17276 11203
rect 17224 11160 17276 11169
rect 18144 11160 18196 11212
rect 18696 11203 18748 11212
rect 18696 11169 18719 11203
rect 18719 11169 18748 11203
rect 18696 11160 18748 11169
rect 17316 11135 17368 11144
rect 9864 11024 9916 11076
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 12164 11024 12216 11076
rect 11888 10956 11940 11008
rect 15292 10956 15344 11008
rect 16304 10956 16356 11008
rect 19064 10956 19116 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 9864 10795 9916 10804
rect 9864 10761 9873 10795
rect 9873 10761 9907 10795
rect 9907 10761 9916 10795
rect 9864 10752 9916 10761
rect 10784 10795 10836 10804
rect 10784 10761 10793 10795
rect 10793 10761 10827 10795
rect 10827 10761 10836 10795
rect 10784 10752 10836 10761
rect 10876 10752 10928 10804
rect 13820 10795 13872 10804
rect 11704 10616 11756 10668
rect 9128 10548 9180 10600
rect 8944 10480 8996 10532
rect 5080 10412 5132 10464
rect 11796 10548 11848 10600
rect 12624 10480 12676 10532
rect 12900 10480 12952 10532
rect 13820 10761 13829 10795
rect 13829 10761 13863 10795
rect 13863 10761 13872 10795
rect 13820 10752 13872 10761
rect 15476 10795 15528 10804
rect 15476 10761 15485 10795
rect 15485 10761 15519 10795
rect 15519 10761 15528 10795
rect 15476 10752 15528 10761
rect 19432 10752 19484 10804
rect 20628 10752 20680 10804
rect 16304 10684 16356 10736
rect 18144 10616 18196 10668
rect 19064 10616 19116 10668
rect 14188 10548 14240 10600
rect 18604 10548 18656 10600
rect 19800 10480 19852 10532
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 12440 10412 12492 10464
rect 16948 10412 17000 10464
rect 20352 10412 20404 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 9036 10208 9088 10260
rect 10232 10208 10284 10260
rect 11888 10208 11940 10260
rect 14004 10251 14056 10260
rect 14004 10217 14013 10251
rect 14013 10217 14047 10251
rect 14047 10217 14056 10251
rect 14004 10208 14056 10217
rect 17224 10208 17276 10260
rect 18972 10251 19024 10260
rect 18972 10217 18981 10251
rect 18981 10217 19015 10251
rect 19015 10217 19024 10251
rect 18972 10208 19024 10217
rect 11704 10140 11756 10192
rect 13268 10140 13320 10192
rect 11796 10072 11848 10124
rect 16304 10115 16356 10124
rect 1768 10004 1820 10056
rect 8484 10047 8536 10056
rect 8484 10013 8493 10047
rect 8493 10013 8527 10047
rect 8527 10013 8536 10047
rect 8484 10004 8536 10013
rect 8944 10004 8996 10056
rect 10232 10004 10284 10056
rect 11060 10004 11112 10056
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 20812 10140 20864 10192
rect 17316 10072 17368 10124
rect 18880 10115 18932 10124
rect 18880 10081 18889 10115
rect 18889 10081 18923 10115
rect 18923 10081 18932 10115
rect 18880 10072 18932 10081
rect 9220 9936 9272 9988
rect 10416 9868 10468 9920
rect 12624 9979 12676 9988
rect 12624 9945 12633 9979
rect 12633 9945 12667 9979
rect 12667 9945 12676 9979
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 16212 10004 16264 10056
rect 12624 9936 12676 9945
rect 13544 9868 13596 9920
rect 16672 9868 16724 9920
rect 17684 9911 17736 9920
rect 17684 9877 17693 9911
rect 17693 9877 17727 9911
rect 17727 9877 17736 9911
rect 17684 9868 17736 9877
rect 17776 9868 17828 9920
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 8944 9707 8996 9716
rect 8944 9673 8953 9707
rect 8953 9673 8987 9707
rect 8987 9673 8996 9707
rect 8944 9664 8996 9673
rect 11704 9664 11756 9716
rect 20812 9707 20864 9716
rect 20812 9673 20821 9707
rect 20821 9673 20855 9707
rect 20855 9673 20864 9707
rect 20812 9664 20864 9673
rect 9220 9596 9272 9648
rect 12440 9571 12492 9580
rect 12440 9537 12449 9571
rect 12449 9537 12483 9571
rect 12483 9537 12492 9571
rect 12440 9528 12492 9537
rect 8576 9392 8628 9444
rect 12164 9460 12216 9512
rect 13544 9503 13596 9512
rect 13544 9469 13553 9503
rect 13553 9469 13587 9503
rect 13587 9469 13596 9503
rect 13544 9460 13596 9469
rect 15476 9460 15528 9512
rect 11152 9392 11204 9444
rect 17684 9460 17736 9512
rect 18788 9460 18840 9512
rect 19432 9503 19484 9512
rect 19432 9469 19441 9503
rect 19441 9469 19475 9503
rect 19475 9469 19484 9503
rect 19432 9460 19484 9469
rect 20628 9460 20680 9512
rect 16304 9392 16356 9444
rect 16672 9392 16724 9444
rect 11060 9324 11112 9376
rect 11980 9324 12032 9376
rect 12256 9324 12308 9376
rect 12624 9324 12676 9376
rect 14280 9324 14332 9376
rect 17132 9367 17184 9376
rect 17132 9333 17141 9367
rect 17141 9333 17175 9367
rect 17175 9333 17184 9367
rect 17132 9324 17184 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 8484 9120 8536 9172
rect 9772 9163 9824 9172
rect 9772 9129 9781 9163
rect 9781 9129 9815 9163
rect 9815 9129 9824 9163
rect 9772 9120 9824 9129
rect 11244 9120 11296 9172
rect 11796 9120 11848 9172
rect 16948 9120 17000 9172
rect 19248 9163 19300 9172
rect 6552 8984 6604 9036
rect 10140 9027 10192 9036
rect 10140 8993 10149 9027
rect 10149 8993 10183 9027
rect 10183 8993 10192 9027
rect 10140 8984 10192 8993
rect 12072 9052 12124 9104
rect 17132 9052 17184 9104
rect 19248 9129 19257 9163
rect 19257 9129 19291 9163
rect 19291 9129 19300 9163
rect 19248 9120 19300 9129
rect 7012 8959 7064 8968
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 7012 8916 7064 8925
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 10232 8959 10284 8968
rect 8576 8916 8628 8925
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 7288 8848 7340 8900
rect 13452 8984 13504 9036
rect 15292 9027 15344 9036
rect 15292 8993 15301 9027
rect 15301 8993 15335 9027
rect 15335 8993 15344 9027
rect 15292 8984 15344 8993
rect 16396 8984 16448 9036
rect 18880 8984 18932 9036
rect 19248 8984 19300 9036
rect 11060 8916 11112 8968
rect 11152 8848 11204 8900
rect 11980 8916 12032 8968
rect 13728 8916 13780 8968
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 12808 8848 12860 8900
rect 15752 8916 15804 8968
rect 16488 8916 16540 8968
rect 4344 8780 4396 8832
rect 12072 8780 12124 8832
rect 12624 8780 12676 8832
rect 19064 8916 19116 8968
rect 18144 8848 18196 8900
rect 18880 8780 18932 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 2320 8576 2372 8628
rect 7288 8576 7340 8628
rect 8576 8576 8628 8628
rect 11152 8576 11204 8628
rect 12624 8619 12676 8628
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 13728 8576 13780 8628
rect 15292 8576 15344 8628
rect 16764 8576 16816 8628
rect 16488 8508 16540 8560
rect 19432 8576 19484 8628
rect 9220 8440 9272 8492
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 17132 8440 17184 8492
rect 6644 8236 6696 8288
rect 7748 8304 7800 8356
rect 11060 8304 11112 8356
rect 14280 8372 14332 8424
rect 16120 8372 16172 8424
rect 16212 8372 16264 8424
rect 17776 8372 17828 8424
rect 18696 8372 18748 8424
rect 18604 8304 18656 8356
rect 19340 8304 19392 8356
rect 13544 8236 13596 8288
rect 15752 8279 15804 8288
rect 15752 8245 15761 8279
rect 15761 8245 15795 8279
rect 15795 8245 15804 8279
rect 15752 8236 15804 8245
rect 20536 8279 20588 8288
rect 20536 8245 20545 8279
rect 20545 8245 20579 8279
rect 20579 8245 20588 8279
rect 20536 8236 20588 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 7748 8032 7800 8084
rect 11060 8075 11112 8084
rect 11060 8041 11069 8075
rect 11069 8041 11103 8075
rect 11103 8041 11112 8075
rect 11060 8032 11112 8041
rect 10140 7964 10192 8016
rect 10324 7964 10376 8016
rect 16396 8032 16448 8084
rect 18052 8032 18104 8084
rect 11980 7964 12032 8016
rect 12716 7964 12768 8016
rect 16856 7964 16908 8016
rect 18144 8007 18196 8016
rect 18144 7973 18178 8007
rect 18178 7973 18196 8007
rect 18144 7964 18196 7973
rect 6644 7939 6696 7948
rect 6644 7905 6653 7939
rect 6653 7905 6687 7939
rect 6687 7905 6696 7939
rect 6644 7896 6696 7905
rect 7472 7896 7524 7948
rect 9220 7896 9272 7948
rect 10416 7896 10468 7948
rect 15844 7828 15896 7880
rect 12900 7692 12952 7744
rect 13268 7735 13320 7744
rect 13268 7701 13277 7735
rect 13277 7701 13311 7735
rect 13311 7701 13320 7735
rect 13268 7692 13320 7701
rect 16120 7692 16172 7744
rect 16304 7735 16356 7744
rect 16304 7701 16313 7735
rect 16313 7701 16347 7735
rect 16347 7701 16356 7735
rect 16304 7692 16356 7701
rect 20536 7896 20588 7948
rect 16580 7760 16632 7812
rect 17776 7760 17828 7812
rect 18144 7692 18196 7744
rect 19340 7692 19392 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 7104 7531 7156 7540
rect 7104 7497 7113 7531
rect 7113 7497 7147 7531
rect 7147 7497 7156 7531
rect 7104 7488 7156 7497
rect 9312 7488 9364 7540
rect 9588 7488 9640 7540
rect 10232 7488 10284 7540
rect 18696 7488 18748 7540
rect 20168 7488 20220 7540
rect 20720 7488 20772 7540
rect 22100 7488 22152 7540
rect 5816 7352 5868 7404
rect 7748 7395 7800 7404
rect 7012 7284 7064 7336
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 7748 7352 7800 7361
rect 10416 7352 10468 7404
rect 13268 7352 13320 7404
rect 13544 7352 13596 7404
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 10784 7284 10836 7336
rect 12716 7284 12768 7336
rect 7380 7216 7432 7268
rect 11152 7216 11204 7268
rect 11980 7216 12032 7268
rect 16212 7284 16264 7336
rect 17960 7284 18012 7336
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 20536 7284 20588 7336
rect 14372 7216 14424 7268
rect 16580 7216 16632 7268
rect 7564 7191 7616 7200
rect 7564 7157 7573 7191
rect 7573 7157 7607 7191
rect 7607 7157 7616 7191
rect 7564 7148 7616 7157
rect 9772 7191 9824 7200
rect 9772 7157 9781 7191
rect 9781 7157 9815 7191
rect 9815 7157 9824 7191
rect 9772 7148 9824 7157
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 12532 7148 12584 7200
rect 14096 7148 14148 7200
rect 15384 7191 15436 7200
rect 15384 7157 15393 7191
rect 15393 7157 15427 7191
rect 15427 7157 15436 7191
rect 15384 7148 15436 7157
rect 15936 7148 15988 7200
rect 17408 7148 17460 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 7564 6944 7616 6996
rect 12256 6944 12308 6996
rect 12532 6987 12584 6996
rect 12532 6953 12541 6987
rect 12541 6953 12575 6987
rect 12575 6953 12584 6987
rect 12532 6944 12584 6953
rect 17224 6987 17276 6996
rect 17224 6953 17233 6987
rect 17233 6953 17267 6987
rect 17267 6953 17276 6987
rect 17224 6944 17276 6953
rect 19156 6944 19208 6996
rect 7104 6876 7156 6928
rect 12440 6919 12492 6928
rect 12440 6885 12449 6919
rect 12449 6885 12483 6919
rect 12483 6885 12492 6919
rect 14004 6919 14056 6928
rect 12440 6876 12492 6885
rect 14004 6885 14013 6919
rect 14013 6885 14047 6919
rect 14047 6885 14056 6919
rect 14004 6876 14056 6885
rect 15476 6876 15528 6928
rect 16304 6876 16356 6928
rect 20076 6876 20128 6928
rect 7472 6808 7524 6860
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 12164 6808 12216 6860
rect 17316 6851 17368 6860
rect 8208 6740 8260 6792
rect 9864 6740 9916 6792
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 11060 6740 11112 6792
rect 12716 6783 12768 6792
rect 12716 6749 12725 6783
rect 12725 6749 12759 6783
rect 12759 6749 12768 6783
rect 12716 6740 12768 6749
rect 9956 6672 10008 6724
rect 13636 6715 13688 6724
rect 5724 6604 5776 6656
rect 10784 6604 10836 6656
rect 11796 6647 11848 6656
rect 11796 6613 11805 6647
rect 11805 6613 11839 6647
rect 11839 6613 11848 6647
rect 11796 6604 11848 6613
rect 13636 6681 13645 6715
rect 13645 6681 13679 6715
rect 13679 6681 13688 6715
rect 13636 6672 13688 6681
rect 15384 6740 15436 6792
rect 16028 6740 16080 6792
rect 17316 6817 17325 6851
rect 17325 6817 17359 6851
rect 17359 6817 17368 6851
rect 17316 6808 17368 6817
rect 18880 6851 18932 6860
rect 18880 6817 18889 6851
rect 18889 6817 18923 6851
rect 18923 6817 18932 6851
rect 18880 6808 18932 6817
rect 17408 6783 17460 6792
rect 17132 6672 17184 6724
rect 17408 6749 17417 6783
rect 17417 6749 17451 6783
rect 17451 6749 17460 6783
rect 17408 6740 17460 6749
rect 19340 6740 19392 6792
rect 19616 6672 19668 6724
rect 15200 6604 15252 6656
rect 16580 6604 16632 6656
rect 16856 6604 16908 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 8208 6443 8260 6452
rect 8208 6409 8217 6443
rect 8217 6409 8251 6443
rect 8251 6409 8260 6443
rect 8208 6400 8260 6409
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 6644 6264 6696 6316
rect 10784 6196 10836 6248
rect 12624 6400 12676 6452
rect 12716 6400 12768 6452
rect 13912 6400 13964 6452
rect 16948 6400 17000 6452
rect 17040 6400 17092 6452
rect 17684 6400 17736 6452
rect 12164 6332 12216 6384
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 17684 6264 17736 6316
rect 7748 6128 7800 6180
rect 10324 6128 10376 6180
rect 11796 6128 11848 6180
rect 13268 6196 13320 6248
rect 16028 6239 16080 6248
rect 16028 6205 16062 6239
rect 16062 6205 16080 6239
rect 12900 6128 12952 6180
rect 16028 6196 16080 6205
rect 17040 6196 17092 6248
rect 17224 6196 17276 6248
rect 17776 6196 17828 6248
rect 18052 6239 18104 6248
rect 18052 6205 18061 6239
rect 18061 6205 18095 6239
rect 18095 6205 18104 6239
rect 18052 6196 18104 6205
rect 20444 6196 20496 6248
rect 12624 6060 12676 6112
rect 13912 6060 13964 6112
rect 15568 6060 15620 6112
rect 16488 6128 16540 6180
rect 17408 6128 17460 6180
rect 18788 6060 18840 6112
rect 19340 6060 19392 6112
rect 19708 6060 19760 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 7196 5899 7248 5908
rect 7196 5865 7205 5899
rect 7205 5865 7239 5899
rect 7239 5865 7248 5899
rect 7196 5856 7248 5865
rect 10048 5856 10100 5908
rect 10416 5856 10468 5908
rect 15660 5899 15712 5908
rect 6920 5720 6972 5772
rect 10600 5720 10652 5772
rect 10784 5763 10836 5772
rect 10784 5729 10793 5763
rect 10793 5729 10827 5763
rect 10827 5729 10836 5763
rect 10784 5720 10836 5729
rect 11060 5763 11112 5772
rect 11060 5729 11094 5763
rect 11094 5729 11112 5763
rect 11060 5720 11112 5729
rect 15660 5865 15669 5899
rect 15669 5865 15703 5899
rect 15703 5865 15712 5899
rect 15660 5856 15712 5865
rect 18788 5856 18840 5908
rect 15476 5720 15528 5772
rect 16212 5720 16264 5772
rect 16856 5763 16908 5772
rect 16856 5729 16865 5763
rect 16865 5729 16899 5763
rect 16899 5729 16908 5763
rect 16856 5720 16908 5729
rect 19340 5720 19392 5772
rect 6092 5652 6144 5704
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 14188 5652 14240 5704
rect 14372 5652 14424 5704
rect 16488 5652 16540 5704
rect 16672 5584 16724 5636
rect 18052 5652 18104 5704
rect 9864 5559 9916 5568
rect 9864 5525 9873 5559
rect 9873 5525 9907 5559
rect 9907 5525 9916 5559
rect 9864 5516 9916 5525
rect 11796 5516 11848 5568
rect 14924 5516 14976 5568
rect 19432 5516 19484 5568
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 7748 5312 7800 5364
rect 10324 5312 10376 5364
rect 10692 5312 10744 5364
rect 11796 5312 11848 5364
rect 12440 5355 12492 5364
rect 12440 5321 12449 5355
rect 12449 5321 12483 5355
rect 12483 5321 12492 5355
rect 12440 5312 12492 5321
rect 15936 5312 15988 5364
rect 14556 5244 14608 5296
rect 19892 5244 19944 5296
rect 6644 5176 6696 5228
rect 9220 5219 9272 5228
rect 9220 5185 9229 5219
rect 9229 5185 9263 5219
rect 9263 5185 9272 5219
rect 9220 5176 9272 5185
rect 13268 5176 13320 5228
rect 14924 5176 14976 5228
rect 16028 5176 16080 5228
rect 19340 5176 19392 5228
rect 19800 5176 19852 5228
rect 20076 5219 20128 5228
rect 20076 5185 20085 5219
rect 20085 5185 20119 5219
rect 20119 5185 20128 5219
rect 20076 5176 20128 5185
rect 20168 5219 20220 5228
rect 20168 5185 20177 5219
rect 20177 5185 20211 5219
rect 20211 5185 20220 5219
rect 20168 5176 20220 5185
rect 6920 5040 6972 5092
rect 8208 5040 8260 5092
rect 6092 4972 6144 5024
rect 14464 5108 14516 5160
rect 14648 5108 14700 5160
rect 10692 5040 10744 5092
rect 11060 5040 11112 5092
rect 15200 5108 15252 5160
rect 17592 5108 17644 5160
rect 19248 5108 19300 5160
rect 19156 5040 19208 5092
rect 11704 4972 11756 5024
rect 14096 4972 14148 5024
rect 14740 4972 14792 5024
rect 19432 4972 19484 5024
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 7656 4811 7708 4820
rect 7656 4777 7665 4811
rect 7665 4777 7699 4811
rect 7699 4777 7708 4811
rect 7656 4768 7708 4777
rect 8392 4768 8444 4820
rect 10140 4768 10192 4820
rect 11704 4811 11756 4820
rect 11704 4777 11713 4811
rect 11713 4777 11747 4811
rect 11747 4777 11756 4811
rect 11704 4768 11756 4777
rect 11980 4768 12032 4820
rect 17960 4768 18012 4820
rect 7656 4632 7708 4684
rect 4804 4564 4856 4616
rect 12992 4632 13044 4684
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 8392 4564 8444 4616
rect 10692 4564 10744 4616
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 11704 4496 11756 4548
rect 6736 4471 6788 4480
rect 6736 4437 6745 4471
rect 6745 4437 6779 4471
rect 6779 4437 6788 4471
rect 6736 4428 6788 4437
rect 8484 4428 8536 4480
rect 14280 4471 14332 4480
rect 14280 4437 14289 4471
rect 14289 4437 14323 4471
rect 14323 4437 14332 4471
rect 14280 4428 14332 4437
rect 15200 4632 15252 4684
rect 15752 4700 15804 4752
rect 17868 4675 17920 4684
rect 17868 4641 17877 4675
rect 17877 4641 17911 4675
rect 17911 4641 17920 4675
rect 17868 4632 17920 4641
rect 19064 4632 19116 4684
rect 17960 4607 18012 4616
rect 17960 4573 17969 4607
rect 17969 4573 18003 4607
rect 18003 4573 18012 4607
rect 17960 4564 18012 4573
rect 16488 4496 16540 4548
rect 18972 4564 19024 4616
rect 19800 4607 19852 4616
rect 19800 4573 19809 4607
rect 19809 4573 19843 4607
rect 19843 4573 19852 4607
rect 19800 4564 19852 4573
rect 16304 4428 16356 4480
rect 17500 4471 17552 4480
rect 17500 4437 17509 4471
rect 17509 4437 17543 4471
rect 17543 4437 17552 4471
rect 17500 4428 17552 4437
rect 20076 4428 20128 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 8208 4267 8260 4276
rect 8208 4233 8217 4267
rect 8217 4233 8251 4267
rect 8251 4233 8260 4267
rect 8208 4224 8260 4233
rect 16488 4267 16540 4276
rect 16488 4233 16497 4267
rect 16497 4233 16531 4267
rect 16531 4233 16540 4267
rect 16488 4224 16540 4233
rect 19340 4224 19392 4276
rect 20168 4224 20220 4276
rect 6644 4088 6696 4140
rect 8208 4088 8260 4140
rect 9220 4088 9272 4140
rect 2872 3952 2924 4004
rect 9772 4020 9824 4072
rect 10508 4020 10560 4072
rect 10600 4020 10652 4072
rect 12808 4020 12860 4072
rect 18052 4156 18104 4208
rect 14096 4020 14148 4072
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 8576 3952 8628 4004
rect 16120 4088 16172 4140
rect 17224 4088 17276 4140
rect 15752 4020 15804 4072
rect 16396 4020 16448 4072
rect 15384 3995 15436 4004
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 7196 3884 7248 3936
rect 8760 3884 8812 3936
rect 10232 3884 10284 3936
rect 11244 3927 11296 3936
rect 11244 3893 11253 3927
rect 11253 3893 11287 3927
rect 11287 3893 11296 3927
rect 11244 3884 11296 3893
rect 12440 3884 12492 3936
rect 13544 3927 13596 3936
rect 13544 3893 13553 3927
rect 13553 3893 13587 3927
rect 13587 3893 13596 3927
rect 13544 3884 13596 3893
rect 15384 3961 15418 3995
rect 15418 3961 15436 3995
rect 15384 3952 15436 3961
rect 15476 3952 15528 4004
rect 16764 3952 16816 4004
rect 17132 3952 17184 4004
rect 19340 3995 19392 4004
rect 19340 3961 19374 3995
rect 19374 3961 19392 3995
rect 19340 3952 19392 3961
rect 17592 3884 17644 3936
rect 19984 3884 20036 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 5632 3680 5684 3732
rect 6460 3680 6512 3732
rect 7196 3680 7248 3732
rect 7564 3680 7616 3732
rect 8484 3723 8536 3732
rect 8484 3689 8493 3723
rect 8493 3689 8527 3723
rect 8527 3689 8536 3723
rect 8484 3680 8536 3689
rect 6000 3612 6052 3664
rect 9680 3680 9732 3732
rect 13360 3680 13412 3732
rect 15476 3680 15528 3732
rect 15752 3680 15804 3732
rect 17500 3680 17552 3732
rect 17592 3680 17644 3732
rect 19984 3680 20036 3732
rect 9220 3612 9272 3664
rect 10600 3612 10652 3664
rect 11244 3612 11296 3664
rect 5816 3587 5868 3596
rect 5816 3553 5825 3587
rect 5825 3553 5859 3587
rect 5859 3553 5868 3587
rect 5816 3544 5868 3553
rect 8208 3544 8260 3596
rect 8392 3587 8444 3596
rect 8392 3553 8401 3587
rect 8401 3553 8435 3587
rect 8435 3553 8444 3587
rect 8392 3544 8444 3553
rect 8576 3544 8628 3596
rect 8852 3544 8904 3596
rect 9312 3476 9364 3528
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 3332 3408 3384 3460
rect 4804 3408 4856 3460
rect 4988 3451 5040 3460
rect 4988 3417 4997 3451
rect 4997 3417 5031 3451
rect 5031 3417 5040 3451
rect 4988 3408 5040 3417
rect 5540 3340 5592 3392
rect 8760 3340 8812 3392
rect 12256 3408 12308 3460
rect 11980 3383 12032 3392
rect 11980 3349 11989 3383
rect 11989 3349 12023 3383
rect 12023 3349 12032 3383
rect 16764 3612 16816 3664
rect 16948 3612 17000 3664
rect 14280 3544 14332 3596
rect 15660 3544 15712 3596
rect 17132 3544 17184 3596
rect 19432 3587 19484 3596
rect 19432 3553 19441 3587
rect 19441 3553 19475 3587
rect 19475 3553 19484 3587
rect 19432 3544 19484 3553
rect 20352 3544 20404 3596
rect 21548 3544 21600 3596
rect 12808 3519 12860 3528
rect 12808 3485 12817 3519
rect 12817 3485 12851 3519
rect 12851 3485 12860 3519
rect 12808 3476 12860 3485
rect 16304 3519 16356 3528
rect 16304 3485 16313 3519
rect 16313 3485 16347 3519
rect 16347 3485 16356 3519
rect 16304 3476 16356 3485
rect 16396 3476 16448 3528
rect 14096 3408 14148 3460
rect 11980 3340 12032 3349
rect 12992 3340 13044 3392
rect 19708 3408 19760 3460
rect 18604 3383 18656 3392
rect 18604 3349 18613 3383
rect 18613 3349 18647 3383
rect 18647 3349 18656 3383
rect 18604 3340 18656 3349
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 9312 3179 9364 3188
rect 3884 3068 3936 3120
rect 9312 3145 9321 3179
rect 9321 3145 9355 3179
rect 9355 3145 9364 3179
rect 9312 3136 9364 3145
rect 10968 3136 11020 3188
rect 12532 3136 12584 3188
rect 15200 3136 15252 3188
rect 15660 3179 15712 3188
rect 15660 3145 15669 3179
rect 15669 3145 15703 3179
rect 15703 3145 15712 3179
rect 15660 3136 15712 3145
rect 15752 3136 15804 3188
rect 6736 3000 6788 3052
rect 10508 3068 10560 3120
rect 11060 3000 11112 3052
rect 11244 3000 11296 3052
rect 11888 3068 11940 3120
rect 12992 3000 13044 3052
rect 13544 3068 13596 3120
rect 17960 3136 18012 3188
rect 19616 3179 19668 3188
rect 19616 3145 19625 3179
rect 19625 3145 19659 3179
rect 19659 3145 19668 3179
rect 19616 3136 19668 3145
rect 13636 3000 13688 3052
rect 13728 3000 13780 3052
rect 14280 3000 14332 3052
rect 7380 2932 7432 2984
rect 15936 2932 15988 2984
rect 16488 3000 16540 3052
rect 17408 3000 17460 3052
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 18052 2932 18104 2984
rect 18788 2932 18840 2984
rect 19432 3068 19484 3120
rect 19708 3068 19760 3120
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 20168 3043 20220 3052
rect 20168 3009 20177 3043
rect 20177 3009 20211 3043
rect 20211 3009 20220 3043
rect 20168 3000 20220 3009
rect 20260 2932 20312 2984
rect 204 2796 256 2848
rect 5540 2796 5592 2848
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 8668 2864 8720 2916
rect 11980 2864 12032 2916
rect 10232 2796 10284 2848
rect 11152 2839 11204 2848
rect 11152 2805 11161 2839
rect 11161 2805 11195 2839
rect 11195 2805 11204 2839
rect 11152 2796 11204 2805
rect 12992 2839 13044 2848
rect 12992 2805 13001 2839
rect 13001 2805 13035 2839
rect 13035 2805 13044 2839
rect 14648 2864 14700 2916
rect 18144 2864 18196 2916
rect 19892 2864 19944 2916
rect 12992 2796 13044 2805
rect 14464 2839 14516 2848
rect 14464 2805 14473 2839
rect 14473 2805 14507 2839
rect 14507 2805 14516 2839
rect 14464 2796 14516 2805
rect 15200 2796 15252 2848
rect 16212 2796 16264 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 8392 2592 8444 2644
rect 10232 2635 10284 2644
rect 10232 2601 10241 2635
rect 10241 2601 10275 2635
rect 10275 2601 10284 2635
rect 10232 2592 10284 2601
rect 12992 2592 13044 2644
rect 17868 2592 17920 2644
rect 8208 2524 8260 2576
rect 11704 2524 11756 2576
rect 7012 2499 7064 2508
rect 7012 2465 7021 2499
rect 7021 2465 7055 2499
rect 7055 2465 7064 2499
rect 7012 2456 7064 2465
rect 11244 2456 11296 2508
rect 13452 2499 13504 2508
rect 13452 2465 13461 2499
rect 13461 2465 13495 2499
rect 13495 2465 13504 2499
rect 13452 2456 13504 2465
rect 15384 2524 15436 2576
rect 17408 2524 17460 2576
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 8760 2388 8812 2440
rect 10508 2431 10560 2440
rect 10508 2397 10517 2431
rect 10517 2397 10551 2431
rect 10551 2397 10560 2431
rect 10508 2388 10560 2397
rect 13728 2431 13780 2440
rect 13728 2397 13737 2431
rect 13737 2397 13771 2431
rect 13771 2397 13780 2431
rect 13728 2388 13780 2397
rect 16672 2456 16724 2508
rect 17040 2499 17092 2508
rect 17040 2465 17049 2499
rect 17049 2465 17083 2499
rect 17083 2465 17092 2499
rect 17040 2456 17092 2465
rect 17132 2431 17184 2440
rect 17132 2397 17141 2431
rect 17141 2397 17175 2431
rect 17175 2397 17184 2431
rect 17132 2388 17184 2397
rect 17960 2456 18012 2508
rect 18972 2456 19024 2508
rect 19248 2456 19300 2508
rect 5724 2320 5776 2372
rect 7196 2295 7248 2304
rect 7196 2261 7205 2295
rect 7205 2261 7239 2295
rect 7239 2261 7248 2295
rect 7196 2252 7248 2261
rect 11152 2320 11204 2372
rect 19524 2431 19576 2440
rect 19524 2397 19533 2431
rect 19533 2397 19567 2431
rect 19567 2397 19576 2431
rect 19524 2388 19576 2397
rect 20168 2388 20220 2440
rect 11704 2252 11756 2304
rect 13544 2252 13596 2304
rect 17960 2252 18012 2304
rect 19064 2295 19116 2304
rect 19064 2261 19073 2295
rect 19073 2261 19107 2295
rect 19107 2261 19116 2295
rect 19064 2252 19116 2261
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 7196 2048 7248 2100
rect 20444 2048 20496 2100
rect 9772 1980 9824 2032
rect 19524 1980 19576 2032
rect 7012 1912 7064 1964
rect 14004 1912 14056 1964
rect 19064 1912 19116 1964
rect 17132 1844 17184 1896
rect 17316 1844 17368 1896
rect 13452 1776 13504 1828
rect 18972 1776 19024 1828
rect 18696 1708 18748 1760
rect 9864 1640 9916 1692
rect 18328 1640 18380 1692
rect 12164 1096 12216 1148
rect 17776 1096 17828 1148
rect 19432 552 19484 604
rect 19708 552 19760 604
<< metal2 >>
rect 2870 22520 2926 23000
rect 8574 22522 8630 23000
rect 8312 22520 8630 22522
rect 14370 22520 14426 23000
rect 18050 22672 18106 22681
rect 18050 22607 18106 22616
rect 2884 20058 2912 22520
rect 8312 22494 8616 22520
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4816 19514 4844 19654
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 662 12200 718 12209
rect 662 12135 718 12144
rect 204 2848 256 2854
rect 204 2790 256 2796
rect 216 480 244 2790
rect 676 480 704 12135
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 1216 11756 1268 11762
rect 1216 11698 1268 11704
rect 1228 480 1256 11698
rect 4066 11520 4122 11529
rect 4066 11455 4122 11464
rect 4080 11286 4108 11455
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1780 480 1808 9998
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2332 480 2360 8570
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2884 480 2912 3946
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3344 480 3372 3402
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 3896 480 3924 3062
rect 4356 1442 4384 8774
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4816 3466 4844 4558
rect 4986 3496 5042 3505
rect 4804 3460 4856 3466
rect 4986 3431 4988 3440
rect 4804 3402 4856 3408
rect 5040 3431 5042 3440
rect 4988 3402 5040 3408
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 5092 2632 5120 10406
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 6322 5764 6598
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5552 2854 5580 3334
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5000 2604 5120 2632
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4356 1414 4476 1442
rect 4448 480 4476 1414
rect 5000 480 5028 2604
rect 5644 1034 5672 3674
rect 5736 2378 5764 3878
rect 5828 3602 5856 7346
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6104 5030 6132 5646
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6458 4040 6514 4049
rect 6458 3975 6514 3984
rect 6472 3738 6500 3975
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5814 2952 5870 2961
rect 5814 2887 5870 2896
rect 5828 2854 5856 2887
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5552 1006 5672 1034
rect 5552 480 5580 1006
rect 6012 480 6040 3606
rect 6564 480 6592 8978
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 7954 6684 8230
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6656 6322 6684 7890
rect 7024 7342 7052 8910
rect 7116 7546 7144 14894
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6656 5234 6684 6258
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6656 4146 6684 5170
rect 6932 5098 6960 5714
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6656 3074 6684 4082
rect 6748 3641 6776 4422
rect 6734 3632 6790 3641
rect 6734 3567 6790 3576
rect 7010 3224 7066 3233
rect 7010 3159 7012 3168
rect 7064 3159 7066 3168
rect 7012 3130 7064 3136
rect 6656 3058 6776 3074
rect 6656 3052 6788 3058
rect 6656 3046 6736 3052
rect 6736 2994 6788 3000
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7024 1970 7052 2450
rect 7012 1964 7064 1970
rect 7012 1906 7064 1912
rect 7116 480 7144 6870
rect 7208 5914 7236 14418
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7300 8634 7328 8842
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7208 3738 7236 3878
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7392 2990 7420 7210
rect 7484 6866 7512 7890
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 7002 7604 7142
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7668 5794 7696 14282
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8312 11558 8340 22494
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8944 10532 8996 10538
rect 8944 10474 8996 10480
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 8956 10062 8984 10474
rect 9048 10266 9076 14894
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9232 11694 9260 12786
rect 9586 12200 9642 12209
rect 9586 12135 9642 12144
rect 9600 12102 9628 12135
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9128 10600 9180 10606
rect 9232 10588 9260 11630
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9180 10560 9260 10588
rect 9128 10542 9180 10548
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8496 9178 8524 9998
rect 8956 9722 8984 9998
rect 9232 9994 9260 10560
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 9232 9654 9260 9930
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8588 8974 8616 9386
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8588 8634 8616 8910
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 9232 8498 9260 9590
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7760 8090 7788 8298
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7760 7410 7788 8026
rect 9232 7954 9260 8434
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8220 6458 8248 6734
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7576 5766 7696 5794
rect 7576 3738 7604 5766
rect 7760 5710 7788 6122
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7668 4826 7696 5646
rect 7760 5370 7788 5646
rect 7748 5364 7800 5370
rect 7748 5306 7800 5312
rect 9232 5234 9260 7890
rect 9324 7546 9628 7562
rect 9312 7540 9640 7546
rect 9364 7534 9588 7540
rect 9312 7482 9364 7488
rect 9588 7482 9640 7488
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7208 2106 7236 2246
rect 7196 2100 7248 2106
rect 7196 2042 7248 2048
rect 7668 480 7696 4626
rect 8220 4622 8248 5034
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8404 4622 8432 4762
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8220 4282 8248 4558
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 8220 3602 8248 4082
rect 8496 3738 8524 4422
rect 9232 4146 9260 5170
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8588 3602 8616 3946
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8392 3596 8444 3602
rect 8392 3538 8444 3544
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 8404 2650 8432 3538
rect 8772 3398 8800 3878
rect 9692 3738 9720 11154
rect 9784 9178 9812 18770
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9876 11082 9904 11562
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9876 10810 9904 11018
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9784 4078 9812 7142
rect 9876 6798 9904 7142
rect 9864 6792 9916 6798
rect 9862 6760 9864 6769
rect 9916 6760 9918 6769
rect 9968 6730 9996 18158
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10152 12850 10180 13262
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10244 10266 10272 17002
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10520 12442 10548 15506
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10612 12238 10640 12650
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10336 11354 10364 12174
rect 10612 11898 10640 12174
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10230 10160 10286 10169
rect 10230 10095 10286 10104
rect 10244 10062 10272 10095
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10428 9926 10456 11154
rect 10796 10810 10824 19246
rect 14016 18970 14044 19246
rect 14384 19242 14412 22520
rect 17774 21720 17830 21729
rect 17774 21655 17830 21664
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 14372 19236 14424 19242
rect 14372 19178 14424 19184
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14004 18964 14056 18970
rect 14004 18906 14056 18912
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 10968 14000 11020 14006
rect 10968 13942 11020 13948
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10152 8022 10180 8978
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10244 7546 10272 8910
rect 10324 8016 10376 8022
rect 10324 7958 10376 7964
rect 10782 7984 10838 7993
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10336 7426 10364 7958
rect 10416 7948 10468 7954
rect 10782 7919 10838 7928
rect 10416 7890 10468 7896
rect 10244 7398 10364 7426
rect 10428 7410 10456 7890
rect 10416 7404 10468 7410
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 9862 6695 9918 6704
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 10060 5914 10088 6802
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8864 3233 8892 3538
rect 8850 3224 8906 3233
rect 8850 3159 8906 3168
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 8220 480 8248 2518
rect 8680 2446 8708 2858
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8772 480 8800 2382
rect 9232 480 9260 3606
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9324 3194 9352 3470
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9772 2032 9824 2038
rect 9772 1974 9824 1980
rect 9784 480 9812 1974
rect 9876 1698 9904 5510
rect 10152 4826 10180 6734
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10244 3942 10272 7398
rect 10416 7346 10468 7352
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 6186 10364 6734
rect 10428 6458 10456 7346
rect 10796 7342 10824 7919
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10796 6254 10824 6598
rect 10784 6248 10836 6254
rect 10598 6216 10654 6225
rect 10324 6180 10376 6186
rect 10784 6190 10836 6196
rect 10598 6151 10654 6160
rect 10324 6122 10376 6128
rect 10336 5370 10364 6122
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10428 2904 10456 5850
rect 10612 5778 10640 6151
rect 10796 5778 10824 6190
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10704 5098 10732 5306
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10704 4622 10732 5034
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10520 3126 10548 4014
rect 10612 3670 10640 4014
rect 10600 3664 10652 3670
rect 10796 3618 10824 5714
rect 10600 3606 10652 3612
rect 10704 3590 10824 3618
rect 10600 3528 10652 3534
rect 10704 3482 10732 3590
rect 10652 3476 10732 3482
rect 10600 3470 10732 3476
rect 10612 3454 10732 3470
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10336 2876 10456 2904
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10244 2650 10272 2790
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 9864 1692 9916 1698
rect 9864 1634 9916 1640
rect 10336 480 10364 2876
rect 10520 2446 10548 3062
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10888 480 10916 10746
rect 10980 3194 11008 13942
rect 12544 13870 12572 14350
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11992 12646 12020 13330
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11992 12238 12020 12582
rect 12360 12442 12388 13670
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12636 12356 12664 17070
rect 13004 16726 13032 17682
rect 13280 17202 13308 18158
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 12992 16720 13044 16726
rect 12992 16662 13044 16668
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12728 14074 12756 16594
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13004 13530 13032 13874
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12544 12328 12664 12356
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11900 11098 11928 12174
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11992 11218 12020 11290
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11900 11070 12020 11098
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 11072 9382 11100 9998
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8362 11100 8910
rect 11164 8906 11192 9386
rect 11256 9178 11284 10406
rect 11716 10198 11744 10610
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11808 10441 11836 10542
rect 11794 10432 11850 10441
rect 11794 10367 11850 10376
rect 11900 10266 11928 10950
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11716 9722 11744 10134
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11808 9178 11836 10066
rect 11992 9466 12020 11070
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12176 9518 12204 11018
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 9586 12480 10406
rect 12544 9602 12572 12328
rect 12912 12306 12940 12718
rect 13004 12714 13032 13466
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12636 11286 12664 11562
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12728 11286 12756 11494
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 12912 10538 12940 12242
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13464 11354 13492 11494
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 12636 9994 12664 10474
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12440 9580 12492 9586
rect 12544 9574 12664 9602
rect 12440 9522 12492 9528
rect 11900 9438 12020 9466
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11152 8900 11204 8906
rect 11152 8842 11204 8848
rect 11164 8634 11192 8842
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 11072 8090 11100 8298
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11072 5778 11100 6734
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 11072 3058 11100 5034
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11164 2938 11192 7210
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11808 6186 11836 6598
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11808 5370 11836 5510
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4826 11744 4966
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11704 4548 11756 4554
rect 11704 4490 11756 4496
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11256 3670 11284 3878
rect 11244 3664 11296 3670
rect 11244 3606 11296 3612
rect 11256 3058 11284 3606
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11164 2910 11284 2938
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 11164 2378 11192 2790
rect 11256 2514 11284 2910
rect 11716 2582 11744 4490
rect 11900 4049 11928 9438
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11992 8974 12020 9318
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11992 8022 12020 8910
rect 12084 8838 12112 9046
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11980 7268 12032 7274
rect 11980 7210 12032 7216
rect 11992 4826 12020 7210
rect 12176 6866 12204 9454
rect 12636 9382 12664 9574
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12268 7002 12296 9318
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 8634 12664 8774
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12728 7342 12756 7958
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 7002 12572 7142
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11886 4040 11942 4049
rect 11886 3975 11942 3984
rect 11992 3398 12020 4558
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11716 1170 11744 2246
rect 11440 1142 11744 1170
rect 11440 480 11468 1142
rect 11900 480 11928 3062
rect 11992 2922 12020 3334
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 12176 1154 12204 6326
rect 12452 5370 12480 6870
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12728 6458 12756 6734
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12636 6118 12664 6394
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12820 4078 12848 8842
rect 12912 7750 12940 10474
rect 13268 10192 13320 10198
rect 13266 10160 13268 10169
rect 13320 10160 13322 10169
rect 13266 10095 13322 10104
rect 13556 9926 13584 11494
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 12912 6186 12940 7686
rect 13280 7410 13308 7686
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13280 6254 13308 7346
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12912 5930 12940 6122
rect 12912 5902 13032 5930
rect 13004 4690 13032 5902
rect 13280 5234 13308 6190
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12256 3460 12308 3466
rect 12256 3402 12308 3408
rect 12268 3097 12296 3402
rect 12254 3088 12310 3097
rect 12254 3023 12310 3032
rect 12164 1148 12216 1154
rect 12164 1090 12216 1096
rect 12452 480 12480 3878
rect 12808 3528 12860 3534
rect 13004 3482 13032 4626
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 12860 3476 13032 3482
rect 12808 3470 13032 3476
rect 12820 3454 13032 3470
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12544 3097 12572 3130
rect 12530 3088 12586 3097
rect 13004 3058 13032 3334
rect 12530 3023 12586 3032
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 13004 2650 13032 2790
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13372 1306 13400 3674
rect 13464 2514 13492 8978
rect 13556 8498 13584 9454
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13556 8294 13584 8434
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13556 7410 13584 8230
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13648 6730 13676 14962
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13832 11762 13860 12242
rect 13924 11898 13952 18770
rect 14200 15858 14228 19110
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14200 15830 14412 15858
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13832 10810 13860 11698
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 14200 10606 14228 12582
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14292 11286 14320 12038
rect 14280 11280 14332 11286
rect 14280 11222 14332 11228
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14002 10432 14058 10441
rect 14002 10367 14058 10376
rect 14016 10266 14044 10367
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14200 10062 14228 10542
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14292 8974 14320 9318
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 13740 8634 13768 8910
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 14292 8430 14320 8910
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14384 7274 14412 15830
rect 14752 15638 14780 16594
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 14740 15632 14792 15638
rect 14740 15574 14792 15580
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14660 11898 14688 13806
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 15212 13394 15240 18906
rect 15856 18766 15884 19926
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15212 12986 15240 13330
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 15120 11762 15148 12310
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 14462 9072 14518 9081
rect 14462 9007 14518 9016
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14004 6928 14056 6934
rect 14004 6870 14056 6876
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13924 6118 13952 6394
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 3126 13584 3878
rect 13634 3224 13690 3233
rect 13634 3159 13690 3168
rect 13544 3120 13596 3126
rect 13544 3062 13596 3068
rect 13648 3058 13676 3159
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 13464 1834 13492 2450
rect 13740 2446 13768 2994
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13452 1828 13504 1834
rect 13452 1770 13504 1776
rect 13004 1278 13400 1306
rect 13004 480 13032 1278
rect 13556 480 13584 2246
rect 14016 1970 14044 6870
rect 14108 5692 14136 7142
rect 14384 5710 14412 7210
rect 14188 5704 14240 5710
rect 14108 5664 14188 5692
rect 14108 5030 14136 5664
rect 14188 5646 14240 5652
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14476 5166 14504 9007
rect 14556 5296 14608 5302
rect 14556 5238 14608 5244
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14108 4078 14136 4966
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14096 4072 14148 4078
rect 14094 4040 14096 4049
rect 14148 4040 14150 4049
rect 14094 3975 14150 3984
rect 14292 3602 14320 4422
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14096 3460 14148 3466
rect 14096 3402 14148 3408
rect 14004 1964 14056 1970
rect 14004 1906 14056 1912
rect 14108 480 14136 3402
rect 14292 3058 14320 3538
rect 14462 3088 14518 3097
rect 14280 3052 14332 3058
rect 14462 3023 14518 3032
rect 14280 2994 14332 3000
rect 14476 2854 14504 3023
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14568 480 14596 5238
rect 14660 5166 14688 11698
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15304 11014 15332 14350
rect 16592 14074 16620 18770
rect 16672 16720 16724 16726
rect 16672 16662 16724 16668
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15396 12102 15424 13330
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15396 11762 15424 12038
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15488 10810 15516 11698
rect 15580 11694 15608 13670
rect 15948 13530 15976 13670
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 16500 13190 16528 13874
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16500 12782 16528 13126
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15672 11354 15700 12718
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 16500 12306 16528 12582
rect 16488 12300 16540 12306
rect 16488 12242 16540 12248
rect 16684 11898 16712 16662
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17328 13938 17356 14418
rect 17788 14278 17816 21655
rect 17960 20324 18012 20330
rect 17960 20266 18012 20272
rect 17972 19310 18000 20266
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 17958 18864 18014 18873
rect 17958 18799 18014 18808
rect 17972 18426 18000 18799
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17972 14958 18000 15982
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 18064 14770 18092 22607
rect 20074 22520 20130 23000
rect 18970 22264 19026 22273
rect 18970 22199 19026 22208
rect 18786 20768 18842 20777
rect 18282 20700 18578 20720
rect 18786 20703 18842 20712
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18800 20058 18828 20703
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18616 18902 18644 19858
rect 18984 19174 19012 22199
rect 19062 21312 19118 21321
rect 19062 21247 19118 21256
rect 19076 20602 19104 21247
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 19800 20392 19852 20398
rect 19800 20334 19852 20340
rect 19614 19408 19670 19417
rect 19614 19343 19670 19352
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18604 18896 18656 18902
rect 18604 18838 18656 18844
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18970 18048 19026 18057
rect 18970 17983 19026 17992
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18984 17338 19012 17983
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18788 17128 18840 17134
rect 18602 17096 18658 17105
rect 18788 17070 18840 17076
rect 18602 17031 18658 17040
rect 18616 16794 18644 17031
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18800 16726 18828 17070
rect 18788 16720 18840 16726
rect 18788 16662 18840 16668
rect 18602 16552 18658 16561
rect 18602 16487 18658 16496
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18616 16250 18644 16487
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18786 16144 18842 16153
rect 18786 16079 18842 16088
rect 18144 15972 18196 15978
rect 18144 15914 18196 15920
rect 17972 14742 18092 14770
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17880 13530 17908 14350
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17866 13288 17922 13297
rect 17866 13223 17922 13232
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17328 12306 17356 12582
rect 17880 12442 17908 13223
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15488 9518 15516 10746
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15304 8634 15332 8978
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15764 8294 15792 8910
rect 16132 8430 16160 11290
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16316 10742 16344 10950
rect 16304 10736 16356 10742
rect 16304 10678 16356 10684
rect 16316 10130 16344 10678
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16224 8430 16252 9998
rect 16316 9450 16344 10066
rect 16684 9926 16712 11494
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 15396 6798 15424 7142
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14936 5234 14964 5510
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 15212 5166 15240 6598
rect 15488 5778 15516 6870
rect 15658 6760 15714 6769
rect 15658 6695 15714 6704
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 14660 2922 14688 5102
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14648 2916 14700 2922
rect 14648 2858 14700 2864
rect 14752 1442 14780 4966
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15108 4072 15160 4078
rect 15212 4060 15240 4626
rect 15160 4032 15240 4060
rect 15108 4014 15160 4020
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15476 4004 15528 4010
rect 15476 3946 15528 3952
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15212 2854 15240 3130
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 15396 2582 15424 3946
rect 15488 3738 15516 3946
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15580 3074 15608 6054
rect 15672 5914 15700 6695
rect 15764 6322 15792 8230
rect 16408 8090 16436 8978
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16500 8566 16528 8910
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 16500 7834 16528 8502
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15764 4758 15792 6258
rect 15752 4752 15804 4758
rect 15752 4694 15804 4700
rect 15764 4078 15792 4694
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15672 3194 15700 3538
rect 15764 3194 15792 3674
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15856 3074 15884 7822
rect 16500 7818 16620 7834
rect 16500 7812 16632 7818
rect 16500 7806 16580 7812
rect 16580 7754 16632 7760
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15948 5370 15976 7142
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16040 6254 16068 6734
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 16040 5234 16068 6190
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16132 4146 16160 7686
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 16224 5778 16252 7278
rect 16316 6934 16344 7686
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16592 6662 16620 7210
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16488 6180 16540 6186
rect 16488 6122 16540 6128
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16500 5710 16528 6122
rect 16684 5794 16712 9386
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16592 5766 16712 5794
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16488 4548 16540 4554
rect 16488 4490 16540 4496
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16316 3534 16344 4422
rect 16500 4282 16528 4490
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16408 3534 16436 4014
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 15580 3046 15700 3074
rect 15856 3046 15976 3074
rect 16500 3058 16528 4218
rect 16592 3233 16620 5766
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16578 3224 16634 3233
rect 16578 3159 16634 3168
rect 15384 2576 15436 2582
rect 15384 2518 15436 2524
rect 14752 1414 15148 1442
rect 15120 480 15148 1414
rect 15672 480 15700 3046
rect 15948 2990 15976 3046
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 16224 480 16252 2790
rect 16684 2514 16712 5578
rect 16776 4010 16804 8570
rect 16868 8022 16896 11494
rect 17224 11212 17276 11218
rect 17224 11154 17276 11160
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16960 9178 16988 10406
rect 17236 10266 17264 11154
rect 17328 11150 17356 12242
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 17144 9110 17172 9318
rect 17132 9104 17184 9110
rect 17132 9046 17184 9052
rect 17144 8498 17172 9046
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 16856 8016 16908 8022
rect 16856 7958 16908 7964
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16868 5778 16896 6598
rect 17052 6458 17080 7346
rect 17236 7002 17264 10202
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17132 6724 17184 6730
rect 17132 6666 17184 6672
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16960 3670 16988 6394
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16948 3664 17000 3670
rect 16948 3606 17000 3612
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 16776 480 16804 3606
rect 17052 2553 17080 6190
rect 17144 4010 17172 6666
rect 17236 6254 17264 6938
rect 17328 6866 17356 10066
rect 17420 7206 17448 12310
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17696 9518 17724 9862
rect 17684 9512 17736 9518
rect 17498 9480 17554 9489
rect 17684 9454 17736 9460
rect 17498 9415 17554 9424
rect 17512 7426 17540 9415
rect 17788 8430 17816 9862
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17512 7398 17724 7426
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17132 4004 17184 4010
rect 17132 3946 17184 3952
rect 17144 3602 17172 3946
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 17038 2544 17094 2553
rect 17038 2479 17040 2488
rect 17092 2479 17094 2488
rect 17040 2450 17092 2456
rect 17052 2419 17080 2450
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17144 1902 17172 2382
rect 17132 1896 17184 1902
rect 17132 1838 17184 1844
rect 17236 1034 17264 4082
rect 17328 1902 17356 6802
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17420 6186 17448 6734
rect 17696 6610 17724 7398
rect 17604 6582 17724 6610
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 17604 5166 17632 6582
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17696 6322 17724 6394
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17788 6254 17816 7754
rect 17972 7342 18000 14742
rect 18156 14550 18184 15914
rect 18800 15706 18828 16079
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18616 14890 18644 15506
rect 19062 15192 19118 15201
rect 19062 15127 19064 15136
rect 19116 15127 19118 15136
rect 19064 15098 19116 15104
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18604 14884 18656 14890
rect 18604 14826 18656 14832
rect 18696 14884 18748 14890
rect 18696 14826 18748 14832
rect 18144 14544 18196 14550
rect 18144 14486 18196 14492
rect 18708 14482 18736 14826
rect 18892 14550 18920 14894
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18512 13864 18564 13870
rect 18616 13841 18644 14214
rect 18512 13806 18564 13812
rect 18602 13832 18658 13841
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18064 11354 18092 13262
rect 18156 12714 18184 13262
rect 18524 13258 18552 13806
rect 18602 13767 18658 13776
rect 19076 13410 19104 14758
rect 19168 13530 19196 19246
rect 19628 18426 19656 19343
rect 19812 18902 19840 20334
rect 20088 19854 20116 22520
rect 20166 20360 20222 20369
rect 20166 20295 20222 20304
rect 20180 20262 20208 20295
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20076 19848 20128 19854
rect 19890 19816 19946 19825
rect 20076 19790 20128 19796
rect 19890 19751 19892 19760
rect 19944 19751 19946 19760
rect 19892 19722 19944 19728
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 19800 18896 19852 18902
rect 19800 18838 19852 18844
rect 20732 18578 20760 19450
rect 20640 18550 20760 18578
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 20640 18306 20668 18550
rect 20718 18456 20774 18465
rect 20718 18391 20720 18400
rect 20772 18391 20774 18400
rect 20720 18362 20772 18368
rect 20640 18278 20760 18306
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 19892 17536 19944 17542
rect 19890 17504 19892 17513
rect 19944 17504 19946 17513
rect 19890 17439 19946 17448
rect 20548 17202 20576 18158
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 19260 15609 19288 15846
rect 19246 15600 19302 15609
rect 19246 15535 19302 15544
rect 19984 15564 20036 15570
rect 19984 15506 20036 15512
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19904 14657 19932 15302
rect 19890 14648 19946 14657
rect 19890 14583 19946 14592
rect 19996 13938 20024 15506
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19076 13382 19196 13410
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18602 12880 18658 12889
rect 18602 12815 18658 12824
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 18156 12442 18184 12650
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18156 10674 18184 11154
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18144 10668 18196 10674
rect 18144 10610 18196 10616
rect 18616 10606 18644 12815
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18708 11218 18736 12582
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18786 11928 18842 11937
rect 18786 11863 18842 11872
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 18694 10976 18750 10985
rect 18694 10911 18750 10920
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17972 6338 18000 7278
rect 18064 6769 18092 8026
rect 18156 8022 18184 8842
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18708 8430 18736 10911
rect 18800 9518 18828 11863
rect 18892 10130 18920 12242
rect 18970 11384 19026 11393
rect 18970 11319 19026 11328
rect 18984 10266 19012 11319
rect 19076 11014 19104 12718
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 19076 10674 19104 10950
rect 19064 10668 19116 10674
rect 19064 10610 19116 10616
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18892 9042 18920 10066
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18786 8664 18842 8673
rect 18786 8599 18842 8608
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18144 8016 18196 8022
rect 18144 7958 18196 7964
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18156 7177 18184 7686
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18142 7168 18198 7177
rect 18142 7103 18198 7112
rect 18050 6760 18106 6769
rect 18050 6695 18106 6704
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 17972 6310 18184 6338
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 18052 6248 18104 6254
rect 18052 6190 18104 6196
rect 18064 5710 18092 6190
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 17958 5264 18014 5273
rect 17958 5199 18014 5208
rect 17592 5160 17644 5166
rect 17592 5102 17644 5108
rect 17972 4826 18000 5199
rect 18050 4856 18106 4865
rect 17960 4820 18012 4826
rect 18050 4791 18106 4800
rect 17960 4762 18012 4768
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17512 3738 17540 4422
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17604 3738 17632 3878
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17420 2582 17448 2994
rect 17880 2650 17908 4626
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17972 3194 18000 4558
rect 18064 4214 18092 4791
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 18050 3904 18106 3913
rect 18050 3839 18106 3848
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18064 2990 18092 3839
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 18156 2922 18184 6310
rect 18616 5817 18644 8298
rect 18694 7712 18750 7721
rect 18694 7647 18750 7656
rect 18708 7546 18736 7647
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18800 6118 18828 8599
rect 18892 6866 18920 8774
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18602 5808 18658 5817
rect 18602 5743 18658 5752
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18694 4448 18750 4457
rect 18282 4380 18578 4400
rect 18694 4383 18750 4392
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18616 3058 18644 3334
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 17972 2310 18000 2450
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 17316 1896 17368 1902
rect 17316 1838 17368 1844
rect 17328 1601 17356 1838
rect 18708 1766 18736 4383
rect 18800 2990 18828 5850
rect 19076 4978 19104 8910
rect 19168 7002 19196 13382
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19352 11762 19380 13330
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19444 10810 19472 13262
rect 19706 12336 19762 12345
rect 19706 12271 19708 12280
rect 19760 12271 19762 12280
rect 19708 12242 19760 12248
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19536 11762 19564 12038
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19812 11354 19840 13262
rect 20548 12850 20576 15982
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20640 14249 20668 15846
rect 20626 14240 20682 14249
rect 20626 14175 20682 14184
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19812 10538 19840 11290
rect 19800 10532 19852 10538
rect 19800 10474 19852 10480
rect 19246 10432 19302 10441
rect 19246 10367 19302 10376
rect 19260 9178 19288 10367
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 19260 5166 19288 8978
rect 19444 8634 19472 9454
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19352 7750 19380 8298
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19352 6798 19380 7686
rect 19444 7410 19472 8570
rect 20180 7546 20208 11494
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19352 5778 19380 6054
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19352 5234 19380 5714
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19248 5160 19300 5166
rect 19444 5114 19472 5510
rect 19248 5102 19300 5108
rect 19156 5092 19208 5098
rect 19156 5034 19208 5040
rect 18892 4950 19104 4978
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18696 1760 18748 1766
rect 18696 1702 18748 1708
rect 18328 1692 18380 1698
rect 18328 1634 18380 1640
rect 17314 1592 17370 1601
rect 17314 1527 17370 1536
rect 17776 1148 17828 1154
rect 17776 1090 17828 1096
rect 17236 1006 17356 1034
rect 17328 480 17356 1006
rect 17788 480 17816 1090
rect 18340 480 18368 1634
rect 18800 649 18828 2926
rect 18786 640 18842 649
rect 18786 575 18842 584
rect 18892 480 18920 4950
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 18984 2514 19012 4558
rect 18972 2508 19024 2514
rect 18972 2450 19024 2456
rect 19076 2394 19104 4626
rect 18984 2366 19104 2394
rect 18984 1834 19012 2366
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 19076 1970 19104 2246
rect 19168 2009 19196 5034
rect 19260 3097 19288 5102
rect 19352 5086 19472 5114
rect 19352 4282 19380 5086
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19352 4010 19380 4218
rect 19340 4004 19392 4010
rect 19340 3946 19392 3952
rect 19444 3602 19472 4966
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19430 3496 19486 3505
rect 19430 3431 19486 3440
rect 19444 3126 19472 3431
rect 19628 3194 19656 6666
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19720 3466 19748 6054
rect 19892 5296 19944 5302
rect 19892 5238 19944 5244
rect 19800 5228 19852 5234
rect 19800 5170 19852 5176
rect 19812 4622 19840 5170
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19708 3460 19760 3466
rect 19708 3402 19760 3408
rect 19616 3188 19668 3194
rect 19616 3130 19668 3136
rect 19432 3120 19484 3126
rect 19246 3088 19302 3097
rect 19432 3062 19484 3068
rect 19708 3120 19760 3126
rect 19708 3062 19760 3068
rect 19246 3023 19302 3032
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 19154 2000 19210 2009
rect 19064 1964 19116 1970
rect 19154 1935 19210 1944
rect 19064 1906 19116 1912
rect 18972 1828 19024 1834
rect 18972 1770 19024 1776
rect 18984 1057 19012 1770
rect 18970 1048 19026 1057
rect 18970 983 19026 992
rect 202 0 258 480
rect 662 0 718 480
rect 1214 0 1270 480
rect 1766 0 1822 480
rect 2318 0 2374 480
rect 2870 0 2926 480
rect 3330 0 3386 480
rect 3882 0 3938 480
rect 4434 0 4490 480
rect 4986 0 5042 480
rect 5538 0 5594 480
rect 5998 0 6054 480
rect 6550 0 6606 480
rect 7102 0 7158 480
rect 7654 0 7710 480
rect 8206 0 8262 480
rect 8758 0 8814 480
rect 9218 0 9274 480
rect 9770 0 9826 480
rect 10322 0 10378 480
rect 10874 0 10930 480
rect 11426 0 11482 480
rect 11886 0 11942 480
rect 12438 0 12494 480
rect 12990 0 13046 480
rect 13542 0 13598 480
rect 14094 0 14150 480
rect 14554 0 14610 480
rect 15106 0 15162 480
rect 15658 0 15714 480
rect 16210 0 16266 480
rect 16762 0 16818 480
rect 17314 0 17370 480
rect 17774 0 17830 480
rect 18326 0 18382 480
rect 18878 0 18934 480
rect 19260 241 19288 2450
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19536 2038 19564 2382
rect 19524 2032 19576 2038
rect 19524 1974 19576 1980
rect 19720 610 19748 3062
rect 19904 2922 19932 5238
rect 20088 5234 20116 6870
rect 20180 5234 20208 7482
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19996 3942 20024 4966
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19432 604 19484 610
rect 19432 546 19484 552
rect 19708 604 19760 610
rect 19708 546 19760 552
rect 19444 480 19472 546
rect 19996 480 20024 3674
rect 20088 3058 20116 4422
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 20180 3058 20208 4218
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 20180 2446 20208 2994
rect 20272 2990 20300 12718
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20640 10810 20668 12174
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 3602 20392 10406
rect 20442 10024 20498 10033
rect 20442 9959 20498 9968
rect 20456 6254 20484 9959
rect 20640 9518 20668 10746
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20536 8288 20588 8294
rect 20536 8230 20588 8236
rect 20548 7954 20576 8230
rect 20536 7948 20588 7954
rect 20536 7890 20588 7896
rect 20548 7342 20576 7890
rect 20732 7546 20760 18278
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20824 10198 20852 11698
rect 20812 10192 20864 10198
rect 20812 10134 20864 10140
rect 20824 9722 20852 10134
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 22100 7540 22152 7546
rect 22100 7482 22152 7488
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 21548 3596 21600 3602
rect 21548 3538 21600 3544
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 20994 2952 21050 2961
rect 20994 2887 21050 2896
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 20444 2100 20496 2106
rect 20444 2042 20496 2048
rect 20456 480 20484 2042
rect 21008 480 21036 2887
rect 21560 480 21588 3538
rect 22112 480 22140 7482
rect 22650 3224 22706 3233
rect 22650 3159 22706 3168
rect 22664 480 22692 3159
rect 19246 232 19302 241
rect 19246 167 19302 176
rect 19430 0 19486 480
rect 19982 0 20038 480
rect 20442 0 20498 480
rect 20994 0 21050 480
rect 21546 0 21602 480
rect 22098 0 22154 480
rect 22650 0 22706 480
<< via2 >>
rect 18050 22616 18106 22672
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 662 12144 718 12200
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4066 11464 4122 11520
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4986 3460 5042 3496
rect 4986 3440 4988 3460
rect 4988 3440 5040 3460
rect 5040 3440 5042 3460
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 6458 3984 6514 4040
rect 5814 2896 5870 2952
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 6734 3576 6790 3632
rect 7010 3188 7066 3224
rect 7010 3168 7012 3188
rect 7012 3168 7064 3188
rect 7064 3168 7066 3188
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 9586 12144 9642 12200
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 9862 6740 9864 6760
rect 9864 6740 9916 6760
rect 9916 6740 9918 6760
rect 9862 6704 9918 6740
rect 10230 10104 10286 10160
rect 17774 21664 17830 21720
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 10782 7928 10838 7984
rect 8850 3168 8906 3224
rect 10598 6160 10654 6216
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11794 10376 11850 10432
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11886 3984 11942 4040
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 13266 10140 13268 10160
rect 13268 10140 13320 10160
rect 13320 10140 13322 10160
rect 13266 10104 13322 10140
rect 12254 3032 12310 3088
rect 12530 3032 12586 3088
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14002 10376 14058 10432
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14462 9016 14518 9072
rect 13634 3168 13690 3224
rect 14094 4020 14096 4040
rect 14096 4020 14148 4040
rect 14148 4020 14150 4040
rect 14094 3984 14150 4020
rect 14462 3032 14518 3088
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 17958 18808 18014 18864
rect 18970 22208 19026 22264
rect 18786 20712 18842 20768
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 19062 21256 19118 21312
rect 19614 19352 19670 19408
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18970 17992 19026 18048
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18602 17040 18658 17096
rect 18602 16496 18658 16552
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18786 16088 18842 16144
rect 17866 13232 17922 13288
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 15658 6704 15714 6760
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 16578 3168 16634 3224
rect 17498 9424 17554 9480
rect 17038 2508 17094 2544
rect 17038 2488 17040 2508
rect 17040 2488 17092 2508
rect 17092 2488 17094 2508
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 19062 15156 19118 15192
rect 19062 15136 19064 15156
rect 19064 15136 19116 15156
rect 19116 15136 19118 15156
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18602 13776 18658 13832
rect 20166 20304 20222 20360
rect 19890 19780 19946 19816
rect 19890 19760 19892 19780
rect 19892 19760 19944 19780
rect 19944 19760 19946 19780
rect 20718 18420 20774 18456
rect 20718 18400 20720 18420
rect 20720 18400 20772 18420
rect 20772 18400 20774 18420
rect 19890 17484 19892 17504
rect 19892 17484 19944 17504
rect 19944 17484 19946 17504
rect 19890 17448 19946 17484
rect 19246 15544 19302 15600
rect 19890 14592 19946 14648
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18602 12824 18658 12880
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18786 11872 18842 11928
rect 18694 10920 18750 10976
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18970 11328 19026 11384
rect 18786 8608 18842 8664
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18142 7112 18198 7168
rect 18050 6704 18106 6760
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 17958 5208 18014 5264
rect 18050 4800 18106 4856
rect 18050 3848 18106 3904
rect 18694 7656 18750 7712
rect 18602 5752 18658 5808
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18694 4392 18750 4448
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 19706 12300 19762 12336
rect 19706 12280 19708 12300
rect 19708 12280 19760 12300
rect 19760 12280 19762 12300
rect 20626 14184 20682 14240
rect 19246 10376 19302 10432
rect 17314 1536 17370 1592
rect 18786 584 18842 640
rect 19430 3440 19486 3496
rect 19246 3032 19302 3088
rect 19154 1944 19210 2000
rect 18970 992 19026 1048
rect 20442 9968 20498 10024
rect 20994 2896 21050 2952
rect 22650 3168 22706 3224
rect 19246 176 19302 232
<< metal3 >>
rect 18045 22674 18111 22677
rect 22520 22674 23000 22704
rect 18045 22672 23000 22674
rect 18045 22616 18050 22672
rect 18106 22616 23000 22672
rect 18045 22614 23000 22616
rect 18045 22611 18111 22614
rect 22520 22584 23000 22614
rect 18965 22266 19031 22269
rect 22520 22266 23000 22296
rect 18965 22264 23000 22266
rect 18965 22208 18970 22264
rect 19026 22208 23000 22264
rect 18965 22206 23000 22208
rect 18965 22203 19031 22206
rect 22520 22176 23000 22206
rect 17769 21722 17835 21725
rect 22520 21722 23000 21752
rect 17769 21720 23000 21722
rect 17769 21664 17774 21720
rect 17830 21664 23000 21720
rect 17769 21662 23000 21664
rect 17769 21659 17835 21662
rect 22520 21632 23000 21662
rect 19057 21314 19123 21317
rect 22520 21314 23000 21344
rect 19057 21312 23000 21314
rect 19057 21256 19062 21312
rect 19118 21256 23000 21312
rect 19057 21254 23000 21256
rect 19057 21251 19123 21254
rect 22520 21224 23000 21254
rect 18781 20770 18847 20773
rect 22520 20770 23000 20800
rect 18781 20768 23000 20770
rect 18781 20712 18786 20768
rect 18842 20712 23000 20768
rect 18781 20710 23000 20712
rect 18781 20707 18847 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 22520 20680 23000 20710
rect 18270 20639 18590 20640
rect 20161 20362 20227 20365
rect 22520 20362 23000 20392
rect 20161 20360 23000 20362
rect 20161 20304 20166 20360
rect 20222 20304 23000 20360
rect 20161 20302 23000 20304
rect 20161 20299 20227 20302
rect 22520 20272 23000 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 19885 19818 19951 19821
rect 22520 19818 23000 19848
rect 19885 19816 23000 19818
rect 19885 19760 19890 19816
rect 19946 19760 23000 19816
rect 19885 19758 23000 19760
rect 19885 19755 19951 19758
rect 22520 19728 23000 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 19609 19410 19675 19413
rect 22520 19410 23000 19440
rect 19609 19408 23000 19410
rect 19609 19352 19614 19408
rect 19670 19352 23000 19408
rect 19609 19350 23000 19352
rect 19609 19347 19675 19350
rect 22520 19320 23000 19350
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 17953 18866 18019 18869
rect 22520 18866 23000 18896
rect 17953 18864 23000 18866
rect 17953 18808 17958 18864
rect 18014 18808 23000 18864
rect 17953 18806 23000 18808
rect 17953 18803 18019 18806
rect 22520 18776 23000 18806
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 20713 18458 20779 18461
rect 22520 18458 23000 18488
rect 20713 18456 23000 18458
rect 20713 18400 20718 18456
rect 20774 18400 23000 18456
rect 20713 18398 23000 18400
rect 20713 18395 20779 18398
rect 22520 18368 23000 18398
rect 18965 18050 19031 18053
rect 22520 18050 23000 18080
rect 18965 18048 23000 18050
rect 18965 17992 18970 18048
rect 19026 17992 23000 18048
rect 18965 17990 23000 17992
rect 18965 17987 19031 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22520 17960 23000 17990
rect 14805 17919 15125 17920
rect 19885 17506 19951 17509
rect 22520 17506 23000 17536
rect 19885 17504 23000 17506
rect 19885 17448 19890 17504
rect 19946 17448 23000 17504
rect 19885 17446 23000 17448
rect 19885 17443 19951 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 22520 17416 23000 17446
rect 18270 17375 18590 17376
rect 18597 17098 18663 17101
rect 22520 17098 23000 17128
rect 18597 17096 23000 17098
rect 18597 17040 18602 17096
rect 18658 17040 23000 17096
rect 18597 17038 23000 17040
rect 18597 17035 18663 17038
rect 22520 17008 23000 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 18597 16554 18663 16557
rect 22520 16554 23000 16584
rect 18597 16552 23000 16554
rect 18597 16496 18602 16552
rect 18658 16496 23000 16552
rect 18597 16494 23000 16496
rect 18597 16491 18663 16494
rect 22520 16464 23000 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 18781 16146 18847 16149
rect 22520 16146 23000 16176
rect 18781 16144 23000 16146
rect 18781 16088 18786 16144
rect 18842 16088 23000 16144
rect 18781 16086 23000 16088
rect 18781 16083 18847 16086
rect 22520 16056 23000 16086
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 19241 15602 19307 15605
rect 22520 15602 23000 15632
rect 19241 15600 23000 15602
rect 19241 15544 19246 15600
rect 19302 15544 23000 15600
rect 19241 15542 23000 15544
rect 19241 15539 19307 15542
rect 22520 15512 23000 15542
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 19057 15194 19123 15197
rect 22520 15194 23000 15224
rect 19057 15192 23000 15194
rect 19057 15136 19062 15192
rect 19118 15136 23000 15192
rect 19057 15134 23000 15136
rect 19057 15131 19123 15134
rect 22520 15104 23000 15134
rect 7874 14720 8194 14721
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 19885 14650 19951 14653
rect 22520 14650 23000 14680
rect 19885 14648 23000 14650
rect 19885 14592 19890 14648
rect 19946 14592 23000 14648
rect 19885 14590 23000 14592
rect 19885 14587 19951 14590
rect 22520 14560 23000 14590
rect 20621 14242 20687 14245
rect 22520 14242 23000 14272
rect 20621 14240 23000 14242
rect 20621 14184 20626 14240
rect 20682 14184 23000 14240
rect 20621 14182 23000 14184
rect 20621 14179 20687 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 22520 14152 23000 14182
rect 18270 14111 18590 14112
rect 18597 13834 18663 13837
rect 22520 13834 23000 13864
rect 18597 13832 23000 13834
rect 18597 13776 18602 13832
rect 18658 13776 23000 13832
rect 18597 13774 23000 13776
rect 18597 13771 18663 13774
rect 22520 13744 23000 13774
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 17861 13290 17927 13293
rect 22520 13290 23000 13320
rect 17861 13288 23000 13290
rect 17861 13232 17866 13288
rect 17922 13232 23000 13288
rect 17861 13230 23000 13232
rect 17861 13227 17927 13230
rect 22520 13200 23000 13230
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 18597 12882 18663 12885
rect 22520 12882 23000 12912
rect 18597 12880 23000 12882
rect 18597 12824 18602 12880
rect 18658 12824 23000 12880
rect 18597 12822 23000 12824
rect 18597 12819 18663 12822
rect 22520 12792 23000 12822
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 19701 12338 19767 12341
rect 22520 12338 23000 12368
rect 19701 12336 23000 12338
rect 19701 12280 19706 12336
rect 19762 12280 23000 12336
rect 19701 12278 23000 12280
rect 19701 12275 19767 12278
rect 22520 12248 23000 12278
rect 657 12202 723 12205
rect 9581 12202 9647 12205
rect 657 12200 9647 12202
rect 657 12144 662 12200
rect 718 12144 9586 12200
rect 9642 12144 9647 12200
rect 657 12142 9647 12144
rect 657 12139 723 12142
rect 9581 12139 9647 12142
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 18781 11930 18847 11933
rect 22520 11930 23000 11960
rect 18781 11928 23000 11930
rect 18781 11872 18786 11928
rect 18842 11872 23000 11928
rect 18781 11870 23000 11872
rect 18781 11867 18847 11870
rect 22520 11840 23000 11870
rect 0 11522 480 11552
rect 4061 11522 4127 11525
rect 0 11520 4127 11522
rect 0 11464 4066 11520
rect 4122 11464 4127 11520
rect 0 11462 4127 11464
rect 0 11432 480 11462
rect 4061 11459 4127 11462
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 18965 11386 19031 11389
rect 22520 11386 23000 11416
rect 18965 11384 23000 11386
rect 18965 11328 18970 11384
rect 19026 11328 23000 11384
rect 18965 11326 23000 11328
rect 18965 11323 19031 11326
rect 22520 11296 23000 11326
rect 18689 10978 18755 10981
rect 22520 10978 23000 11008
rect 18689 10976 23000 10978
rect 18689 10920 18694 10976
rect 18750 10920 23000 10976
rect 18689 10918 23000 10920
rect 18689 10915 18755 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 22520 10888 23000 10918
rect 18270 10847 18590 10848
rect 11789 10434 11855 10437
rect 13997 10434 14063 10437
rect 11789 10432 14063 10434
rect 11789 10376 11794 10432
rect 11850 10376 14002 10432
rect 14058 10376 14063 10432
rect 11789 10374 14063 10376
rect 11789 10371 11855 10374
rect 13997 10371 14063 10374
rect 19241 10434 19307 10437
rect 22520 10434 23000 10464
rect 19241 10432 23000 10434
rect 19241 10376 19246 10432
rect 19302 10376 23000 10432
rect 19241 10374 23000 10376
rect 19241 10371 19307 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 22520 10344 23000 10374
rect 14805 10303 15125 10304
rect 10225 10162 10291 10165
rect 13261 10162 13327 10165
rect 10225 10160 13327 10162
rect 10225 10104 10230 10160
rect 10286 10104 13266 10160
rect 13322 10104 13327 10160
rect 10225 10102 13327 10104
rect 10225 10099 10291 10102
rect 13261 10099 13327 10102
rect 20437 10026 20503 10029
rect 22520 10026 23000 10056
rect 20437 10024 23000 10026
rect 20437 9968 20442 10024
rect 20498 9968 23000 10024
rect 20437 9966 23000 9968
rect 20437 9963 20503 9966
rect 22520 9936 23000 9966
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 17493 9482 17559 9485
rect 22520 9482 23000 9512
rect 17493 9480 23000 9482
rect 17493 9424 17498 9480
rect 17554 9424 23000 9480
rect 17493 9422 23000 9424
rect 17493 9419 17559 9422
rect 22520 9392 23000 9422
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 14457 9074 14523 9077
rect 22520 9074 23000 9104
rect 14457 9072 23000 9074
rect 14457 9016 14462 9072
rect 14518 9016 23000 9072
rect 14457 9014 23000 9016
rect 14457 9011 14523 9014
rect 22520 8984 23000 9014
rect 4409 8736 4729 8737
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 18781 8666 18847 8669
rect 22520 8666 23000 8696
rect 18781 8664 23000 8666
rect 18781 8608 18786 8664
rect 18842 8608 23000 8664
rect 18781 8606 23000 8608
rect 18781 8603 18847 8606
rect 22520 8576 23000 8606
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 22520 8122 23000 8152
rect 15334 8062 23000 8122
rect 10777 7986 10843 7989
rect 15334 7986 15394 8062
rect 22520 8032 23000 8062
rect 10777 7984 15394 7986
rect 10777 7928 10782 7984
rect 10838 7928 15394 7984
rect 10777 7926 15394 7928
rect 10777 7923 10843 7926
rect 18689 7714 18755 7717
rect 22520 7714 23000 7744
rect 18689 7712 23000 7714
rect 18689 7656 18694 7712
rect 18750 7656 23000 7712
rect 18689 7654 23000 7656
rect 18689 7651 18755 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 22520 7624 23000 7654
rect 18270 7583 18590 7584
rect 18137 7170 18203 7173
rect 22520 7170 23000 7200
rect 18137 7168 23000 7170
rect 18137 7112 18142 7168
rect 18198 7112 23000 7168
rect 18137 7110 23000 7112
rect 18137 7107 18203 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 22520 7080 23000 7110
rect 14805 7039 15125 7040
rect 9857 6762 9923 6765
rect 15653 6762 15719 6765
rect 9857 6760 15719 6762
rect 9857 6704 9862 6760
rect 9918 6704 15658 6760
rect 15714 6704 15719 6760
rect 9857 6702 15719 6704
rect 9857 6699 9923 6702
rect 15653 6699 15719 6702
rect 18045 6762 18111 6765
rect 22520 6762 23000 6792
rect 18045 6760 23000 6762
rect 18045 6704 18050 6760
rect 18106 6704 23000 6760
rect 18045 6702 23000 6704
rect 18045 6699 18111 6702
rect 22520 6672 23000 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 10593 6218 10659 6221
rect 22520 6218 23000 6248
rect 10593 6216 23000 6218
rect 10593 6160 10598 6216
rect 10654 6160 23000 6216
rect 10593 6158 23000 6160
rect 10593 6155 10659 6158
rect 22520 6128 23000 6158
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 18597 5810 18663 5813
rect 22520 5810 23000 5840
rect 18597 5808 23000 5810
rect 18597 5752 18602 5808
rect 18658 5752 23000 5808
rect 18597 5750 23000 5752
rect 18597 5747 18663 5750
rect 22520 5720 23000 5750
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 17953 5266 18019 5269
rect 22520 5266 23000 5296
rect 17953 5264 23000 5266
rect 17953 5208 17958 5264
rect 18014 5208 23000 5264
rect 17953 5206 23000 5208
rect 17953 5203 18019 5206
rect 22520 5176 23000 5206
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 18045 4858 18111 4861
rect 22520 4858 23000 4888
rect 18045 4856 23000 4858
rect 18045 4800 18050 4856
rect 18106 4800 23000 4856
rect 18045 4798 23000 4800
rect 18045 4795 18111 4798
rect 22520 4768 23000 4798
rect 18689 4450 18755 4453
rect 22520 4450 23000 4480
rect 18689 4448 23000 4450
rect 18689 4392 18694 4448
rect 18750 4392 23000 4448
rect 18689 4390 23000 4392
rect 18689 4387 18755 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 22520 4360 23000 4390
rect 18270 4319 18590 4320
rect 6453 4042 6519 4045
rect 11881 4042 11947 4045
rect 6453 4040 11947 4042
rect 6453 3984 6458 4040
rect 6514 3984 11886 4040
rect 11942 3984 11947 4040
rect 6453 3982 11947 3984
rect 6453 3979 6519 3982
rect 11881 3979 11947 3982
rect 14089 4042 14155 4045
rect 14089 4040 15394 4042
rect 14089 3984 14094 4040
rect 14150 3984 15394 4040
rect 14089 3982 15394 3984
rect 14089 3979 14155 3982
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 3775 15125 3776
rect 15334 3770 15394 3982
rect 18045 3906 18111 3909
rect 22520 3906 23000 3936
rect 18045 3904 23000 3906
rect 18045 3848 18050 3904
rect 18106 3848 23000 3904
rect 18045 3846 23000 3848
rect 18045 3843 18111 3846
rect 22520 3816 23000 3846
rect 15334 3710 19626 3770
rect 6729 3634 6795 3637
rect 6729 3632 19442 3634
rect 6729 3576 6734 3632
rect 6790 3576 19442 3632
rect 6729 3574 19442 3576
rect 6729 3571 6795 3574
rect 19382 3501 19442 3574
rect 4981 3498 5047 3501
rect 4981 3496 18890 3498
rect 4981 3440 4986 3496
rect 5042 3440 18890 3496
rect 4981 3438 18890 3440
rect 19382 3496 19491 3501
rect 19382 3440 19430 3496
rect 19486 3440 19491 3496
rect 19382 3438 19491 3440
rect 19566 3498 19626 3710
rect 22520 3498 23000 3528
rect 19566 3438 23000 3498
rect 4981 3435 5047 3438
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 7005 3226 7071 3229
rect 8845 3226 8911 3229
rect 7005 3224 8911 3226
rect 7005 3168 7010 3224
rect 7066 3168 8850 3224
rect 8906 3168 8911 3224
rect 7005 3166 8911 3168
rect 7005 3163 7071 3166
rect 8845 3163 8911 3166
rect 13629 3226 13695 3229
rect 16573 3226 16639 3229
rect 13629 3224 16639 3226
rect 13629 3168 13634 3224
rect 13690 3168 16578 3224
rect 16634 3168 16639 3224
rect 13629 3166 16639 3168
rect 18830 3226 18890 3438
rect 19425 3435 19491 3438
rect 22520 3408 23000 3438
rect 22645 3226 22711 3229
rect 18830 3224 22711 3226
rect 18830 3168 22650 3224
rect 22706 3168 22711 3224
rect 18830 3166 22711 3168
rect 13629 3163 13695 3166
rect 16573 3163 16639 3166
rect 22645 3163 22711 3166
rect 12249 3090 12315 3093
rect 12525 3090 12591 3093
rect 12249 3088 12591 3090
rect 12249 3032 12254 3088
rect 12310 3032 12530 3088
rect 12586 3032 12591 3088
rect 12249 3030 12591 3032
rect 12249 3027 12315 3030
rect 12525 3027 12591 3030
rect 14457 3090 14523 3093
rect 19241 3090 19307 3093
rect 14457 3088 21282 3090
rect 14457 3032 14462 3088
rect 14518 3032 19246 3088
rect 19302 3032 21282 3088
rect 14457 3030 21282 3032
rect 14457 3027 14523 3030
rect 19241 3027 19307 3030
rect 5809 2954 5875 2957
rect 20989 2954 21055 2957
rect 5809 2952 21055 2954
rect 5809 2896 5814 2952
rect 5870 2896 20994 2952
rect 21050 2896 21055 2952
rect 5809 2894 21055 2896
rect 21222 2954 21282 3030
rect 22520 2954 23000 2984
rect 21222 2894 23000 2954
rect 5809 2891 5875 2894
rect 20989 2891 21055 2894
rect 22520 2864 23000 2894
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 17033 2546 17099 2549
rect 22520 2546 23000 2576
rect 17033 2544 23000 2546
rect 17033 2488 17038 2544
rect 17094 2488 23000 2544
rect 17033 2486 23000 2488
rect 17033 2483 17099 2486
rect 22520 2456 23000 2486
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 19149 2002 19215 2005
rect 22520 2002 23000 2032
rect 19149 2000 23000 2002
rect 19149 1944 19154 2000
rect 19210 1944 23000 2000
rect 19149 1942 23000 1944
rect 19149 1939 19215 1942
rect 22520 1912 23000 1942
rect 17309 1594 17375 1597
rect 22520 1594 23000 1624
rect 17309 1592 23000 1594
rect 17309 1536 17314 1592
rect 17370 1536 23000 1592
rect 17309 1534 23000 1536
rect 17309 1531 17375 1534
rect 22520 1504 23000 1534
rect 18965 1050 19031 1053
rect 22520 1050 23000 1080
rect 18965 1048 23000 1050
rect 18965 992 18970 1048
rect 19026 992 23000 1048
rect 18965 990 23000 992
rect 18965 987 19031 990
rect 22520 960 23000 990
rect 18781 642 18847 645
rect 22520 642 23000 672
rect 18781 640 23000 642
rect 18781 584 18786 640
rect 18842 584 23000 640
rect 18781 582 23000 584
rect 18781 579 18847 582
rect 22520 552 23000 582
rect 19241 234 19307 237
rect 22520 234 23000 264
rect 19241 232 23000 234
rect 19241 176 19246 232
rect 19302 176 23000 232
rect 19241 174 23000 176
rect 19241 171 19307 174
rect 22520 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18590 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 19616 18590 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 18528 18590 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 17440 18590 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 16352 18590 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 15264 18590 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 14176 18590 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 13088 18590 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 12000 18590 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 10912 18590 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 9824 18590 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 8736 18590 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 7648 18590 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 6560 18590 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 5472 18590 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 4384 18590 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 3296 18590 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 2208 18590 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2128 18590 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _33_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4600 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_35
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_41
timestamp 1604681595
transform 1 0 4876 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _72_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5612 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54
timestamp 1604681595
transform 1 0 6072 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 6992 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68
timestamp 1604681595
transform 1 0 7360 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_66
timestamp 1604681595
transform 1 0 7176 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9844 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp 1604681595
transform 1 0 10672 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_90
timestamp 1604681595
transform 1 0 9384 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_102
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _90_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12512 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13064 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 14076 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129
timestamp 1604681595
transform 1 0 12972 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_139
timestamp 1604681595
transform 1 0 13892 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_133
timestamp 1604681595
transform 1 0 13340 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15640 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_160
timestamp 1604681595
transform 1 0 15824 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_150
timestamp 1604681595
transform 1 0 14904 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_178
timestamp 1604681595
transform 1 0 17480 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_167
timestamp 1604681595
transform 1 0 16468 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1604681595
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19044 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_0_204
timestamp 1604681595
transform 1 0 19872 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_193
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1604681595
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1604681595
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_210
timestamp 1604681595
transform 1 0 20424 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_222
timestamp 1604681595
transform 1 0 21528 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1604681595
transform 1 0 4784 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1604681595
transform 1 0 5796 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_43
timestamp 1604681595
transform 1 0 5060 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_55
timestamp 1604681595
transform 1 0 6164 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 6900 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_67
timestamp 1604681595
transform 1 0 7268 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10580 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_119
timestamp 1604681595
transform 1 0 12052 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12788 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_2_143
timestamp 1604681595
transform 1 0 14260 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15640 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 17204 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_2_167
timestamp 1604681595
transform 1 0 16468 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 19412 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_191
timestamp 1604681595
transform 1 0 18676 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_205
timestamp 1604681595
transform 1 0 19964 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1604681595
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1604681595
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_47
timestamp 1604681595
transform 1 0 5428 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_78
timestamp 1604681595
transform 1 0 8280 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9844 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_90
timestamp 1604681595
transform 1 0 9384 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_94
timestamp 1604681595
transform 1 0 9752 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_111
timestamp 1604681595
transform 1 0 11316 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1604681595
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_127
timestamp 1604681595
transform 1 0 12788 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_144
timestamp 1604681595
transform 1 0 14352 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15088 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_168
timestamp 1604681595
transform 1 0 16560 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_180
timestamp 1604681595
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_187
timestamp 1604681595
transform 1 0 18308 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_211
timestamp 1604681595
transform 1 0 20516 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 6532 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7636 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_63
timestamp 1604681595
transform 1 0 6900 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_102
timestamp 1604681595
transform 1 0 10488 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11316 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_110
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_120
timestamp 1604681595
transform 1 0 12144 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12880 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_4_144
timestamp 1604681595
transform 1 0 14352 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1604681595
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_170
timestamp 1604681595
transform 1 0 16744 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_187
timestamp 1604681595
transform 1 0 18308 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_195
timestamp 1604681595
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1604681595
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_47
timestamp 1604681595
transform 1 0 5428 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_53
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_78
timestamp 1604681595
transform 1 0 8280 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9200 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_104
timestamp 1604681595
transform 1 0 10672 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_116
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1604681595
transform 1 0 14168 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_132
timestamp 1604681595
transform 1 0 13248 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_140
timestamp 1604681595
transform 1 0 13984 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_146
timestamp 1604681595
transform 1 0 14536 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_163
timestamp 1604681595
transform 1 0 16100 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_193
timestamp 1604681595
transform 1 0 18860 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_210
timestamp 1604681595
transform 1 0 20424 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1604681595
transform 1 0 21528 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 6164 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_47
timestamp 1604681595
transform 1 0 5428 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_58
timestamp 1604681595
transform 1 0 6440 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_47
timestamp 1604681595
transform 1 0 5428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_53
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_75
timestamp 1604681595
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_78
timestamp 1604681595
transform 1 0 8280 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1604681595
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1604681595
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_97
timestamp 1604681595
transform 1 0 10028 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_102
timestamp 1604681595
transform 1 0 10488 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1604681595
transform 1 0 12236 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_6_133
timestamp 1604681595
transform 1 0 13340 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_145
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_139
timestamp 1604681595
transform 1 0 13892 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_163
timestamp 1604681595
transform 1 0 16100 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_151
timestamp 1604681595
transform 1 0 14996 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18124 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16836 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_177
timestamp 1604681595
transform 1 0 17388 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1604681595
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_200
timestamp 1604681595
transform 1 0 19504 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1604681595
transform 1 0 20516 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1604681595
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1604681595
transform 1 0 20884 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_64
timestamp 1604681595
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_76
timestamp 1604681595
transform 1 0 8096 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12052 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 11776 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_114
timestamp 1604681595
transform 1 0 11592 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_128
timestamp 1604681595
transform 1 0 12880 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_163
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16836 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_180
timestamp 1604681595
transform 1 0 17664 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18400 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1604681595
transform 1 0 19228 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1604681595
transform 1 0 20332 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7084 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9384 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_99
timestamp 1604681595
transform 1 0 10212 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_107
timestamp 1604681595
transform 1 0 10948 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13984 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_9_132
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_156
timestamp 1604681595
transform 1 0 15456 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_164
timestamp 1604681595
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_175
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19412 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_9_190
timestamp 1604681595
transform 1 0 18584 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_198
timestamp 1604681595
transform 1 0 19320 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_215
timestamp 1604681595
transform 1 0 20884 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 5612 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6624 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_44
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_48
timestamp 1604681595
transform 1 0 5520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_52
timestamp 1604681595
transform 1 0 5888 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_76
timestamp 1604681595
transform 1 0 8096 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_109
timestamp 1604681595
transform 1 0 11132 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_133
timestamp 1604681595
transform 1 0 13340 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16284 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_157
timestamp 1604681595
transform 1 0 15548 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17848 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_174
timestamp 1604681595
transform 1 0 17112 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_198
timestamp 1604681595
transform 1 0 19320 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_210
timestamp 1604681595
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6992 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1604681595
transform 1 0 8464 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9844 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_92
timestamp 1604681595
transform 1 0 9568 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_111
timestamp 1604681595
transform 1 0 11316 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 1604681595
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_127
timestamp 1604681595
transform 1 0 12788 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16100 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_151
timestamp 1604681595
transform 1 0 14996 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_162
timestamp 1604681595
transform 1 0 16008 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_172
timestamp 1604681595
transform 1 0 16928 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_180
timestamp 1604681595
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_188
timestamp 1604681595
transform 1 0 18400 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_212
timestamp 1604681595
transform 1 0 20608 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1604681595
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_67
timestamp 1604681595
transform 1 0 7268 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_103
timestamp 1604681595
transform 1 0 10580 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11316 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_120
timestamp 1604681595
transform 1 0 12144 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_132
timestamp 1604681595
transform 1 0 13248 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_160
timestamp 1604681595
transform 1 0 15824 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16560 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_184
timestamp 1604681595
transform 1 0 18032 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18768 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1604681595
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1604681595
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1604681595
transform 1 0 6992 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7544 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_67
timestamp 1604681595
transform 1 0 7268 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 9844 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_94
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_102
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11224 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12696 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_126
timestamp 1604681595
transform 1 0 12696 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_134
timestamp 1604681595
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_135
timestamp 1604681595
transform 1 0 13524 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16284 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_151
timestamp 1604681595
transform 1 0 14996 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_157
timestamp 1604681595
transform 1 0 15548 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _89_
timestamp 1604681595
transform 1 0 18308 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_175
timestamp 1604681595
transform 1 0 17204 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_181
timestamp 1604681595
transform 1 0 17756 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19412 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18492 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_191
timestamp 1604681595
transform 1 0 18676 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_198
timestamp 1604681595
transform 1 0 19320 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1604681595
transform 1 0 20884 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1604681595
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1604681595
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8464 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_96
timestamp 1604681595
transform 1 0 9936 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_104
timestamp 1604681595
transform 1 0 10672 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14076 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_139
timestamp 1604681595
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_157
timestamp 1604681595
transform 1 0 15548 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_165
timestamp 1604681595
transform 1 0 16284 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 18308 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19412 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_191
timestamp 1604681595
transform 1 0 18676 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1604681595
transform 1 0 20884 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_103
timestamp 1604681595
transform 1 0 10580 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 11776 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_115
timestamp 1604681595
transform 1 0 11684 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_119
timestamp 1604681595
transform 1 0 12052 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13064 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_16_127
timestamp 1604681595
transform 1 0 12788 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1604681595
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_157
timestamp 1604681595
transform 1 0 15548 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16744 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 16560 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_179
timestamp 1604681595
transform 1 0 17572 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_187
timestamp 1604681595
transform 1 0 18308 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18400 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_204
timestamp 1604681595
transform 1 0 19872 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1604681595
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1604681595
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_104
timestamp 1604681595
transform 1 0 10672 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_116
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13064 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1604681595
transform 1 0 12972 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_139
timestamp 1604681595
transform 1 0 13892 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14628 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_156
timestamp 1604681595
transform 1 0 15456 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_173
timestamp 1604681595
transform 1 0 17020 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_187
timestamp 1604681595
transform 1 0 18308 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19044 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_204
timestamp 1604681595
transform 1 0 19872 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 20608 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_215
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9844 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_84
timestamp 1604681595
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_104
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11408 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_121
timestamp 1604681595
transform 1 0 12236 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12972 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 15640 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_162
timestamp 1604681595
transform 1 0 16008 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16744 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_186
timestamp 1604681595
transform 1 0 18216 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_194
timestamp 1604681595
transform 1 0 18952 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_206
timestamp 1604681595
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11316 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_105
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 14168 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12788 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_19_143
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_127
timestamp 1604681595
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_139
timestamp 1604681595
transform 1 0 13892 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 15456 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_155
timestamp 1604681595
transform 1 0 15364 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17572 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_170
timestamp 1604681595
transform 1 0 16744 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_178
timestamp 1604681595
transform 1 0 17480 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_200
timestamp 1604681595
transform 1 0 19504 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_188
timestamp 1604681595
transform 1 0 18400 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_196
timestamp 1604681595
transform 1 0 19136 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_206
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 1604681595
transform 1 0 20792 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_222
timestamp 1604681595
transform 1 0 21528 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1604681595
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_144
timestamp 1604681595
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1604681595
transform 1 0 14536 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15548 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1604681595
transform 1 0 14812 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_166
timestamp 1604681595
transform 1 0 16376 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1604681595
transform 1 0 17480 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1604681595
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18492 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19780 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_188
timestamp 1604681595
transform 1 0 18400 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_195
timestamp 1604681595
transform 1 0 19044 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_209
timestamp 1604681595
transform 1 0 20332 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1604681595
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_74
timestamp 1604681595
transform 1 0 7912 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_81
timestamp 1604681595
transform 1 0 8556 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1604681595
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1604681595
transform 1 0 12512 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_117
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_123
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_127
timestamp 1604681595
transform 1 0 12788 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_139
timestamp 1604681595
transform 1 0 13892 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 16284 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_157
timestamp 1604681595
transform 1 0 15548 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 17296 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_168
timestamp 1604681595
transform 1 0 16560 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_180
timestamp 1604681595
transform 1 0 17664 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 18400 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_192
timestamp 1604681595
transform 1 0 18768 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7728 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_70
timestamp 1604681595
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_78
timestamp 1604681595
transform 1 0 8280 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_92
timestamp 1604681595
transform 1 0 9568 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_104
timestamp 1604681595
transform 1 0 10672 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_116
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604681595
transform 1 0 16928 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_171
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 18860 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19964 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_192
timestamp 1604681595
transform 1 0 18768 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_197
timestamp 1604681595
transform 1 0 19228 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_211
timestamp 1604681595
transform 1 0 20516 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 1604681595
transform 1 0 10396 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_108
timestamp 1604681595
transform 1 0 11040 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_120
timestamp 1604681595
transform 1 0 12144 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_132
timestamp 1604681595
transform 1 0 13248 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_144
timestamp 1604681595
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1604681595
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_194
timestamp 1604681595
transform 1 0 18952 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1604681595
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 18308 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1604681595
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 19412 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_191
timestamp 1604681595
transform 1 0 18676 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_203
timestamp 1604681595
transform 1 0 19780 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 1604681595
transform 1 0 20884 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12512 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_117
timestamp 1604681595
transform 1 0 11868 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_125
timestamp 1604681595
transform 1 0 12604 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12696 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_132
timestamp 1604681595
transform 1 0 13248 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_144
timestamp 1604681595
transform 1 0 14352 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_130
timestamp 1604681595
transform 1 0 13064 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_142
timestamp 1604681595
transform 1 0 14168 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1604681595
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_154
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_166
timestamp 1604681595
transform 1 0 16376 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_186
timestamp 1604681595
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1604681595
transform 1 0 17480 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1604681595
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 18768 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 18400 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19872 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_192
timestamp 1604681595
transform 1 0 18768 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_206
timestamp 1604681595
transform 1 0 20056 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_210
timestamp 1604681595
transform 1 0 20424 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_222
timestamp 1604681595
transform 1 0 21528 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_206
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10396 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_107
timestamp 1604681595
transform 1 0 10948 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1604681595
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 13248 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_131
timestamp 1604681595
transform 1 0 13156 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_136
timestamp 1604681595
transform 1 0 13616 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_148
timestamp 1604681595
transform 1 0 14720 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_160
timestamp 1604681595
transform 1 0 15824 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_172
timestamp 1604681595
transform 1 0 16928 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_180
timestamp 1604681595
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 19412 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_203
timestamp 1604681595
transform 1 0 19780 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_215
timestamp 1604681595
transform 1 0 20884 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10304 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_99
timestamp 1604681595
transform 1 0 10212 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_106
timestamp 1604681595
transform 1 0 10856 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_118
timestamp 1604681595
transform 1 0 11960 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13800 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_130
timestamp 1604681595
transform 1 0 13064 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_144
timestamp 1604681595
transform 1 0 14352 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1604681595
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_190
timestamp 1604681595
transform 1 0 18584 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_198
timestamp 1604681595
transform 1 0 19320 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13984 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_129
timestamp 1604681595
transform 1 0 12972 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_137
timestamp 1604681595
transform 1 0 13708 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_156
timestamp 1604681595
transform 1 0 15456 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_168
timestamp 1604681595
transform 1 0 16560 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1604681595
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 18768 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19872 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_210
timestamp 1604681595
transform 1 0 20424 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1604681595
transform 1 0 21528 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1604681595
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_38
timestamp 1604681595
transform 1 0 4600 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_50
timestamp 1604681595
transform 1 0 5704 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_62
timestamp 1604681595
transform 1 0 6808 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_74
timestamp 1604681595
transform 1 0 7912 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_86
timestamp 1604681595
transform 1 0 9016 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1604681595
transform 1 0 17572 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_178
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_182
timestamp 1604681595
transform 1 0 17848 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_194
timestamp 1604681595
transform 1 0 18952 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1604681595
transform 1 0 5152 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_56
timestamp 1604681595
transform 1 0 6256 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_63
timestamp 1604681595
transform 1 0 6900 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_75
timestamp 1604681595
transform 1 0 8004 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_87
timestamp 1604681595
transform 1 0 9108 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_106
timestamp 1604681595
transform 1 0 10856 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1604681595
transform 1 0 12604 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1604681595
transform 1 0 13708 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1604681595
transform 1 0 14812 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1604681595
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_180
timestamp 1604681595
transform 1 0 17664 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_187
timestamp 1604681595
transform 1 0 18308 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 18860 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 19964 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_197
timestamp 1604681595
transform 1 0 19228 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_209
timestamp 1604681595
transform 1 0 20332 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 130 592
<< labels >>
rlabel metal2 s 22098 0 22154 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 2870 22520 2926 23000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 22650 0 22706 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 20074 22520 20130 23000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_1_
port 4 nsew default input
rlabel metal2 s 14370 22520 14426 23000 6 ccff_head
port 5 nsew default input
rlabel metal3 s 0 11432 480 11552 6 ccff_tail
port 6 nsew default tristate
rlabel metal3 s 22520 3816 23000 3936 6 chanx_right_in[0]
port 7 nsew default input
rlabel metal3 s 22520 8576 23000 8696 6 chanx_right_in[10]
port 8 nsew default input
rlabel metal3 s 22520 8984 23000 9104 6 chanx_right_in[11]
port 9 nsew default input
rlabel metal3 s 22520 9392 23000 9512 6 chanx_right_in[12]
port 10 nsew default input
rlabel metal3 s 22520 9936 23000 10056 6 chanx_right_in[13]
port 11 nsew default input
rlabel metal3 s 22520 10344 23000 10464 6 chanx_right_in[14]
port 12 nsew default input
rlabel metal3 s 22520 10888 23000 11008 6 chanx_right_in[15]
port 13 nsew default input
rlabel metal3 s 22520 11296 23000 11416 6 chanx_right_in[16]
port 14 nsew default input
rlabel metal3 s 22520 11840 23000 11960 6 chanx_right_in[17]
port 15 nsew default input
rlabel metal3 s 22520 12248 23000 12368 6 chanx_right_in[18]
port 16 nsew default input
rlabel metal3 s 22520 12792 23000 12912 6 chanx_right_in[19]
port 17 nsew default input
rlabel metal3 s 22520 4360 23000 4480 6 chanx_right_in[1]
port 18 nsew default input
rlabel metal3 s 22520 4768 23000 4888 6 chanx_right_in[2]
port 19 nsew default input
rlabel metal3 s 22520 5176 23000 5296 6 chanx_right_in[3]
port 20 nsew default input
rlabel metal3 s 22520 5720 23000 5840 6 chanx_right_in[4]
port 21 nsew default input
rlabel metal3 s 22520 6128 23000 6248 6 chanx_right_in[5]
port 22 nsew default input
rlabel metal3 s 22520 6672 23000 6792 6 chanx_right_in[6]
port 23 nsew default input
rlabel metal3 s 22520 7080 23000 7200 6 chanx_right_in[7]
port 24 nsew default input
rlabel metal3 s 22520 7624 23000 7744 6 chanx_right_in[8]
port 25 nsew default input
rlabel metal3 s 22520 8032 23000 8152 6 chanx_right_in[9]
port 26 nsew default input
rlabel metal3 s 22520 13200 23000 13320 6 chanx_right_out[0]
port 27 nsew default tristate
rlabel metal3 s 22520 17960 23000 18080 6 chanx_right_out[10]
port 28 nsew default tristate
rlabel metal3 s 22520 18368 23000 18488 6 chanx_right_out[11]
port 29 nsew default tristate
rlabel metal3 s 22520 18776 23000 18896 6 chanx_right_out[12]
port 30 nsew default tristate
rlabel metal3 s 22520 19320 23000 19440 6 chanx_right_out[13]
port 31 nsew default tristate
rlabel metal3 s 22520 19728 23000 19848 6 chanx_right_out[14]
port 32 nsew default tristate
rlabel metal3 s 22520 20272 23000 20392 6 chanx_right_out[15]
port 33 nsew default tristate
rlabel metal3 s 22520 20680 23000 20800 6 chanx_right_out[16]
port 34 nsew default tristate
rlabel metal3 s 22520 21224 23000 21344 6 chanx_right_out[17]
port 35 nsew default tristate
rlabel metal3 s 22520 21632 23000 21752 6 chanx_right_out[18]
port 36 nsew default tristate
rlabel metal3 s 22520 22176 23000 22296 6 chanx_right_out[19]
port 37 nsew default tristate
rlabel metal3 s 22520 13744 23000 13864 6 chanx_right_out[1]
port 38 nsew default tristate
rlabel metal3 s 22520 14152 23000 14272 6 chanx_right_out[2]
port 39 nsew default tristate
rlabel metal3 s 22520 14560 23000 14680 6 chanx_right_out[3]
port 40 nsew default tristate
rlabel metal3 s 22520 15104 23000 15224 6 chanx_right_out[4]
port 41 nsew default tristate
rlabel metal3 s 22520 15512 23000 15632 6 chanx_right_out[5]
port 42 nsew default tristate
rlabel metal3 s 22520 16056 23000 16176 6 chanx_right_out[6]
port 43 nsew default tristate
rlabel metal3 s 22520 16464 23000 16584 6 chanx_right_out[7]
port 44 nsew default tristate
rlabel metal3 s 22520 17008 23000 17128 6 chanx_right_out[8]
port 45 nsew default tristate
rlabel metal3 s 22520 17416 23000 17536 6 chanx_right_out[9]
port 46 nsew default tristate
rlabel metal2 s 662 0 718 480 6 chany_bottom_in[0]
port 47 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_in[10]
port 48 nsew default input
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[11]
port 49 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[12]
port 50 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[13]
port 51 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[14]
port 52 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chany_bottom_in[15]
port 53 nsew default input
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_in[16]
port 54 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[17]
port 55 nsew default input
rlabel metal2 s 10322 0 10378 480 6 chany_bottom_in[18]
port 56 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[19]
port 57 nsew default input
rlabel metal2 s 1214 0 1270 480 6 chany_bottom_in[1]
port 58 nsew default input
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_in[2]
port 59 nsew default input
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_in[3]
port 60 nsew default input
rlabel metal2 s 2870 0 2926 480 6 chany_bottom_in[4]
port 61 nsew default input
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_in[5]
port 62 nsew default input
rlabel metal2 s 3882 0 3938 480 6 chany_bottom_in[6]
port 63 nsew default input
rlabel metal2 s 4434 0 4490 480 6 chany_bottom_in[7]
port 64 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[8]
port 65 nsew default input
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_in[9]
port 66 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chany_bottom_out[0]
port 67 nsew default tristate
rlabel metal2 s 16762 0 16818 480 6 chany_bottom_out[10]
port 68 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_out[11]
port 69 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_out[12]
port 70 nsew default tristate
rlabel metal2 s 18326 0 18382 480 6 chany_bottom_out[13]
port 71 nsew default tristate
rlabel metal2 s 18878 0 18934 480 6 chany_bottom_out[14]
port 72 nsew default tristate
rlabel metal2 s 19430 0 19486 480 6 chany_bottom_out[15]
port 73 nsew default tristate
rlabel metal2 s 19982 0 20038 480 6 chany_bottom_out[16]
port 74 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[17]
port 75 nsew default tristate
rlabel metal2 s 20994 0 21050 480 6 chany_bottom_out[18]
port 76 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[19]
port 77 nsew default tristate
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_out[1]
port 78 nsew default tristate
rlabel metal2 s 12438 0 12494 480 6 chany_bottom_out[2]
port 79 nsew default tristate
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_out[3]
port 80 nsew default tristate
rlabel metal2 s 13542 0 13598 480 6 chany_bottom_out[4]
port 81 nsew default tristate
rlabel metal2 s 14094 0 14150 480 6 chany_bottom_out[5]
port 82 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[6]
port 83 nsew default tristate
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_out[7]
port 84 nsew default tristate
rlabel metal2 s 15658 0 15714 480 6 chany_bottom_out[8]
port 85 nsew default tristate
rlabel metal2 s 16210 0 16266 480 6 chany_bottom_out[9]
port 86 nsew default tristate
rlabel metal2 s 8574 22520 8630 23000 6 prog_clk
port 87 nsew default input
rlabel metal3 s 22520 144 23000 264 6 right_bottom_grid_pin_34_
port 88 nsew default input
rlabel metal3 s 22520 552 23000 672 6 right_bottom_grid_pin_35_
port 89 nsew default input
rlabel metal3 s 22520 960 23000 1080 6 right_bottom_grid_pin_36_
port 90 nsew default input
rlabel metal3 s 22520 1504 23000 1624 6 right_bottom_grid_pin_37_
port 91 nsew default input
rlabel metal3 s 22520 1912 23000 2032 6 right_bottom_grid_pin_38_
port 92 nsew default input
rlabel metal3 s 22520 2456 23000 2576 6 right_bottom_grid_pin_39_
port 93 nsew default input
rlabel metal3 s 22520 2864 23000 2984 6 right_bottom_grid_pin_40_
port 94 nsew default input
rlabel metal3 s 22520 3408 23000 3528 6 right_bottom_grid_pin_41_
port 95 nsew default input
rlabel metal3 s 22520 22584 23000 22704 6 right_top_grid_pin_1_
port 96 nsew default input
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 97 nsew default input
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 98 nsew default input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
