magic
tech EFS8A
magscale 1 2
timestamp 1602042383
<< locali >>
rect 5675 14433 5710 14467
rect 5123 12257 5158 12291
rect 14519 10761 14657 10795
rect 14139 10081 14266 10115
rect 5491 6817 5526 6851
rect 13771 6817 13806 6851
rect 6319 5729 6354 5763
rect 10241 5729 10402 5763
rect 12943 5729 12978 5763
rect 10241 5559 10275 5729
rect 1547 3689 1593 3723
rect 1443 3553 1478 3587
rect 7021 3553 7182 3587
rect 7021 3519 7055 3553
<< viali >>
rect 11437 18377 11471 18411
rect 1476 18173 1510 18207
rect 1869 18173 1903 18207
rect 2488 18173 2522 18207
rect 2881 18173 2915 18207
rect 5156 18173 5190 18207
rect 5549 18173 5583 18207
rect 8100 18173 8134 18207
rect 8493 18173 8527 18207
rect 11044 18173 11078 18207
rect 13896 18173 13930 18207
rect 14289 18173 14323 18207
rect 7021 18105 7055 18139
rect 1547 18037 1581 18071
rect 2559 18037 2593 18071
rect 4077 18037 4111 18071
rect 5227 18037 5261 18071
rect 8171 18037 8205 18071
rect 9965 18037 9999 18071
rect 11115 18037 11149 18071
rect 13967 18037 14001 18071
rect 8125 17833 8159 17867
rect 10241 17833 10275 17867
rect 13369 17833 13403 17867
rect 4905 17765 4939 17799
rect 11529 17765 11563 17799
rect 1409 17697 1443 17731
rect 3040 17697 3074 17731
rect 7941 17697 7975 17731
rect 10057 17697 10091 17731
rect 13185 17697 13219 17731
rect 16440 17697 16474 17731
rect 4261 17629 4295 17663
rect 5825 17629 5859 17663
rect 12173 17629 12207 17663
rect 15393 17629 15427 17663
rect 6377 17561 6411 17595
rect 1593 17493 1627 17527
rect 3111 17493 3145 17527
rect 16543 17493 16577 17527
rect 1593 17289 1627 17323
rect 3249 17289 3283 17323
rect 3985 17289 4019 17323
rect 8217 17289 8251 17323
rect 8585 17289 8619 17323
rect 10333 17289 10367 17323
rect 11529 17289 11563 17323
rect 14473 17289 14507 17323
rect 16221 17289 16255 17323
rect 16497 17289 16531 17323
rect 4169 17153 4203 17187
rect 4813 17153 4847 17187
rect 9137 17153 9171 17187
rect 10609 17153 10643 17187
rect 13461 17153 13495 17187
rect 14749 17153 14783 17187
rect 15117 17153 15151 17187
rect 5784 17085 5818 17119
rect 6193 17085 6227 17119
rect 16313 17085 16347 17119
rect 2053 17017 2087 17051
rect 2237 17017 2271 17051
rect 2881 17017 2915 17051
rect 5871 17017 5905 17051
rect 7021 17017 7055 17051
rect 7297 17017 7331 17051
rect 7941 17017 7975 17051
rect 8861 17017 8895 17051
rect 11253 17017 11287 17051
rect 13185 17017 13219 17051
rect 6653 16949 6687 16983
rect 10057 16949 10091 16983
rect 12909 16949 12943 16983
rect 16865 16949 16899 16983
rect 4353 16745 4387 16779
rect 4721 16745 4755 16779
rect 6193 16745 6227 16779
rect 13185 16745 13219 16779
rect 13691 16745 13725 16779
rect 1777 16677 1811 16711
rect 11621 16677 11655 16711
rect 15761 16677 15795 16711
rect 4537 16609 4571 16643
rect 6009 16609 6043 16643
rect 13620 16609 13654 16643
rect 2237 16541 2271 16575
rect 8125 16541 8159 16575
rect 8493 16541 8527 16575
rect 10057 16541 10091 16575
rect 10333 16541 10367 16575
rect 11897 16541 11931 16575
rect 16313 16473 16347 16507
rect 1685 16201 1719 16235
rect 3893 16201 3927 16235
rect 5089 16201 5123 16235
rect 5641 16201 5675 16235
rect 5871 16201 5905 16235
rect 10885 16201 10919 16235
rect 12679 16201 12713 16235
rect 13645 16201 13679 16235
rect 15117 16201 15151 16235
rect 15485 16201 15519 16235
rect 9229 16133 9263 16167
rect 11621 16133 11655 16167
rect 16313 16133 16347 16167
rect 2145 16065 2179 16099
rect 4169 16065 4203 16099
rect 4445 16065 4479 16099
rect 6285 16065 6319 16099
rect 7205 16065 7239 16099
rect 9505 16065 9539 16099
rect 10149 16065 10183 16099
rect 15761 16065 15795 16099
rect 5800 15997 5834 16031
rect 8125 15997 8159 16031
rect 8468 15997 8502 16031
rect 11044 15997 11078 16031
rect 12576 15997 12610 16031
rect 13001 15997 13035 16031
rect 1869 15929 1903 15963
rect 6653 15929 6687 15963
rect 6929 15929 6963 15963
rect 2789 15861 2823 15895
rect 8539 15861 8573 15895
rect 8953 15861 8987 15895
rect 10425 15861 10459 15895
rect 11115 15861 11149 15895
rect 2421 15589 2455 15623
rect 6101 15589 6135 15623
rect 7849 15589 7883 15623
rect 11161 15589 11195 15623
rect 1777 15453 1811 15487
rect 4077 15453 4111 15487
rect 6561 15453 6595 15487
rect 8125 15453 8159 15487
rect 10517 15453 10551 15487
rect 15853 15453 15887 15487
rect 16129 15453 16163 15487
rect 1777 15113 1811 15147
rect 6193 15113 6227 15147
rect 7849 15113 7883 15147
rect 10425 15113 10459 15147
rect 10747 15113 10781 15147
rect 15853 15113 15887 15147
rect 16267 15113 16301 15147
rect 5733 15045 5767 15079
rect 1961 14977 1995 15011
rect 2881 14977 2915 15011
rect 4261 14977 4295 15011
rect 6837 14977 6871 15011
rect 9597 14977 9631 15011
rect 10676 14909 10710 14943
rect 16196 14909 16230 14943
rect 2605 14841 2639 14875
rect 3433 14841 3467 14875
rect 3617 14841 3651 14875
rect 4997 14841 5031 14875
rect 5181 14841 5215 14875
rect 11069 14773 11103 14807
rect 16589 14773 16623 14807
rect 2605 14569 2639 14603
rect 5779 14569 5813 14603
rect 6791 14569 6825 14603
rect 2237 14501 2271 14535
rect 5641 14433 5675 14467
rect 6720 14433 6754 14467
rect 1593 14365 1627 14399
rect 4169 14365 4203 14399
rect 4721 14297 4755 14331
rect 4077 14025 4111 14059
rect 4307 14025 4341 14059
rect 7113 14025 7147 14059
rect 5641 13957 5675 13991
rect 1869 13889 1903 13923
rect 2697 13889 2731 13923
rect 2973 13889 3007 13923
rect 4721 13889 4755 13923
rect 1444 13821 1478 13855
rect 1547 13821 1581 13855
rect 4236 13821 4270 13855
rect 5216 13821 5250 13855
rect 6009 13821 6043 13855
rect 5319 13753 5353 13787
rect 2237 13685 2271 13719
rect 1593 13481 1627 13515
rect 4215 13481 4249 13515
rect 1409 13345 1443 13379
rect 2580 13345 2614 13379
rect 4112 13345 4146 13379
rect 16104 13345 16138 13379
rect 2053 13141 2087 13175
rect 2651 13141 2685 13175
rect 16175 13141 16209 13175
rect 1547 12937 1581 12971
rect 16129 12937 16163 12971
rect 3065 12869 3099 12903
rect 16497 12869 16531 12903
rect 2329 12801 2363 12835
rect 2513 12801 2547 12835
rect 3985 12801 4019 12835
rect 1476 12733 1510 12767
rect 1869 12733 1903 12767
rect 5089 12733 5123 12767
rect 13680 12733 13714 12767
rect 14105 12733 14139 12767
rect 16313 12733 16347 12767
rect 16865 12733 16899 12767
rect 4445 12597 4479 12631
rect 5273 12597 5307 12631
rect 5733 12597 5767 12631
rect 13783 12597 13817 12631
rect 15301 12597 15335 12631
rect 2605 12393 2639 12427
rect 6239 12393 6273 12427
rect 5227 12325 5261 12359
rect 15393 12325 15427 12359
rect 1961 12257 1995 12291
rect 5089 12257 5123 12291
rect 6168 12257 6202 12291
rect 4077 12189 4111 12223
rect 15761 12189 15795 12223
rect 2145 12121 2179 12155
rect 1593 12053 1627 12087
rect 2513 11849 2547 11883
rect 6193 11849 6227 11883
rect 14197 11849 14231 11883
rect 15117 11849 15151 11883
rect 15485 11849 15519 11883
rect 4445 11781 4479 11815
rect 1501 11713 1535 11747
rect 3709 11713 3743 11747
rect 3893 11713 3927 11747
rect 15761 11713 15795 11747
rect 16221 11713 16255 11747
rect 14013 11645 14047 11679
rect 14565 11645 14599 11679
rect 2145 11577 2179 11611
rect 5089 11509 5123 11543
rect 2329 11237 2363 11271
rect 15761 11237 15795 11271
rect 1685 11101 1719 11135
rect 16221 11101 16255 11135
rect 14657 10761 14691 10795
rect 15301 10693 15335 10727
rect 3893 10625 3927 10659
rect 14933 10625 14967 10659
rect 16129 10625 16163 10659
rect 4788 10557 4822 10591
rect 5181 10557 5215 10591
rect 14448 10557 14482 10591
rect 1685 10489 1719 10523
rect 2329 10489 2363 10523
rect 2973 10489 3007 10523
rect 3249 10489 3283 10523
rect 15853 10489 15887 10523
rect 2605 10421 2639 10455
rect 4859 10421 4893 10455
rect 15577 10421 15611 10455
rect 1409 10217 1443 10251
rect 1961 10217 1995 10251
rect 14335 10217 14369 10251
rect 2456 10081 2490 10115
rect 14105 10081 14139 10115
rect 15393 10013 15427 10047
rect 15945 9945 15979 9979
rect 2329 9877 2363 9911
rect 2559 9877 2593 9911
rect 15393 9673 15427 9707
rect 2421 9605 2455 9639
rect 1501 9537 1535 9571
rect 14473 9537 14507 9571
rect 15945 9537 15979 9571
rect 3040 9469 3074 9503
rect 3433 9469 3467 9503
rect 2145 9401 2179 9435
rect 15577 9401 15611 9435
rect 3111 9333 3145 9367
rect 14289 9333 14323 9367
rect 1593 9129 1627 9163
rect 2053 9129 2087 9163
rect 1409 8993 1443 9027
rect 2513 8925 2547 8959
rect 16037 8925 16071 8959
rect 16313 8925 16347 8959
rect 15577 8857 15611 8891
rect 12633 8585 12667 8619
rect 16037 8585 16071 8619
rect 16451 8585 16485 8619
rect 16865 8585 16899 8619
rect 1869 8449 1903 8483
rect 2053 8449 2087 8483
rect 2697 8449 2731 8483
rect 3592 8381 3626 8415
rect 3985 8381 4019 8415
rect 12449 8381 12483 8415
rect 16380 8381 16414 8415
rect 3663 8245 3697 8279
rect 13093 8245 13127 8279
rect 1777 8041 1811 8075
rect 13231 8041 13265 8075
rect 13128 7905 13162 7939
rect 2237 7837 2271 7871
rect 2697 7837 2731 7871
rect 12081 7837 12115 7871
rect 16037 7837 16071 7871
rect 16313 7837 16347 7871
rect 12173 7497 12207 7531
rect 14289 7497 14323 7531
rect 16037 7497 16071 7531
rect 16451 7497 16485 7531
rect 1777 7361 1811 7395
rect 2421 7361 2455 7395
rect 2789 7361 2823 7395
rect 5549 7361 5583 7395
rect 12541 7361 12575 7395
rect 12909 7361 12943 7395
rect 13461 7361 13495 7395
rect 14105 7293 14139 7327
rect 14657 7293 14691 7327
rect 16380 7293 16414 7327
rect 5089 7225 5123 7259
rect 5273 7225 5307 7259
rect 16865 7157 16899 7191
rect 5595 6953 5629 6987
rect 13875 6953 13909 6987
rect 12909 6885 12943 6919
rect 5457 6817 5491 6851
rect 13737 6817 13771 6851
rect 1869 6749 1903 6783
rect 2329 6749 2363 6783
rect 12265 6749 12299 6783
rect 13737 6341 13771 6375
rect 1547 6273 1581 6307
rect 2237 6273 2271 6307
rect 9321 6273 9355 6307
rect 12817 6273 12851 6307
rect 1460 6205 1494 6239
rect 1869 6137 1903 6171
rect 9045 6137 9079 6171
rect 12265 6137 12299 6171
rect 12541 6137 12575 6171
rect 5549 6069 5583 6103
rect 7941 6069 7975 6103
rect 8769 6069 8803 6103
rect 11897 6069 11931 6103
rect 13047 5865 13081 5899
rect 8769 5797 8803 5831
rect 6285 5729 6319 5763
rect 12909 5729 12943 5763
rect 8125 5661 8159 5695
rect 10471 5661 10505 5695
rect 11437 5661 11471 5695
rect 11897 5661 11931 5695
rect 6423 5525 6457 5559
rect 10241 5525 10275 5559
rect 6285 5321 6319 5355
rect 7021 5321 7055 5355
rect 8217 5321 8251 5355
rect 9597 5321 9631 5355
rect 11437 5321 11471 5355
rect 13001 5321 13035 5355
rect 7849 5253 7883 5287
rect 7297 5185 7331 5219
rect 9413 5117 9447 5151
rect 10568 5117 10602 5151
rect 10057 5049 10091 5083
rect 10655 5049 10689 5083
rect 10333 4981 10367 5015
rect 11069 4981 11103 5015
rect 7757 4709 7791 4743
rect 8401 4709 8435 4743
rect 12516 4641 12550 4675
rect 9689 4573 9723 4607
rect 10701 4573 10735 4607
rect 1593 4437 1627 4471
rect 12587 4437 12621 4471
rect 7665 4233 7699 4267
rect 1501 4097 1535 4131
rect 2145 4097 2179 4131
rect 8493 4097 8527 4131
rect 8677 4097 8711 4131
rect 10517 4097 10551 4131
rect 10701 4097 10735 4131
rect 7481 4029 7515 4063
rect 14908 4029 14942 4063
rect 15301 4029 15335 4063
rect 15920 4029 15954 4063
rect 9321 3961 9355 3995
rect 11345 3961 11379 3995
rect 7389 3893 7423 3927
rect 8033 3893 8067 3927
rect 12449 3893 12483 3927
rect 13001 3893 13035 3927
rect 14979 3893 15013 3927
rect 15991 3893 16025 3927
rect 16405 3893 16439 3927
rect 1593 3689 1627 3723
rect 7251 3689 7285 3723
rect 8263 3621 8297 3655
rect 10425 3621 10459 3655
rect 15393 3621 15427 3655
rect 1409 3553 1443 3587
rect 8176 3553 8210 3587
rect 13804 3553 13838 3587
rect 7021 3485 7055 3519
rect 9781 3485 9815 3519
rect 11345 3485 11379 3519
rect 11621 3485 11655 3519
rect 15761 3485 15795 3519
rect 13875 3349 13909 3383
rect 1593 3145 1627 3179
rect 8033 3145 8067 3179
rect 9045 3145 9079 3179
rect 11345 3145 11379 3179
rect 12265 3145 12299 3179
rect 15393 3145 15427 3179
rect 16681 3145 16715 3179
rect 8677 3077 8711 3111
rect 12633 3009 12667 3043
rect 14197 3009 14231 3043
rect 14841 3009 14875 3043
rect 15761 3009 15795 3043
rect 8192 2941 8226 2975
rect 9188 2941 9222 2975
rect 9275 2873 9309 2907
rect 9965 2873 9999 2907
rect 10241 2873 10275 2907
rect 10885 2873 10919 2907
rect 13277 2873 13311 2907
rect 16405 2873 16439 2907
rect 7205 2805 7239 2839
rect 8263 2805 8297 2839
rect 9689 2805 9723 2839
rect 13829 2805 13863 2839
rect 12357 2601 12391 2635
rect 14197 2601 14231 2635
rect 11437 2533 11471 2567
rect 12817 2533 12851 2567
rect 16313 2533 16347 2567
rect 8585 2465 8619 2499
rect 9137 2465 9171 2499
rect 14432 2465 14466 2499
rect 10609 2397 10643 2431
rect 10793 2397 10827 2431
rect 14519 2397 14553 2431
rect 15301 2397 15335 2431
rect 15669 2397 15703 2431
rect 8769 2329 8803 2363
rect 13369 2329 13403 2363
rect 14933 2329 14967 2363
<< metal1 >>
rect 12526 20544 12532 20596
rect 12584 20584 12590 20596
rect 13354 20584 13360 20596
rect 12584 20556 13360 20584
rect 12584 20544 12590 20556
rect 13354 20544 13360 20556
rect 13412 20544 13418 20596
rect 15286 19660 15292 19712
rect 15344 19700 15350 19712
rect 16390 19700 16396 19712
rect 15344 19672 16396 19700
rect 15344 19660 15350 19672
rect 16390 19660 16396 19672
rect 16448 19660 16454 19712
rect 1104 18522 17756 18544
rect 1104 18470 4135 18522
rect 4187 18470 4199 18522
rect 4251 18470 4263 18522
rect 4315 18470 4327 18522
rect 4379 18470 10441 18522
rect 10493 18470 10505 18522
rect 10557 18470 10569 18522
rect 10621 18470 10633 18522
rect 10685 18470 16748 18522
rect 16800 18470 16812 18522
rect 16864 18470 16876 18522
rect 16928 18470 16940 18522
rect 16992 18470 17756 18522
rect 1104 18448 17756 18470
rect 11422 18408 11428 18420
rect 11383 18380 11428 18408
rect 11422 18368 11428 18380
rect 11480 18368 11486 18420
rect 1464 18207 1522 18213
rect 1464 18173 1476 18207
rect 1510 18204 1522 18207
rect 1857 18207 1915 18213
rect 1857 18204 1869 18207
rect 1510 18176 1869 18204
rect 1510 18173 1522 18176
rect 1464 18167 1522 18173
rect 1857 18173 1869 18176
rect 1903 18204 1915 18207
rect 2130 18204 2136 18216
rect 1903 18176 2136 18204
rect 1903 18173 1915 18176
rect 1857 18167 1915 18173
rect 2130 18164 2136 18176
rect 2188 18164 2194 18216
rect 2476 18207 2534 18213
rect 2476 18173 2488 18207
rect 2522 18204 2534 18207
rect 2682 18204 2688 18216
rect 2522 18176 2688 18204
rect 2522 18173 2534 18176
rect 2476 18167 2534 18173
rect 2682 18164 2688 18176
rect 2740 18204 2746 18216
rect 2869 18207 2927 18213
rect 2869 18204 2881 18207
rect 2740 18176 2881 18204
rect 2740 18164 2746 18176
rect 2869 18173 2881 18176
rect 2915 18173 2927 18207
rect 2869 18167 2927 18173
rect 4890 18164 4896 18216
rect 4948 18204 4954 18216
rect 5144 18207 5202 18213
rect 5144 18204 5156 18207
rect 4948 18176 5156 18204
rect 4948 18164 4954 18176
rect 5144 18173 5156 18176
rect 5190 18204 5202 18207
rect 5537 18207 5595 18213
rect 5537 18204 5549 18207
rect 5190 18176 5549 18204
rect 5190 18173 5202 18176
rect 5144 18167 5202 18173
rect 5537 18173 5549 18176
rect 5583 18173 5595 18207
rect 5537 18167 5595 18173
rect 8088 18207 8146 18213
rect 8088 18173 8100 18207
rect 8134 18204 8146 18207
rect 8478 18204 8484 18216
rect 8134 18176 8484 18204
rect 8134 18173 8146 18176
rect 8088 18167 8146 18173
rect 8478 18164 8484 18176
rect 8536 18164 8542 18216
rect 11032 18207 11090 18213
rect 11032 18173 11044 18207
rect 11078 18204 11090 18207
rect 11422 18204 11428 18216
rect 11078 18176 11428 18204
rect 11078 18173 11090 18176
rect 11032 18167 11090 18173
rect 11422 18164 11428 18176
rect 11480 18164 11486 18216
rect 11606 18164 11612 18216
rect 11664 18204 11670 18216
rect 13884 18207 13942 18213
rect 13884 18204 13896 18207
rect 11664 18176 13896 18204
rect 11664 18164 11670 18176
rect 13884 18173 13896 18176
rect 13930 18204 13942 18207
rect 14277 18207 14335 18213
rect 14277 18204 14289 18207
rect 13930 18176 14289 18204
rect 13930 18173 13942 18176
rect 13884 18167 13942 18173
rect 14277 18173 14289 18176
rect 14323 18173 14335 18207
rect 14277 18167 14335 18173
rect 7009 18139 7067 18145
rect 7009 18105 7021 18139
rect 7055 18136 7067 18139
rect 8570 18136 8576 18148
rect 7055 18108 8576 18136
rect 7055 18105 7067 18108
rect 7009 18099 7067 18105
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 8662 18096 8668 18148
rect 8720 18136 8726 18148
rect 18414 18136 18420 18148
rect 8720 18108 18420 18136
rect 8720 18096 8726 18108
rect 18414 18096 18420 18108
rect 18472 18096 18478 18148
rect 1394 18028 1400 18080
rect 1452 18068 1458 18080
rect 1535 18071 1593 18077
rect 1535 18068 1547 18071
rect 1452 18040 1547 18068
rect 1452 18028 1458 18040
rect 1535 18037 1547 18040
rect 1581 18037 1593 18071
rect 1535 18031 1593 18037
rect 2038 18028 2044 18080
rect 2096 18068 2102 18080
rect 2547 18071 2605 18077
rect 2547 18068 2559 18071
rect 2096 18040 2559 18068
rect 2096 18028 2102 18040
rect 2547 18037 2559 18040
rect 2593 18037 2605 18071
rect 2547 18031 2605 18037
rect 3970 18028 3976 18080
rect 4028 18068 4034 18080
rect 4065 18071 4123 18077
rect 4065 18068 4077 18071
rect 4028 18040 4077 18068
rect 4028 18028 4034 18040
rect 4065 18037 4077 18040
rect 4111 18037 4123 18071
rect 4065 18031 4123 18037
rect 5074 18028 5080 18080
rect 5132 18068 5138 18080
rect 5215 18071 5273 18077
rect 5215 18068 5227 18071
rect 5132 18040 5227 18068
rect 5132 18028 5138 18040
rect 5215 18037 5227 18040
rect 5261 18037 5273 18071
rect 5215 18031 5273 18037
rect 7926 18028 7932 18080
rect 7984 18068 7990 18080
rect 8159 18071 8217 18077
rect 8159 18068 8171 18071
rect 7984 18040 8171 18068
rect 7984 18028 7990 18040
rect 8159 18037 8171 18040
rect 8205 18037 8217 18071
rect 9950 18068 9956 18080
rect 9911 18040 9956 18068
rect 8159 18031 8217 18037
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 11103 18071 11161 18077
rect 11103 18037 11115 18071
rect 11149 18068 11161 18071
rect 11514 18068 11520 18080
rect 11149 18040 11520 18068
rect 11149 18037 11161 18040
rect 11103 18031 11161 18037
rect 11514 18028 11520 18040
rect 11572 18028 11578 18080
rect 13955 18071 14013 18077
rect 13955 18037 13967 18071
rect 14001 18068 14013 18071
rect 14182 18068 14188 18080
rect 14001 18040 14188 18068
rect 14001 18037 14013 18040
rect 13955 18031 14013 18037
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 1104 17978 17756 18000
rect 1104 17926 7288 17978
rect 7340 17926 7352 17978
rect 7404 17926 7416 17978
rect 7468 17926 7480 17978
rect 7532 17926 13595 17978
rect 13647 17926 13659 17978
rect 13711 17926 13723 17978
rect 13775 17926 13787 17978
rect 13839 17926 17756 17978
rect 1104 17904 17756 17926
rect 14 17824 20 17876
rect 72 17864 78 17876
rect 6086 17864 6092 17876
rect 72 17836 6092 17864
rect 72 17824 78 17836
rect 6086 17824 6092 17836
rect 6144 17824 6150 17876
rect 8110 17864 8116 17876
rect 8071 17836 8116 17864
rect 8110 17824 8116 17836
rect 8168 17824 8174 17876
rect 10226 17864 10232 17876
rect 10187 17836 10232 17864
rect 10226 17824 10232 17836
rect 10284 17824 10290 17876
rect 13357 17867 13415 17873
rect 13357 17833 13369 17867
rect 13403 17864 13415 17867
rect 14366 17864 14372 17876
rect 13403 17836 14372 17864
rect 13403 17833 13415 17836
rect 13357 17827 13415 17833
rect 14366 17824 14372 17836
rect 14424 17824 14430 17876
rect 3234 17796 3240 17808
rect 3043 17768 3240 17796
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 3043 17737 3071 17768
rect 3234 17756 3240 17768
rect 3292 17796 3298 17808
rect 4430 17796 4436 17808
rect 3292 17768 4436 17796
rect 3292 17756 3298 17768
rect 4430 17756 4436 17768
rect 4488 17756 4494 17808
rect 4890 17796 4896 17808
rect 4851 17768 4896 17796
rect 4890 17756 4896 17768
rect 4948 17756 4954 17808
rect 11514 17796 11520 17808
rect 11475 17768 11520 17796
rect 11514 17756 11520 17768
rect 11572 17756 11578 17808
rect 3028 17731 3086 17737
rect 3028 17697 3040 17731
rect 3074 17697 3086 17731
rect 7926 17728 7932 17740
rect 7887 17700 7932 17728
rect 3028 17691 3086 17697
rect 7926 17688 7932 17700
rect 7984 17688 7990 17740
rect 10042 17728 10048 17740
rect 10003 17700 10048 17728
rect 10042 17688 10048 17700
rect 10100 17688 10106 17740
rect 12894 17688 12900 17740
rect 12952 17728 12958 17740
rect 13173 17731 13231 17737
rect 13173 17728 13185 17731
rect 12952 17700 13185 17728
rect 12952 17688 12958 17700
rect 13173 17697 13185 17700
rect 13219 17697 13231 17731
rect 13173 17691 13231 17697
rect 16298 17688 16304 17740
rect 16356 17728 16362 17740
rect 16428 17731 16486 17737
rect 16428 17728 16440 17731
rect 16356 17700 16440 17728
rect 16356 17688 16362 17700
rect 16428 17697 16440 17700
rect 16474 17697 16486 17731
rect 16428 17691 16486 17697
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17629 4307 17663
rect 4249 17623 4307 17629
rect 5813 17663 5871 17669
rect 5813 17629 5825 17663
rect 5859 17660 5871 17663
rect 6638 17660 6644 17672
rect 5859 17632 6644 17660
rect 5859 17629 5871 17632
rect 5813 17623 5871 17629
rect 4264 17592 4292 17623
rect 6638 17620 6644 17632
rect 6696 17620 6702 17672
rect 12158 17660 12164 17672
rect 12119 17632 12164 17660
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 15378 17660 15384 17672
rect 15339 17632 15384 17660
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 4430 17592 4436 17604
rect 4264 17564 4436 17592
rect 4430 17552 4436 17564
rect 4488 17592 4494 17604
rect 6365 17595 6423 17601
rect 6365 17592 6377 17595
rect 4488 17564 6377 17592
rect 4488 17552 4494 17564
rect 6365 17561 6377 17564
rect 6411 17561 6423 17595
rect 6365 17555 6423 17561
rect 106 17484 112 17536
rect 164 17524 170 17536
rect 1581 17527 1639 17533
rect 1581 17524 1593 17527
rect 164 17496 1593 17524
rect 164 17484 170 17496
rect 1581 17493 1593 17496
rect 1627 17493 1639 17527
rect 1581 17487 1639 17493
rect 3099 17527 3157 17533
rect 3099 17493 3111 17527
rect 3145 17524 3157 17527
rect 3878 17524 3884 17536
rect 3145 17496 3884 17524
rect 3145 17493 3157 17496
rect 3099 17487 3157 17493
rect 3878 17484 3884 17496
rect 3936 17484 3942 17536
rect 16206 17484 16212 17536
rect 16264 17524 16270 17536
rect 16531 17527 16589 17533
rect 16531 17524 16543 17527
rect 16264 17496 16543 17524
rect 16264 17484 16270 17496
rect 16531 17493 16543 17496
rect 16577 17493 16589 17527
rect 16531 17487 16589 17493
rect 1104 17434 17756 17456
rect 1104 17382 4135 17434
rect 4187 17382 4199 17434
rect 4251 17382 4263 17434
rect 4315 17382 4327 17434
rect 4379 17382 10441 17434
rect 10493 17382 10505 17434
rect 10557 17382 10569 17434
rect 10621 17382 10633 17434
rect 10685 17382 16748 17434
rect 16800 17382 16812 17434
rect 16864 17382 16876 17434
rect 16928 17382 16940 17434
rect 16992 17382 17756 17434
rect 1104 17360 17756 17382
rect 1394 17280 1400 17332
rect 1452 17320 1458 17332
rect 1581 17323 1639 17329
rect 1581 17320 1593 17323
rect 1452 17292 1593 17320
rect 1452 17280 1458 17292
rect 1581 17289 1593 17292
rect 1627 17289 1639 17323
rect 3234 17320 3240 17332
rect 3195 17292 3240 17320
rect 1581 17283 1639 17289
rect 3234 17280 3240 17292
rect 3292 17280 3298 17332
rect 3970 17320 3976 17332
rect 3931 17292 3976 17320
rect 3970 17280 3976 17292
rect 4028 17320 4034 17332
rect 4028 17292 4200 17320
rect 4028 17280 4034 17292
rect 4172 17193 4200 17292
rect 7926 17280 7932 17332
rect 7984 17320 7990 17332
rect 8205 17323 8263 17329
rect 8205 17320 8217 17323
rect 7984 17292 8217 17320
rect 7984 17280 7990 17292
rect 8205 17289 8217 17292
rect 8251 17289 8263 17323
rect 8570 17320 8576 17332
rect 8531 17292 8576 17320
rect 8205 17283 8263 17289
rect 8570 17280 8576 17292
rect 8628 17280 8634 17332
rect 9950 17280 9956 17332
rect 10008 17320 10014 17332
rect 10321 17323 10379 17329
rect 10321 17320 10333 17323
rect 10008 17292 10333 17320
rect 10008 17280 10014 17292
rect 10321 17289 10333 17292
rect 10367 17320 10379 17323
rect 11514 17320 11520 17332
rect 10367 17292 10640 17320
rect 11475 17292 11520 17320
rect 10367 17289 10379 17292
rect 10321 17283 10379 17289
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17153 4215 17187
rect 4157 17147 4215 17153
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17184 4859 17187
rect 4890 17184 4896 17196
rect 4847 17156 4896 17184
rect 4847 17153 4859 17156
rect 4801 17147 4859 17153
rect 4890 17144 4896 17156
rect 4948 17144 4954 17196
rect 8478 17144 8484 17196
rect 8536 17184 8542 17196
rect 10612 17193 10640 17292
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 14182 17280 14188 17332
rect 14240 17320 14246 17332
rect 14461 17323 14519 17329
rect 14461 17320 14473 17323
rect 14240 17292 14473 17320
rect 14240 17280 14246 17292
rect 14461 17289 14473 17292
rect 14507 17289 14519 17323
rect 16206 17320 16212 17332
rect 16167 17292 16212 17320
rect 14461 17283 14519 17289
rect 9125 17187 9183 17193
rect 9125 17184 9137 17187
rect 8536 17156 9137 17184
rect 8536 17144 8542 17156
rect 9125 17153 9137 17156
rect 9171 17153 9183 17187
rect 9125 17147 9183 17153
rect 10597 17187 10655 17193
rect 10597 17153 10609 17187
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 12158 17144 12164 17196
rect 12216 17184 12222 17196
rect 13449 17187 13507 17193
rect 13449 17184 13461 17187
rect 12216 17156 13461 17184
rect 12216 17144 12222 17156
rect 13449 17153 13461 17156
rect 13495 17153 13507 17187
rect 14476 17184 14504 17283
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 16485 17323 16543 17329
rect 16485 17289 16497 17323
rect 16531 17320 16543 17323
rect 17402 17320 17408 17332
rect 16531 17292 17408 17320
rect 16531 17289 16543 17292
rect 16485 17283 16543 17289
rect 17402 17280 17408 17292
rect 17460 17280 17466 17332
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 14476 17156 14749 17184
rect 13449 17147 13507 17153
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 15102 17184 15108 17196
rect 15063 17156 15108 17184
rect 14737 17147 14795 17153
rect 15102 17144 15108 17156
rect 15160 17144 15166 17196
rect 5772 17119 5830 17125
rect 5772 17085 5784 17119
rect 5818 17116 5830 17119
rect 6086 17116 6092 17128
rect 5818 17088 6092 17116
rect 5818 17085 5830 17088
rect 5772 17079 5830 17085
rect 6086 17076 6092 17088
rect 6144 17116 6150 17128
rect 6181 17119 6239 17125
rect 6181 17116 6193 17119
rect 6144 17088 6193 17116
rect 6144 17076 6150 17088
rect 6181 17085 6193 17088
rect 6227 17085 6239 17119
rect 6181 17079 6239 17085
rect 16206 17076 16212 17128
rect 16264 17116 16270 17128
rect 16301 17119 16359 17125
rect 16301 17116 16313 17119
rect 16264 17088 16313 17116
rect 16264 17076 16270 17088
rect 16301 17085 16313 17088
rect 16347 17085 16359 17119
rect 16301 17079 16359 17085
rect 2041 17051 2099 17057
rect 2041 17017 2053 17051
rect 2087 17048 2099 17051
rect 2225 17051 2283 17057
rect 2225 17048 2237 17051
rect 2087 17020 2237 17048
rect 2087 17017 2099 17020
rect 2041 17011 2099 17017
rect 2225 17017 2237 17020
rect 2271 17048 2283 17051
rect 2314 17048 2320 17060
rect 2271 17020 2320 17048
rect 2271 17017 2283 17020
rect 2225 17011 2283 17017
rect 2314 17008 2320 17020
rect 2372 17008 2378 17060
rect 2869 17051 2927 17057
rect 2869 17017 2881 17051
rect 2915 17048 2927 17051
rect 5859 17051 5917 17057
rect 2915 17020 4016 17048
rect 2915 17017 2927 17020
rect 2869 17011 2927 17017
rect 3988 16980 4016 17020
rect 5859 17017 5871 17051
rect 5905 17048 5917 17051
rect 7009 17051 7067 17057
rect 7009 17048 7021 17051
rect 5905 17020 7021 17048
rect 5905 17017 5917 17020
rect 5859 17011 5917 17017
rect 7009 17017 7021 17020
rect 7055 17048 7067 17051
rect 7285 17051 7343 17057
rect 7285 17048 7297 17051
rect 7055 17020 7297 17048
rect 7055 17017 7067 17020
rect 7009 17011 7067 17017
rect 7285 17017 7297 17020
rect 7331 17017 7343 17051
rect 7285 17011 7343 17017
rect 7929 17051 7987 17057
rect 7929 17017 7941 17051
rect 7975 17048 7987 17051
rect 8202 17048 8208 17060
rect 7975 17020 8208 17048
rect 7975 17017 7987 17020
rect 7929 17011 7987 17017
rect 8202 17008 8208 17020
rect 8260 17008 8266 17060
rect 8570 17008 8576 17060
rect 8628 17048 8634 17060
rect 8849 17051 8907 17057
rect 8849 17048 8861 17051
rect 8628 17020 8861 17048
rect 8628 17008 8634 17020
rect 8849 17017 8861 17020
rect 8895 17017 8907 17051
rect 8849 17011 8907 17017
rect 11241 17051 11299 17057
rect 11241 17017 11253 17051
rect 11287 17048 11299 17051
rect 11882 17048 11888 17060
rect 11287 17020 11888 17048
rect 11287 17017 11299 17020
rect 11241 17011 11299 17017
rect 11882 17008 11888 17020
rect 11940 17008 11946 17060
rect 13170 17048 13176 17060
rect 13131 17020 13176 17048
rect 13170 17008 13176 17020
rect 13228 17008 13234 17060
rect 4430 16980 4436 16992
rect 3988 16952 4436 16980
rect 4430 16940 4436 16952
rect 4488 16940 4494 16992
rect 6638 16980 6644 16992
rect 6599 16952 6644 16980
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 10042 16980 10048 16992
rect 9955 16952 10048 16980
rect 10042 16940 10048 16952
rect 10100 16980 10106 16992
rect 10778 16980 10784 16992
rect 10100 16952 10784 16980
rect 10100 16940 10106 16952
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 12894 16980 12900 16992
rect 12855 16952 12900 16980
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 16298 16940 16304 16992
rect 16356 16980 16362 16992
rect 16853 16983 16911 16989
rect 16853 16980 16865 16983
rect 16356 16952 16865 16980
rect 16356 16940 16362 16952
rect 16853 16949 16865 16952
rect 16899 16949 16911 16983
rect 16853 16943 16911 16949
rect 1104 16890 17756 16912
rect 1104 16838 7288 16890
rect 7340 16838 7352 16890
rect 7404 16838 7416 16890
rect 7468 16838 7480 16890
rect 7532 16838 13595 16890
rect 13647 16838 13659 16890
rect 13711 16838 13723 16890
rect 13775 16838 13787 16890
rect 13839 16838 17756 16890
rect 1104 16816 17756 16838
rect 4341 16779 4399 16785
rect 4341 16745 4353 16779
rect 4387 16776 4399 16779
rect 4430 16776 4436 16788
rect 4387 16748 4436 16776
rect 4387 16745 4399 16748
rect 4341 16739 4399 16745
rect 4430 16736 4436 16748
rect 4488 16736 4494 16788
rect 4709 16779 4767 16785
rect 4709 16745 4721 16779
rect 4755 16776 4767 16779
rect 5442 16776 5448 16788
rect 4755 16748 5448 16776
rect 4755 16745 4767 16748
rect 4709 16739 4767 16745
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 6178 16776 6184 16788
rect 6139 16748 6184 16776
rect 6178 16736 6184 16748
rect 6236 16736 6242 16788
rect 12158 16776 12164 16788
rect 11624 16748 12164 16776
rect 11624 16720 11652 16748
rect 12158 16736 12164 16748
rect 12216 16736 12222 16788
rect 13170 16776 13176 16788
rect 13131 16748 13176 16776
rect 13170 16736 13176 16748
rect 13228 16776 13234 16788
rect 13679 16779 13737 16785
rect 13679 16776 13691 16779
rect 13228 16748 13691 16776
rect 13228 16736 13234 16748
rect 13679 16745 13691 16748
rect 13725 16745 13737 16779
rect 18322 16776 18328 16788
rect 13679 16739 13737 16745
rect 13786 16748 18328 16776
rect 1765 16711 1823 16717
rect 1765 16677 1777 16711
rect 1811 16708 1823 16711
rect 2038 16708 2044 16720
rect 1811 16680 2044 16708
rect 1811 16677 1823 16680
rect 1765 16671 1823 16677
rect 2038 16668 2044 16680
rect 2096 16668 2102 16720
rect 11606 16708 11612 16720
rect 11519 16680 11612 16708
rect 11606 16668 11612 16680
rect 11664 16668 11670 16720
rect 4525 16643 4583 16649
rect 4525 16609 4537 16643
rect 4571 16640 4583 16643
rect 5074 16640 5080 16652
rect 4571 16612 5080 16640
rect 4571 16609 4583 16612
rect 4525 16603 4583 16609
rect 5074 16600 5080 16612
rect 5132 16600 5138 16652
rect 5994 16640 6000 16652
rect 5955 16612 6000 16640
rect 5994 16600 6000 16612
rect 6052 16600 6058 16652
rect 13630 16649 13636 16652
rect 13608 16643 13636 16649
rect 13608 16640 13620 16643
rect 13543 16612 13620 16640
rect 13608 16609 13620 16612
rect 13688 16640 13694 16652
rect 13786 16640 13814 16748
rect 18322 16736 18328 16748
rect 18380 16736 18386 16788
rect 15378 16668 15384 16720
rect 15436 16708 15442 16720
rect 15749 16711 15807 16717
rect 15749 16708 15761 16711
rect 15436 16680 15761 16708
rect 15436 16668 15442 16680
rect 15749 16677 15761 16680
rect 15795 16677 15807 16711
rect 15749 16671 15807 16677
rect 13688 16612 13814 16640
rect 13608 16603 13636 16609
rect 13630 16600 13636 16603
rect 13688 16600 13694 16612
rect 2222 16572 2228 16584
rect 2183 16544 2228 16572
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 8113 16575 8171 16581
rect 8113 16541 8125 16575
rect 8159 16572 8171 16575
rect 8202 16572 8208 16584
rect 8159 16544 8208 16572
rect 8159 16541 8171 16544
rect 8113 16535 8171 16541
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 8478 16572 8484 16584
rect 8439 16544 8484 16572
rect 8478 16532 8484 16544
rect 8536 16532 8542 16584
rect 10042 16572 10048 16584
rect 10003 16544 10048 16572
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 10318 16572 10324 16584
rect 10279 16544 10324 16572
rect 10318 16532 10324 16544
rect 10376 16532 10382 16584
rect 11882 16572 11888 16584
rect 11843 16544 11888 16572
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 16298 16504 16304 16516
rect 16259 16476 16304 16504
rect 16298 16464 16304 16476
rect 16356 16464 16362 16516
rect 1104 16346 17756 16368
rect 1104 16294 4135 16346
rect 4187 16294 4199 16346
rect 4251 16294 4263 16346
rect 4315 16294 4327 16346
rect 4379 16294 10441 16346
rect 10493 16294 10505 16346
rect 10557 16294 10569 16346
rect 10621 16294 10633 16346
rect 10685 16294 16748 16346
rect 16800 16294 16812 16346
rect 16864 16294 16876 16346
rect 16928 16294 16940 16346
rect 16992 16294 17756 16346
rect 1104 16272 17756 16294
rect 1673 16235 1731 16241
rect 1673 16201 1685 16235
rect 1719 16232 1731 16235
rect 2038 16232 2044 16244
rect 1719 16204 2044 16232
rect 1719 16201 1731 16204
rect 1673 16195 1731 16201
rect 2038 16192 2044 16204
rect 2096 16192 2102 16244
rect 3878 16232 3884 16244
rect 3839 16204 3884 16232
rect 3878 16192 3884 16204
rect 3936 16232 3942 16244
rect 5074 16232 5080 16244
rect 3936 16204 4200 16232
rect 5035 16204 5080 16232
rect 3936 16192 3942 16204
rect 2130 16096 2136 16108
rect 2091 16068 2136 16096
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 4172 16105 4200 16204
rect 5074 16192 5080 16204
rect 5132 16192 5138 16244
rect 5629 16235 5687 16241
rect 5629 16201 5641 16235
rect 5675 16232 5687 16235
rect 5859 16235 5917 16241
rect 5859 16232 5871 16235
rect 5675 16204 5871 16232
rect 5675 16201 5687 16204
rect 5629 16195 5687 16201
rect 5859 16201 5871 16204
rect 5905 16232 5917 16235
rect 5994 16232 6000 16244
rect 5905 16204 6000 16232
rect 5905 16201 5917 16204
rect 5859 16195 5917 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 10873 16235 10931 16241
rect 10873 16201 10885 16235
rect 10919 16232 10931 16235
rect 11882 16232 11888 16244
rect 10919 16204 11888 16232
rect 10919 16201 10931 16204
rect 10873 16195 10931 16201
rect 9217 16167 9275 16173
rect 9217 16164 9229 16167
rect 4448 16136 9229 16164
rect 4448 16108 4476 16136
rect 9217 16133 9229 16136
rect 9263 16133 9275 16167
rect 9217 16127 9275 16133
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16065 4215 16099
rect 4430 16096 4436 16108
rect 4391 16068 4436 16096
rect 4157 16059 4215 16065
rect 4430 16056 4436 16068
rect 4488 16056 4494 16108
rect 6273 16099 6331 16105
rect 6273 16096 6285 16099
rect 5803 16068 6285 16096
rect 5803 16037 5831 16068
rect 6273 16065 6285 16068
rect 6319 16096 6331 16099
rect 6546 16096 6552 16108
rect 6319 16068 6552 16096
rect 6319 16065 6331 16068
rect 6273 16059 6331 16065
rect 6546 16056 6552 16068
rect 6604 16096 6610 16108
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 6604 16068 7205 16096
rect 6604 16056 6610 16068
rect 7193 16065 7205 16068
rect 7239 16065 7251 16099
rect 9232 16096 9260 16127
rect 9493 16099 9551 16105
rect 9493 16096 9505 16099
rect 9232 16068 9505 16096
rect 7193 16059 7251 16065
rect 9493 16065 9505 16068
rect 9539 16065 9551 16099
rect 9493 16059 9551 16065
rect 10137 16099 10195 16105
rect 10137 16065 10149 16099
rect 10183 16096 10195 16099
rect 10318 16096 10324 16108
rect 10183 16068 10324 16096
rect 10183 16065 10195 16068
rect 10137 16059 10195 16065
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 5788 16031 5846 16037
rect 5788 15997 5800 16031
rect 5834 15997 5846 16031
rect 5788 15991 5846 15997
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 16028 8171 16031
rect 8202 16028 8208 16040
rect 8159 16000 8208 16028
rect 8159 15997 8171 16000
rect 8113 15991 8171 15997
rect 8202 15988 8208 16000
rect 8260 15988 8266 16040
rect 8456 16031 8514 16037
rect 8456 15997 8468 16031
rect 8502 16028 8514 16031
rect 8938 16028 8944 16040
rect 8502 16000 8944 16028
rect 8502 15997 8514 16000
rect 8456 15991 8514 15997
rect 8938 15988 8944 16000
rect 8996 15988 9002 16040
rect 1857 15963 1915 15969
rect 1857 15929 1869 15963
rect 1903 15960 1915 15963
rect 2222 15960 2228 15972
rect 1903 15932 2228 15960
rect 1903 15929 1915 15932
rect 1857 15923 1915 15929
rect 2222 15920 2228 15932
rect 2280 15920 2286 15972
rect 6641 15963 6699 15969
rect 6641 15929 6653 15963
rect 6687 15960 6699 15963
rect 6730 15960 6736 15972
rect 6687 15932 6736 15960
rect 6687 15929 6699 15932
rect 6641 15923 6699 15929
rect 6730 15920 6736 15932
rect 6788 15960 6794 15972
rect 6917 15963 6975 15969
rect 6917 15960 6929 15963
rect 6788 15932 6929 15960
rect 6788 15920 6794 15932
rect 6917 15929 6929 15932
rect 6963 15929 6975 15963
rect 10336 15960 10364 16056
rect 11047 16037 11075 16204
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 12667 16235 12725 16241
rect 12667 16201 12679 16235
rect 12713 16232 12725 16235
rect 12894 16232 12900 16244
rect 12713 16204 12900 16232
rect 12713 16201 12725 16204
rect 12667 16195 12725 16201
rect 12894 16192 12900 16204
rect 12952 16192 12958 16244
rect 13630 16232 13636 16244
rect 13591 16204 13636 16232
rect 13630 16192 13636 16204
rect 13688 16192 13694 16244
rect 15102 16232 15108 16244
rect 15063 16204 15108 16232
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 15378 16192 15384 16244
rect 15436 16232 15442 16244
rect 15473 16235 15531 16241
rect 15473 16232 15485 16235
rect 15436 16204 15485 16232
rect 15436 16192 15442 16204
rect 15473 16201 15485 16204
rect 15519 16201 15531 16235
rect 15473 16195 15531 16201
rect 11606 16164 11612 16176
rect 11567 16136 11612 16164
rect 11606 16124 11612 16136
rect 11664 16124 11670 16176
rect 15120 16096 15148 16192
rect 16298 16164 16304 16176
rect 16259 16136 16304 16164
rect 16298 16124 16304 16136
rect 16356 16124 16362 16176
rect 15749 16099 15807 16105
rect 15749 16096 15761 16099
rect 15120 16068 15761 16096
rect 15749 16065 15761 16068
rect 15795 16096 15807 16099
rect 16114 16096 16120 16108
rect 15795 16068 16120 16096
rect 15795 16065 15807 16068
rect 15749 16059 15807 16065
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 11032 16031 11090 16037
rect 11032 15997 11044 16031
rect 11078 15997 11090 16031
rect 11032 15991 11090 15997
rect 12564 16031 12622 16037
rect 12564 15997 12576 16031
rect 12610 16028 12622 16031
rect 12989 16031 13047 16037
rect 12989 16028 13001 16031
rect 12610 16000 13001 16028
rect 12610 15997 12622 16000
rect 12564 15991 12622 15997
rect 12989 15997 13001 16000
rect 13035 15997 13047 16031
rect 12989 15991 13047 15997
rect 12579 15960 12607 15991
rect 10336 15932 12607 15960
rect 6917 15923 6975 15929
rect 2240 15892 2268 15920
rect 2777 15895 2835 15901
rect 2777 15892 2789 15895
rect 2240 15864 2789 15892
rect 2777 15861 2789 15864
rect 2823 15861 2835 15895
rect 2777 15855 2835 15861
rect 8110 15852 8116 15904
rect 8168 15892 8174 15904
rect 8527 15895 8585 15901
rect 8527 15892 8539 15895
rect 8168 15864 8539 15892
rect 8168 15852 8174 15864
rect 8527 15861 8539 15864
rect 8573 15861 8585 15895
rect 8938 15892 8944 15904
rect 8899 15864 8944 15892
rect 8527 15855 8585 15861
rect 8938 15852 8944 15864
rect 8996 15852 9002 15904
rect 9582 15852 9588 15904
rect 9640 15892 9646 15904
rect 10042 15892 10048 15904
rect 9640 15864 10048 15892
rect 9640 15852 9646 15864
rect 10042 15852 10048 15864
rect 10100 15892 10106 15904
rect 10413 15895 10471 15901
rect 10413 15892 10425 15895
rect 10100 15864 10425 15892
rect 10100 15852 10106 15864
rect 10413 15861 10425 15864
rect 10459 15861 10471 15895
rect 10413 15855 10471 15861
rect 10778 15852 10784 15904
rect 10836 15892 10842 15904
rect 11103 15895 11161 15901
rect 11103 15892 11115 15895
rect 10836 15864 11115 15892
rect 10836 15852 10842 15864
rect 11103 15861 11115 15864
rect 11149 15861 11161 15895
rect 11103 15855 11161 15861
rect 1104 15802 17756 15824
rect 1104 15750 7288 15802
rect 7340 15750 7352 15802
rect 7404 15750 7416 15802
rect 7468 15750 7480 15802
rect 7532 15750 13595 15802
rect 13647 15750 13659 15802
rect 13711 15750 13723 15802
rect 13775 15750 13787 15802
rect 13839 15750 17756 15802
rect 1104 15728 17756 15750
rect 2130 15580 2136 15632
rect 2188 15620 2194 15632
rect 2409 15623 2467 15629
rect 2409 15620 2421 15623
rect 2188 15592 2421 15620
rect 2188 15580 2194 15592
rect 2409 15589 2421 15592
rect 2455 15589 2467 15623
rect 2409 15583 2467 15589
rect 6089 15623 6147 15629
rect 6089 15589 6101 15623
rect 6135 15620 6147 15623
rect 6178 15620 6184 15632
rect 6135 15592 6184 15620
rect 6135 15589 6147 15592
rect 6089 15583 6147 15589
rect 6178 15580 6184 15592
rect 6236 15620 6242 15632
rect 7837 15623 7895 15629
rect 6236 15592 6776 15620
rect 6236 15580 6242 15592
rect 1762 15484 1768 15496
rect 1675 15456 1768 15484
rect 1762 15444 1768 15456
rect 1820 15484 1826 15496
rect 4065 15487 4123 15493
rect 4065 15484 4077 15487
rect 1820 15456 4077 15484
rect 1820 15444 1826 15456
rect 4065 15453 4077 15456
rect 4111 15453 4123 15487
rect 6546 15484 6552 15496
rect 6507 15456 6552 15484
rect 4065 15447 4123 15453
rect 6546 15444 6552 15456
rect 6604 15444 6610 15496
rect 6748 15484 6776 15592
rect 7837 15589 7849 15623
rect 7883 15620 7895 15623
rect 8110 15620 8116 15632
rect 7883 15592 8116 15620
rect 7883 15589 7895 15592
rect 7837 15583 7895 15589
rect 8110 15580 8116 15592
rect 8168 15580 8174 15632
rect 8202 15580 8208 15632
rect 8260 15620 8266 15632
rect 11149 15623 11207 15629
rect 11149 15620 11161 15623
rect 8260 15592 11161 15620
rect 8260 15580 8266 15592
rect 11149 15589 11161 15592
rect 11195 15589 11207 15623
rect 11149 15583 11207 15589
rect 8113 15487 8171 15493
rect 8113 15484 8125 15487
rect 6748 15456 8125 15484
rect 8113 15453 8125 15456
rect 8159 15453 8171 15487
rect 8113 15447 8171 15453
rect 10318 15444 10324 15496
rect 10376 15484 10382 15496
rect 10505 15487 10563 15493
rect 10505 15484 10517 15487
rect 10376 15456 10517 15484
rect 10376 15444 10382 15456
rect 10505 15453 10517 15456
rect 10551 15453 10563 15487
rect 15838 15484 15844 15496
rect 15799 15456 15844 15484
rect 10505 15447 10563 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16114 15484 16120 15496
rect 16075 15456 16120 15484
rect 16114 15444 16120 15456
rect 16172 15444 16178 15496
rect 1104 15258 17756 15280
rect 1104 15206 4135 15258
rect 4187 15206 4199 15258
rect 4251 15206 4263 15258
rect 4315 15206 4327 15258
rect 4379 15206 10441 15258
rect 10493 15206 10505 15258
rect 10557 15206 10569 15258
rect 10621 15206 10633 15258
rect 10685 15206 16748 15258
rect 16800 15206 16812 15258
rect 16864 15206 16876 15258
rect 16928 15206 16940 15258
rect 16992 15206 17756 15258
rect 1104 15184 17756 15206
rect 1762 15144 1768 15156
rect 1723 15116 1768 15144
rect 1762 15104 1768 15116
rect 1820 15104 1826 15156
rect 6178 15144 6184 15156
rect 5736 15116 6184 15144
rect 5736 15085 5764 15116
rect 6178 15104 6184 15116
rect 6236 15104 6242 15156
rect 7837 15147 7895 15153
rect 7837 15113 7849 15147
rect 7883 15144 7895 15147
rect 8110 15144 8116 15156
rect 7883 15116 8116 15144
rect 7883 15113 7895 15116
rect 7837 15107 7895 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 10318 15104 10324 15156
rect 10376 15144 10382 15156
rect 10413 15147 10471 15153
rect 10413 15144 10425 15147
rect 10376 15116 10425 15144
rect 10376 15104 10382 15116
rect 10413 15113 10425 15116
rect 10459 15144 10471 15147
rect 10735 15147 10793 15153
rect 10735 15144 10747 15147
rect 10459 15116 10747 15144
rect 10459 15113 10471 15116
rect 10413 15107 10471 15113
rect 10735 15113 10747 15116
rect 10781 15113 10793 15147
rect 15838 15144 15844 15156
rect 15799 15116 15844 15144
rect 10735 15107 10793 15113
rect 15838 15104 15844 15116
rect 15896 15144 15902 15156
rect 16255 15147 16313 15153
rect 16255 15144 16267 15147
rect 15896 15116 16267 15144
rect 15896 15104 15902 15116
rect 16255 15113 16267 15116
rect 16301 15113 16313 15147
rect 16255 15107 16313 15113
rect 5721 15079 5779 15085
rect 5721 15045 5733 15079
rect 5767 15045 5779 15079
rect 5721 15039 5779 15045
rect 1670 14968 1676 15020
rect 1728 15008 1734 15020
rect 1949 15011 2007 15017
rect 1949 15008 1961 15011
rect 1728 14980 1961 15008
rect 1728 14968 1734 14980
rect 1949 14977 1961 14980
rect 1995 15008 2007 15011
rect 2869 15011 2927 15017
rect 2869 15008 2881 15011
rect 1995 14980 2881 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2869 14977 2881 14980
rect 2915 14977 2927 15011
rect 2869 14971 2927 14977
rect 4249 15011 4307 15017
rect 4249 14977 4261 15011
rect 4295 15008 4307 15011
rect 4430 15008 4436 15020
rect 4295 14980 4436 15008
rect 4295 14977 4307 14980
rect 4249 14971 4307 14977
rect 4430 14968 4436 14980
rect 4488 14968 4494 15020
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 6825 15011 6883 15017
rect 6825 15008 6837 15011
rect 6788 14980 6837 15008
rect 6788 14968 6794 14980
rect 6825 14977 6837 14980
rect 6871 14977 6883 15011
rect 9582 15008 9588 15020
rect 9543 14980 9588 15008
rect 6825 14971 6883 14977
rect 9582 14968 9588 14980
rect 9640 14968 9646 15020
rect 10664 14943 10722 14949
rect 10664 14909 10676 14943
rect 10710 14940 10722 14943
rect 16184 14943 16242 14949
rect 10710 14912 11100 14940
rect 10710 14909 10722 14912
rect 10664 14903 10722 14909
rect 2590 14872 2596 14884
rect 2551 14844 2596 14872
rect 2590 14832 2596 14844
rect 2648 14832 2654 14884
rect 3421 14875 3479 14881
rect 3421 14841 3433 14875
rect 3467 14872 3479 14875
rect 3602 14872 3608 14884
rect 3467 14844 3608 14872
rect 3467 14841 3479 14844
rect 3421 14835 3479 14841
rect 3602 14832 3608 14844
rect 3660 14832 3666 14884
rect 4985 14875 5043 14881
rect 4985 14841 4997 14875
rect 5031 14872 5043 14875
rect 5166 14872 5172 14884
rect 5031 14844 5172 14872
rect 5031 14841 5043 14844
rect 4985 14835 5043 14841
rect 5166 14832 5172 14844
rect 5224 14832 5230 14884
rect 11072 14816 11100 14912
rect 16184 14909 16196 14943
rect 16230 14940 16242 14943
rect 16230 14912 16528 14940
rect 16230 14909 16242 14912
rect 16184 14903 16242 14909
rect 16500 14816 16528 14912
rect 11054 14804 11060 14816
rect 11015 14776 11060 14804
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 16482 14764 16488 14816
rect 16540 14804 16546 14816
rect 16577 14807 16635 14813
rect 16577 14804 16589 14807
rect 16540 14776 16589 14804
rect 16540 14764 16546 14776
rect 16577 14773 16589 14776
rect 16623 14773 16635 14807
rect 16577 14767 16635 14773
rect 1104 14714 17756 14736
rect 1104 14662 7288 14714
rect 7340 14662 7352 14714
rect 7404 14662 7416 14714
rect 7468 14662 7480 14714
rect 7532 14662 13595 14714
rect 13647 14662 13659 14714
rect 13711 14662 13723 14714
rect 13775 14662 13787 14714
rect 13839 14662 17756 14714
rect 1104 14640 17756 14662
rect 2590 14600 2596 14612
rect 2551 14572 2596 14600
rect 2590 14560 2596 14572
rect 2648 14560 2654 14612
rect 5166 14560 5172 14612
rect 5224 14600 5230 14612
rect 5767 14603 5825 14609
rect 5767 14600 5779 14603
rect 5224 14572 5779 14600
rect 5224 14560 5230 14572
rect 5767 14569 5779 14572
rect 5813 14569 5825 14603
rect 5767 14563 5825 14569
rect 6638 14560 6644 14612
rect 6696 14600 6702 14612
rect 6779 14603 6837 14609
rect 6779 14600 6791 14603
rect 6696 14572 6791 14600
rect 6696 14560 6702 14572
rect 6779 14569 6791 14572
rect 6825 14569 6837 14603
rect 6779 14563 6837 14569
rect 2222 14532 2228 14544
rect 2183 14504 2228 14532
rect 2222 14492 2228 14504
rect 2280 14492 2286 14544
rect 5626 14464 5632 14476
rect 5587 14436 5632 14464
rect 5626 14424 5632 14436
rect 5684 14424 5690 14476
rect 6708 14467 6766 14473
rect 6708 14433 6720 14467
rect 6754 14464 6766 14467
rect 7098 14464 7104 14476
rect 6754 14436 7104 14464
rect 6754 14433 6766 14436
rect 6708 14427 6766 14433
rect 7098 14424 7104 14436
rect 7156 14464 7162 14476
rect 12434 14464 12440 14476
rect 7156 14436 12440 14464
rect 7156 14424 7162 14436
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 2222 14396 2228 14408
rect 1627 14368 2228 14396
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 2222 14356 2228 14368
rect 2280 14356 2286 14408
rect 3970 14356 3976 14408
rect 4028 14396 4034 14408
rect 4157 14399 4215 14405
rect 4157 14396 4169 14399
rect 4028 14368 4169 14396
rect 4028 14356 4034 14368
rect 4157 14365 4169 14368
rect 4203 14365 4215 14399
rect 4157 14359 4215 14365
rect 2590 14288 2596 14340
rect 2648 14328 2654 14340
rect 4709 14331 4767 14337
rect 4709 14328 4721 14331
rect 2648 14300 4721 14328
rect 2648 14288 2654 14300
rect 4709 14297 4721 14300
rect 4755 14297 4767 14331
rect 4709 14291 4767 14297
rect 1104 14170 17756 14192
rect 1104 14118 4135 14170
rect 4187 14118 4199 14170
rect 4251 14118 4263 14170
rect 4315 14118 4327 14170
rect 4379 14118 10441 14170
rect 10493 14118 10505 14170
rect 10557 14118 10569 14170
rect 10621 14118 10633 14170
rect 10685 14118 16748 14170
rect 16800 14118 16812 14170
rect 16864 14118 16876 14170
rect 16928 14118 16940 14170
rect 16992 14118 17756 14170
rect 1104 14096 17756 14118
rect 3970 14016 3976 14068
rect 4028 14056 4034 14068
rect 4065 14059 4123 14065
rect 4065 14056 4077 14059
rect 4028 14028 4077 14056
rect 4028 14016 4034 14028
rect 4065 14025 4077 14028
rect 4111 14056 4123 14059
rect 4295 14059 4353 14065
rect 4295 14056 4307 14059
rect 4111 14028 4307 14056
rect 4111 14025 4123 14028
rect 4065 14019 4123 14025
rect 4295 14025 4307 14028
rect 4341 14025 4353 14059
rect 7098 14056 7104 14068
rect 7059 14028 7104 14056
rect 4295 14019 4353 14025
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 106 13948 112 14000
rect 164 13988 170 14000
rect 5626 13988 5632 14000
rect 164 13960 5632 13988
rect 164 13948 170 13960
rect 5626 13948 5632 13960
rect 5684 13948 5690 14000
rect 1857 13923 1915 13929
rect 1857 13920 1869 13923
rect 1447 13892 1869 13920
rect 1118 13812 1124 13864
rect 1176 13852 1182 13864
rect 1447 13861 1475 13892
rect 1857 13889 1869 13892
rect 1903 13889 1915 13923
rect 2682 13920 2688 13932
rect 2643 13892 2688 13920
rect 1857 13883 1915 13889
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 2958 13920 2964 13932
rect 2919 13892 2964 13920
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13920 4767 13923
rect 8662 13920 8668 13932
rect 4755 13892 8668 13920
rect 4755 13889 4767 13892
rect 4709 13883 4767 13889
rect 1432 13855 1490 13861
rect 1432 13852 1444 13855
rect 1176 13824 1444 13852
rect 1176 13812 1182 13824
rect 1432 13821 1444 13824
rect 1478 13821 1490 13855
rect 1432 13815 1490 13821
rect 1535 13855 1593 13861
rect 1535 13821 1547 13855
rect 1581 13852 1593 13855
rect 1670 13852 1676 13864
rect 1581 13824 1676 13852
rect 1581 13821 1593 13824
rect 1535 13815 1593 13821
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 4224 13855 4282 13861
rect 4224 13821 4236 13855
rect 4270 13852 4282 13855
rect 4724 13852 4752 13883
rect 8662 13880 8668 13892
rect 8720 13880 8726 13932
rect 4270 13824 4752 13852
rect 4270 13821 4282 13824
rect 4224 13815 4282 13821
rect 4982 13812 4988 13864
rect 5040 13852 5046 13864
rect 5204 13855 5262 13861
rect 5204 13852 5216 13855
rect 5040 13824 5216 13852
rect 5040 13812 5046 13824
rect 5204 13821 5216 13824
rect 5250 13852 5262 13855
rect 5997 13855 6055 13861
rect 5997 13852 6009 13855
rect 5250 13824 6009 13852
rect 5250 13821 5262 13824
rect 5204 13815 5262 13821
rect 5997 13821 6009 13824
rect 6043 13821 6055 13855
rect 5997 13815 6055 13821
rect 2314 13744 2320 13796
rect 2372 13784 2378 13796
rect 5307 13787 5365 13793
rect 5307 13784 5319 13787
rect 2372 13756 5319 13784
rect 2372 13744 2378 13756
rect 5307 13753 5319 13756
rect 5353 13753 5365 13787
rect 5307 13747 5365 13753
rect 2222 13716 2228 13728
rect 2183 13688 2228 13716
rect 2222 13676 2228 13688
rect 2280 13676 2286 13728
rect 1104 13626 17756 13648
rect 1104 13574 7288 13626
rect 7340 13574 7352 13626
rect 7404 13574 7416 13626
rect 7468 13574 7480 13626
rect 7532 13574 13595 13626
rect 13647 13574 13659 13626
rect 13711 13574 13723 13626
rect 13775 13574 13787 13626
rect 13839 13574 17756 13626
rect 1104 13552 17756 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 3602 13472 3608 13524
rect 3660 13512 3666 13524
rect 4203 13515 4261 13521
rect 4203 13512 4215 13515
rect 3660 13484 4215 13512
rect 3660 13472 3666 13484
rect 4203 13481 4215 13484
rect 4249 13481 4261 13515
rect 4203 13475 4261 13481
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 2038 13376 2044 13388
rect 1443 13348 2044 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 2038 13336 2044 13348
rect 2096 13336 2102 13388
rect 2568 13379 2626 13385
rect 2568 13345 2580 13379
rect 2614 13376 2626 13379
rect 2958 13376 2964 13388
rect 2614 13348 2964 13376
rect 2614 13345 2626 13348
rect 2568 13339 2626 13345
rect 2958 13336 2964 13348
rect 3016 13336 3022 13388
rect 3970 13336 3976 13388
rect 4028 13376 4034 13388
rect 4100 13379 4158 13385
rect 4100 13376 4112 13379
rect 4028 13348 4112 13376
rect 4028 13336 4034 13348
rect 4100 13345 4112 13348
rect 4146 13345 4158 13379
rect 4100 13339 4158 13345
rect 16092 13379 16150 13385
rect 16092 13345 16104 13379
rect 16138 13376 16150 13379
rect 16206 13376 16212 13388
rect 16138 13348 16212 13376
rect 16138 13345 16150 13348
rect 16092 13339 16150 13345
rect 16206 13336 16212 13348
rect 16264 13336 16270 13388
rect 2038 13172 2044 13184
rect 1999 13144 2044 13172
rect 2038 13132 2044 13144
rect 2096 13132 2102 13184
rect 2498 13132 2504 13184
rect 2556 13172 2562 13184
rect 2639 13175 2697 13181
rect 2639 13172 2651 13175
rect 2556 13144 2651 13172
rect 2556 13132 2562 13144
rect 2639 13141 2651 13144
rect 2685 13141 2697 13175
rect 2639 13135 2697 13141
rect 16163 13175 16221 13181
rect 16163 13141 16175 13175
rect 16209 13172 16221 13175
rect 16298 13172 16304 13184
rect 16209 13144 16304 13172
rect 16209 13141 16221 13144
rect 16163 13135 16221 13141
rect 16298 13132 16304 13144
rect 16356 13132 16362 13184
rect 1104 13082 17756 13104
rect 1104 13030 4135 13082
rect 4187 13030 4199 13082
rect 4251 13030 4263 13082
rect 4315 13030 4327 13082
rect 4379 13030 10441 13082
rect 10493 13030 10505 13082
rect 10557 13030 10569 13082
rect 10621 13030 10633 13082
rect 10685 13030 16748 13082
rect 16800 13030 16812 13082
rect 16864 13030 16876 13082
rect 16928 13030 16940 13082
rect 16992 13030 17756 13082
rect 1104 13008 17756 13030
rect 1535 12971 1593 12977
rect 1535 12937 1547 12971
rect 1581 12968 1593 12971
rect 2222 12968 2228 12980
rect 1581 12940 2228 12968
rect 1581 12937 1593 12940
rect 1535 12931 1593 12937
rect 2222 12928 2228 12940
rect 2280 12928 2286 12980
rect 16117 12971 16175 12977
rect 16117 12937 16129 12971
rect 16163 12968 16175 12971
rect 16206 12968 16212 12980
rect 16163 12940 16212 12968
rect 16163 12937 16175 12940
rect 16117 12931 16175 12937
rect 16206 12928 16212 12940
rect 16264 12928 16270 12980
rect 2958 12860 2964 12912
rect 3016 12900 3022 12912
rect 3053 12903 3111 12909
rect 3053 12900 3065 12903
rect 3016 12872 3065 12900
rect 3016 12860 3022 12872
rect 3053 12869 3065 12872
rect 3099 12869 3111 12903
rect 3053 12863 3111 12869
rect 16485 12903 16543 12909
rect 16485 12869 16497 12903
rect 16531 12900 16543 12903
rect 18414 12900 18420 12912
rect 16531 12872 18420 12900
rect 16531 12869 16543 12872
rect 16485 12863 16543 12869
rect 18414 12860 18420 12872
rect 18472 12860 18478 12912
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 2501 12835 2559 12841
rect 2501 12832 2513 12835
rect 2363 12804 2513 12832
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 2501 12801 2513 12804
rect 2547 12832 2559 12835
rect 3973 12835 4031 12841
rect 3973 12832 3985 12835
rect 2547 12804 3985 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 3973 12801 3985 12804
rect 4019 12801 4031 12835
rect 3973 12795 4031 12801
rect 1464 12767 1522 12773
rect 1464 12733 1476 12767
rect 1510 12764 1522 12767
rect 1854 12764 1860 12776
rect 1510 12736 1860 12764
rect 1510 12733 1522 12736
rect 1464 12727 1522 12733
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5123 12736 5764 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5736 12640 5764 12736
rect 13170 12724 13176 12776
rect 13228 12764 13234 12776
rect 13668 12767 13726 12773
rect 13668 12764 13680 12767
rect 13228 12736 13680 12764
rect 13228 12724 13234 12736
rect 13668 12733 13680 12736
rect 13714 12764 13726 12767
rect 14093 12767 14151 12773
rect 14093 12764 14105 12767
rect 13714 12736 14105 12764
rect 13714 12733 13726 12736
rect 13668 12727 13726 12733
rect 14093 12733 14105 12736
rect 14139 12733 14151 12767
rect 16298 12764 16304 12776
rect 16259 12736 16304 12764
rect 14093 12727 14151 12733
rect 16298 12724 16304 12736
rect 16356 12764 16362 12776
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 16356 12736 16865 12764
rect 16356 12724 16362 12736
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 3970 12628 3976 12640
rect 2832 12600 3976 12628
rect 2832 12588 2838 12600
rect 3970 12588 3976 12600
rect 4028 12628 4034 12640
rect 4433 12631 4491 12637
rect 4433 12628 4445 12631
rect 4028 12600 4445 12628
rect 4028 12588 4034 12600
rect 4433 12597 4445 12600
rect 4479 12597 4491 12631
rect 5258 12628 5264 12640
rect 5219 12600 5264 12628
rect 4433 12591 4491 12597
rect 5258 12588 5264 12600
rect 5316 12588 5322 12640
rect 5718 12628 5724 12640
rect 5679 12600 5724 12628
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 13771 12631 13829 12637
rect 13771 12597 13783 12631
rect 13817 12628 13829 12631
rect 15102 12628 15108 12640
rect 13817 12600 15108 12628
rect 13817 12597 13829 12600
rect 13771 12591 13829 12597
rect 15102 12588 15108 12600
rect 15160 12588 15166 12640
rect 15286 12628 15292 12640
rect 15247 12600 15292 12628
rect 15286 12588 15292 12600
rect 15344 12588 15350 12640
rect 1104 12538 17756 12560
rect 1104 12486 7288 12538
rect 7340 12486 7352 12538
rect 7404 12486 7416 12538
rect 7468 12486 7480 12538
rect 7532 12486 13595 12538
rect 13647 12486 13659 12538
rect 13711 12486 13723 12538
rect 13775 12486 13787 12538
rect 13839 12486 17756 12538
rect 1104 12464 17756 12486
rect 2593 12427 2651 12433
rect 2593 12393 2605 12427
rect 2639 12424 2651 12427
rect 2958 12424 2964 12436
rect 2639 12396 2964 12424
rect 2639 12393 2651 12396
rect 2593 12387 2651 12393
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 5718 12384 5724 12436
rect 5776 12424 5782 12436
rect 6227 12427 6285 12433
rect 6227 12424 6239 12427
rect 5776 12396 6239 12424
rect 5776 12384 5782 12396
rect 6227 12393 6239 12396
rect 6273 12393 6285 12427
rect 6227 12387 6285 12393
rect 2038 12316 2044 12368
rect 2096 12356 2102 12368
rect 5215 12359 5273 12365
rect 5215 12356 5227 12359
rect 2096 12328 5227 12356
rect 2096 12316 2102 12328
rect 5215 12325 5227 12328
rect 5261 12325 5273 12359
rect 5215 12319 5273 12325
rect 15102 12316 15108 12368
rect 15160 12356 15166 12368
rect 15381 12359 15439 12365
rect 15381 12356 15393 12359
rect 15160 12328 15393 12356
rect 15160 12316 15166 12328
rect 15381 12325 15393 12328
rect 15427 12325 15439 12359
rect 15381 12319 15439 12325
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 2498 12288 2504 12300
rect 1995 12260 2504 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 5074 12288 5080 12300
rect 5035 12260 5080 12288
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 6156 12291 6214 12297
rect 6156 12257 6168 12291
rect 6202 12288 6214 12291
rect 6270 12288 6276 12300
rect 6202 12260 6276 12288
rect 6202 12257 6214 12260
rect 6156 12251 6214 12257
rect 6270 12248 6276 12260
rect 6328 12248 6334 12300
rect 3878 12180 3884 12232
rect 3936 12220 3942 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 3936 12192 4077 12220
rect 3936 12180 3942 12192
rect 4065 12189 4077 12192
rect 4111 12189 4123 12223
rect 15746 12220 15752 12232
rect 15707 12192 15752 12220
rect 4065 12183 4123 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 106 12112 112 12164
rect 164 12152 170 12164
rect 2133 12155 2191 12161
rect 2133 12152 2145 12155
rect 164 12124 2145 12152
rect 164 12112 170 12124
rect 2133 12121 2145 12124
rect 2179 12121 2191 12155
rect 2133 12115 2191 12121
rect 1578 12084 1584 12096
rect 1539 12056 1584 12084
rect 1578 12044 1584 12056
rect 1636 12044 1642 12096
rect 1104 11994 17756 12016
rect 1104 11942 4135 11994
rect 4187 11942 4199 11994
rect 4251 11942 4263 11994
rect 4315 11942 4327 11994
rect 4379 11942 10441 11994
rect 10493 11942 10505 11994
rect 10557 11942 10569 11994
rect 10621 11942 10633 11994
rect 10685 11942 16748 11994
rect 16800 11942 16812 11994
rect 16864 11942 16876 11994
rect 16928 11942 16940 11994
rect 16992 11942 17756 11994
rect 1104 11920 17756 11942
rect 2498 11880 2504 11892
rect 2459 11852 2504 11880
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 6181 11883 6239 11889
rect 6181 11880 6193 11883
rect 4448 11852 6193 11880
rect 4448 11821 4476 11852
rect 6181 11849 6193 11852
rect 6227 11880 6239 11883
rect 6270 11880 6276 11892
rect 6227 11852 6276 11880
rect 6227 11849 6239 11852
rect 6181 11843 6239 11849
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 14182 11880 14188 11892
rect 14143 11852 14188 11880
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 15102 11880 15108 11892
rect 15063 11852 15108 11880
rect 15102 11840 15108 11852
rect 15160 11840 15166 11892
rect 15286 11840 15292 11892
rect 15344 11880 15350 11892
rect 15473 11883 15531 11889
rect 15473 11880 15485 11883
rect 15344 11852 15485 11880
rect 15344 11840 15350 11852
rect 15473 11849 15485 11852
rect 15519 11880 15531 11883
rect 15519 11852 15792 11880
rect 15519 11849 15531 11852
rect 15473 11843 15531 11849
rect 4433 11815 4491 11821
rect 4433 11812 4445 11815
rect 4126 11784 4445 11812
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11744 1547 11747
rect 1578 11744 1584 11756
rect 1535 11716 1584 11744
rect 1535 11713 1547 11716
rect 1489 11707 1547 11713
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 3697 11747 3755 11753
rect 3697 11713 3709 11747
rect 3743 11744 3755 11747
rect 3878 11744 3884 11756
rect 3743 11716 3884 11744
rect 3743 11713 3755 11716
rect 3697 11707 3755 11713
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 3970 11704 3976 11756
rect 4028 11744 4034 11756
rect 4126 11744 4154 11784
rect 4433 11781 4445 11784
rect 4479 11781 4491 11815
rect 4433 11775 4491 11781
rect 15764 11753 15792 11852
rect 4028 11716 4154 11744
rect 15749 11747 15807 11753
rect 4028 11704 4034 11716
rect 15749 11713 15761 11747
rect 15795 11713 15807 11747
rect 16206 11744 16212 11756
rect 16167 11716 16212 11744
rect 15749 11707 15807 11713
rect 16206 11704 16212 11716
rect 16264 11704 16270 11756
rect 14001 11679 14059 11685
rect 14001 11645 14013 11679
rect 14047 11676 14059 11679
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 14047 11648 14565 11676
rect 14047 11645 14059 11648
rect 14001 11639 14059 11645
rect 14553 11645 14565 11648
rect 14599 11676 14611 11679
rect 14642 11676 14648 11688
rect 14599 11648 14648 11676
rect 14599 11645 14611 11648
rect 14553 11639 14611 11645
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 2133 11611 2191 11617
rect 2133 11577 2145 11611
rect 2179 11608 2191 11611
rect 2314 11608 2320 11620
rect 2179 11580 2320 11608
rect 2179 11577 2191 11580
rect 2133 11571 2191 11577
rect 2314 11568 2320 11580
rect 2372 11608 2378 11620
rect 2372 11580 4154 11608
rect 2372 11568 2378 11580
rect 4126 11540 4154 11580
rect 5074 11540 5080 11552
rect 4126 11512 5080 11540
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 1104 11450 17756 11472
rect 1104 11398 7288 11450
rect 7340 11398 7352 11450
rect 7404 11398 7416 11450
rect 7468 11398 7480 11450
rect 7532 11398 13595 11450
rect 13647 11398 13659 11450
rect 13711 11398 13723 11450
rect 13775 11398 13787 11450
rect 13839 11398 17756 11450
rect 1104 11376 17756 11398
rect 2314 11268 2320 11280
rect 2275 11240 2320 11268
rect 2314 11228 2320 11240
rect 2372 11228 2378 11280
rect 15746 11268 15752 11280
rect 15707 11240 15752 11268
rect 15746 11228 15752 11240
rect 15804 11228 15810 11280
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11132 1731 11135
rect 2130 11132 2136 11144
rect 1719 11104 2136 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 16206 11132 16212 11144
rect 16167 11104 16212 11132
rect 16206 11092 16212 11104
rect 16264 11092 16270 11144
rect 1104 10906 17756 10928
rect 1104 10854 4135 10906
rect 4187 10854 4199 10906
rect 4251 10854 4263 10906
rect 4315 10854 4327 10906
rect 4379 10854 10441 10906
rect 10493 10854 10505 10906
rect 10557 10854 10569 10906
rect 10621 10854 10633 10906
rect 10685 10854 16748 10906
rect 16800 10854 16812 10906
rect 16864 10854 16876 10906
rect 16928 10854 16940 10906
rect 16992 10854 17756 10906
rect 1104 10832 17756 10854
rect 14642 10792 14648 10804
rect 14603 10764 14648 10792
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 15289 10727 15347 10733
rect 15289 10693 15301 10727
rect 15335 10724 15347 10727
rect 15746 10724 15752 10736
rect 15335 10696 15752 10724
rect 15335 10693 15347 10696
rect 15289 10687 15347 10693
rect 15746 10684 15752 10696
rect 15804 10724 15810 10736
rect 15804 10696 16160 10724
rect 15804 10684 15810 10696
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10656 3939 10659
rect 3970 10656 3976 10668
rect 3927 10628 3976 10656
rect 3927 10625 3939 10628
rect 3881 10619 3939 10625
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 14451 10628 14933 10656
rect 4776 10591 4834 10597
rect 4776 10557 4788 10591
rect 4822 10588 4834 10591
rect 5166 10588 5172 10600
rect 4822 10560 5172 10588
rect 4822 10557 4834 10560
rect 4776 10551 4834 10557
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 14451 10597 14479 10628
rect 14921 10625 14933 10628
rect 14967 10656 14979 10659
rect 15930 10656 15936 10668
rect 14967 10628 15936 10656
rect 14967 10625 14979 10628
rect 14921 10619 14979 10625
rect 15930 10616 15936 10628
rect 15988 10616 15994 10668
rect 16132 10665 16160 10696
rect 16117 10659 16175 10665
rect 16117 10625 16129 10659
rect 16163 10625 16175 10659
rect 16117 10619 16175 10625
rect 14436 10591 14494 10597
rect 14436 10557 14448 10591
rect 14482 10557 14494 10591
rect 14436 10551 14494 10557
rect 1670 10520 1676 10532
rect 1631 10492 1676 10520
rect 1670 10480 1676 10492
rect 1728 10480 1734 10532
rect 2314 10520 2320 10532
rect 2275 10492 2320 10520
rect 2314 10480 2320 10492
rect 2372 10520 2378 10532
rect 2961 10523 3019 10529
rect 2961 10520 2973 10523
rect 2372 10492 2973 10520
rect 2372 10480 2378 10492
rect 2961 10489 2973 10492
rect 3007 10520 3019 10523
rect 3237 10523 3295 10529
rect 3237 10520 3249 10523
rect 3007 10492 3249 10520
rect 3007 10489 3019 10492
rect 2961 10483 3019 10489
rect 3237 10489 3249 10492
rect 3283 10489 3295 10523
rect 3237 10483 3295 10489
rect 15841 10523 15899 10529
rect 15841 10489 15853 10523
rect 15887 10489 15899 10523
rect 15841 10483 15899 10489
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 2593 10455 2651 10461
rect 2593 10452 2605 10455
rect 2188 10424 2605 10452
rect 2188 10412 2194 10424
rect 2593 10421 2605 10424
rect 2639 10421 2651 10455
rect 2593 10415 2651 10421
rect 3050 10412 3056 10464
rect 3108 10452 3114 10464
rect 4847 10455 4905 10461
rect 4847 10452 4859 10455
rect 3108 10424 4859 10452
rect 3108 10412 3114 10424
rect 4847 10421 4859 10424
rect 4893 10421 4905 10455
rect 15562 10452 15568 10464
rect 15523 10424 15568 10452
rect 4847 10415 4905 10421
rect 15562 10412 15568 10424
rect 15620 10452 15626 10464
rect 15856 10452 15884 10483
rect 15620 10424 15884 10452
rect 15620 10412 15626 10424
rect 1104 10362 17756 10384
rect 1104 10310 7288 10362
rect 7340 10310 7352 10362
rect 7404 10310 7416 10362
rect 7468 10310 7480 10362
rect 7532 10310 13595 10362
rect 13647 10310 13659 10362
rect 13711 10310 13723 10362
rect 13775 10310 13787 10362
rect 13839 10310 17756 10362
rect 1104 10288 17756 10310
rect 1397 10251 1455 10257
rect 1397 10217 1409 10251
rect 1443 10248 1455 10251
rect 1578 10248 1584 10260
rect 1443 10220 1584 10248
rect 1443 10217 1455 10220
rect 1397 10211 1455 10217
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 1670 10208 1676 10260
rect 1728 10248 1734 10260
rect 1949 10251 2007 10257
rect 1949 10248 1961 10251
rect 1728 10220 1961 10248
rect 1728 10208 1734 10220
rect 1949 10217 1961 10220
rect 1995 10248 2007 10251
rect 3050 10248 3056 10260
rect 1995 10220 3056 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 14323 10251 14381 10257
rect 14323 10217 14335 10251
rect 14369 10248 14381 10251
rect 15562 10248 15568 10260
rect 14369 10220 15568 10248
rect 14369 10217 14381 10220
rect 14323 10211 14381 10217
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 106 10072 112 10124
rect 164 10112 170 10124
rect 2498 10121 2504 10124
rect 2444 10115 2504 10121
rect 2444 10112 2456 10115
rect 164 10084 2456 10112
rect 164 10072 170 10084
rect 2444 10081 2456 10084
rect 2490 10081 2504 10115
rect 2444 10075 2504 10081
rect 2498 10072 2504 10075
rect 2556 10072 2562 10124
rect 14093 10115 14151 10121
rect 14093 10081 14105 10115
rect 14139 10112 14151 10115
rect 14274 10112 14280 10124
rect 14139 10084 14280 10112
rect 14139 10081 14151 10084
rect 14093 10075 14151 10081
rect 14274 10072 14280 10084
rect 14332 10072 14338 10124
rect 15378 10044 15384 10056
rect 15339 10016 15384 10044
rect 15378 10004 15384 10016
rect 15436 10004 15442 10056
rect 15930 9976 15936 9988
rect 15891 9948 15936 9976
rect 15930 9936 15936 9948
rect 15988 9936 15994 9988
rect 1946 9868 1952 9920
rect 2004 9908 2010 9920
rect 2317 9911 2375 9917
rect 2317 9908 2329 9911
rect 2004 9880 2329 9908
rect 2004 9868 2010 9880
rect 2317 9877 2329 9880
rect 2363 9908 2375 9911
rect 2547 9911 2605 9917
rect 2547 9908 2559 9911
rect 2363 9880 2559 9908
rect 2363 9877 2375 9880
rect 2317 9871 2375 9877
rect 2547 9877 2559 9880
rect 2593 9877 2605 9911
rect 2547 9871 2605 9877
rect 1104 9818 17756 9840
rect 1104 9766 4135 9818
rect 4187 9766 4199 9818
rect 4251 9766 4263 9818
rect 4315 9766 4327 9818
rect 4379 9766 10441 9818
rect 10493 9766 10505 9818
rect 10557 9766 10569 9818
rect 10621 9766 10633 9818
rect 10685 9766 16748 9818
rect 16800 9766 16812 9818
rect 16864 9766 16876 9818
rect 16928 9766 16940 9818
rect 16992 9766 17756 9818
rect 1104 9744 17756 9766
rect 15378 9704 15384 9716
rect 15339 9676 15384 9704
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 2406 9636 2412 9648
rect 2367 9608 2412 9636
rect 2406 9596 2412 9608
rect 2464 9596 2470 9648
rect 1489 9571 1547 9577
rect 1489 9537 1501 9571
rect 1535 9568 1547 9571
rect 1946 9568 1952 9580
rect 1535 9540 1952 9568
rect 1535 9537 1547 9540
rect 1489 9531 1547 9537
rect 1946 9528 1952 9540
rect 2004 9528 2010 9580
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 15396 9568 15424 9664
rect 15930 9568 15936 9580
rect 14507 9540 15424 9568
rect 15891 9540 15936 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 15930 9528 15936 9540
rect 15988 9528 15994 9580
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 3028 9503 3086 9509
rect 3028 9500 3040 9503
rect 2740 9472 3040 9500
rect 2740 9460 2746 9472
rect 3028 9469 3040 9472
rect 3074 9500 3086 9503
rect 3421 9503 3479 9509
rect 3421 9500 3433 9503
rect 3074 9472 3433 9500
rect 3074 9469 3086 9472
rect 3028 9463 3086 9469
rect 3421 9469 3433 9472
rect 3467 9469 3479 9503
rect 3421 9463 3479 9469
rect 2130 9432 2136 9444
rect 2091 9404 2136 9432
rect 2130 9392 2136 9404
rect 2188 9392 2194 9444
rect 15562 9432 15568 9444
rect 15523 9404 15568 9432
rect 15562 9392 15568 9404
rect 15620 9392 15626 9444
rect 2498 9324 2504 9376
rect 2556 9364 2562 9376
rect 3099 9367 3157 9373
rect 3099 9364 3111 9367
rect 2556 9336 3111 9364
rect 2556 9324 2562 9336
rect 3099 9333 3111 9336
rect 3145 9333 3157 9367
rect 14274 9364 14280 9376
rect 14235 9336 14280 9364
rect 3099 9327 3157 9333
rect 14274 9324 14280 9336
rect 14332 9324 14338 9376
rect 1104 9274 17756 9296
rect 1104 9222 7288 9274
rect 7340 9222 7352 9274
rect 7404 9222 7416 9274
rect 7468 9222 7480 9274
rect 7532 9222 13595 9274
rect 13647 9222 13659 9274
rect 13711 9222 13723 9274
rect 13775 9222 13787 9274
rect 13839 9222 17756 9274
rect 1104 9200 17756 9222
rect 1486 9120 1492 9172
rect 1544 9160 1550 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 1544 9132 1593 9160
rect 1544 9120 1550 9132
rect 1581 9129 1593 9132
rect 1627 9129 1639 9163
rect 1581 9123 1639 9129
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 2498 9160 2504 9172
rect 2087 9132 2504 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2056 9024 2084 9123
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 1443 8996 2084 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2498 8956 2504 8968
rect 2459 8928 2504 8956
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 16022 8956 16028 8968
rect 15983 8928 16028 8956
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 16298 8956 16304 8968
rect 16259 8928 16304 8956
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 15562 8888 15568 8900
rect 15475 8860 15568 8888
rect 15562 8848 15568 8860
rect 15620 8888 15626 8900
rect 16316 8888 16344 8916
rect 15620 8860 16344 8888
rect 15620 8848 15626 8860
rect 1104 8730 17756 8752
rect 1104 8678 4135 8730
rect 4187 8678 4199 8730
rect 4251 8678 4263 8730
rect 4315 8678 4327 8730
rect 4379 8678 10441 8730
rect 10493 8678 10505 8730
rect 10557 8678 10569 8730
rect 10621 8678 10633 8730
rect 10685 8678 16748 8730
rect 16800 8678 16812 8730
rect 16864 8678 16876 8730
rect 16928 8678 16940 8730
rect 16992 8678 17756 8730
rect 1104 8656 17756 8678
rect 12526 8576 12532 8628
rect 12584 8616 12590 8628
rect 12621 8619 12679 8625
rect 12621 8616 12633 8619
rect 12584 8588 12633 8616
rect 12584 8576 12590 8588
rect 12621 8585 12633 8588
rect 12667 8585 12679 8619
rect 16022 8616 16028 8628
rect 15983 8588 16028 8616
rect 12621 8579 12679 8585
rect 16022 8576 16028 8588
rect 16080 8616 16086 8628
rect 16439 8619 16497 8625
rect 16439 8616 16451 8619
rect 16080 8588 16451 8616
rect 16080 8576 16086 8588
rect 16439 8585 16451 8588
rect 16485 8585 16497 8619
rect 16439 8579 16497 8585
rect 16853 8619 16911 8625
rect 16853 8585 16865 8619
rect 16899 8616 16911 8619
rect 17034 8616 17040 8628
rect 16899 8588 17040 8616
rect 16899 8585 16911 8588
rect 16853 8579 16911 8585
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 1903 8452 2053 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 2041 8449 2053 8452
rect 2087 8480 2099 8483
rect 2498 8480 2504 8492
rect 2087 8452 2504 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2498 8440 2504 8452
rect 2556 8440 2562 8492
rect 2682 8480 2688 8492
rect 2643 8452 2688 8480
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 3580 8415 3638 8421
rect 3580 8381 3592 8415
rect 3626 8412 3638 8415
rect 3970 8412 3976 8424
rect 3626 8384 3976 8412
rect 3626 8381 3638 8384
rect 3580 8375 3638 8381
rect 3970 8372 3976 8384
rect 4028 8372 4034 8424
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 16368 8415 16426 8421
rect 12483 8384 13124 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 13096 8288 13124 8384
rect 16368 8381 16380 8415
rect 16414 8412 16426 8415
rect 16868 8412 16896 8579
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 16414 8384 16896 8412
rect 16414 8381 16426 8384
rect 16368 8375 16426 8381
rect 1762 8236 1768 8288
rect 1820 8276 1826 8288
rect 3651 8279 3709 8285
rect 3651 8276 3663 8279
rect 1820 8248 3663 8276
rect 1820 8236 1826 8248
rect 3651 8245 3663 8248
rect 3697 8245 3709 8279
rect 13078 8276 13084 8288
rect 13039 8248 13084 8276
rect 3651 8239 3709 8245
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 1104 8186 17756 8208
rect 1104 8134 7288 8186
rect 7340 8134 7352 8186
rect 7404 8134 7416 8186
rect 7468 8134 7480 8186
rect 7532 8134 13595 8186
rect 13647 8134 13659 8186
rect 13711 8134 13723 8186
rect 13775 8134 13787 8186
rect 13839 8134 17756 8186
rect 1104 8112 17756 8134
rect 1762 8072 1768 8084
rect 1723 8044 1768 8072
rect 1762 8032 1768 8044
rect 1820 8032 1826 8084
rect 13078 8032 13084 8084
rect 13136 8072 13142 8084
rect 13219 8075 13277 8081
rect 13219 8072 13231 8075
rect 13136 8044 13231 8072
rect 13136 8032 13142 8044
rect 13219 8041 13231 8044
rect 13265 8041 13277 8075
rect 13219 8035 13277 8041
rect 12894 7896 12900 7948
rect 12952 7936 12958 7948
rect 13116 7939 13174 7945
rect 13116 7936 13128 7939
rect 12952 7908 13128 7936
rect 12952 7896 12958 7908
rect 13116 7905 13128 7908
rect 13162 7905 13174 7939
rect 13116 7899 13174 7905
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 2682 7868 2688 7880
rect 2643 7840 2688 7868
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 12066 7868 12072 7880
rect 12027 7840 12072 7868
rect 12066 7828 12072 7840
rect 12124 7828 12130 7880
rect 16022 7868 16028 7880
rect 15983 7840 16028 7868
rect 16022 7828 16028 7840
rect 16080 7828 16086 7880
rect 16298 7868 16304 7880
rect 16259 7840 16304 7868
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 1104 7642 17756 7664
rect 1104 7590 4135 7642
rect 4187 7590 4199 7642
rect 4251 7590 4263 7642
rect 4315 7590 4327 7642
rect 4379 7590 10441 7642
rect 10493 7590 10505 7642
rect 10557 7590 10569 7642
rect 10621 7590 10633 7642
rect 10685 7590 16748 7642
rect 16800 7590 16812 7642
rect 16864 7590 16876 7642
rect 16928 7590 16940 7642
rect 16992 7590 17756 7642
rect 1104 7568 17756 7590
rect 12066 7488 12072 7540
rect 12124 7528 12130 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 12124 7500 12173 7528
rect 12124 7488 12130 7500
rect 12161 7497 12173 7500
rect 12207 7528 12219 7531
rect 14277 7531 14335 7537
rect 12207 7500 12572 7528
rect 12207 7497 12219 7500
rect 12161 7491 12219 7497
rect 1762 7392 1768 7404
rect 1723 7364 1768 7392
rect 1762 7352 1768 7364
rect 1820 7352 1826 7404
rect 2222 7352 2228 7404
rect 2280 7392 2286 7404
rect 12544 7401 12572 7500
rect 14277 7497 14289 7531
rect 14323 7528 14335 7531
rect 15194 7528 15200 7540
rect 14323 7500 15200 7528
rect 14323 7497 14335 7500
rect 14277 7491 14335 7497
rect 15194 7488 15200 7500
rect 15252 7488 15258 7540
rect 16022 7528 16028 7540
rect 15983 7500 16028 7528
rect 16022 7488 16028 7500
rect 16080 7528 16086 7540
rect 16439 7531 16497 7537
rect 16439 7528 16451 7531
rect 16080 7500 16451 7528
rect 16080 7488 16086 7500
rect 16439 7497 16451 7500
rect 16485 7497 16497 7531
rect 16439 7491 16497 7497
rect 2409 7395 2467 7401
rect 2409 7392 2421 7395
rect 2280 7364 2421 7392
rect 2280 7352 2286 7364
rect 2409 7361 2421 7364
rect 2455 7392 2467 7395
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 2455 7364 2789 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 2777 7361 2789 7364
rect 2823 7392 2835 7395
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 2823 7364 5549 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 5537 7361 5549 7364
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7361 12587 7395
rect 12894 7392 12900 7404
rect 12855 7364 12900 7392
rect 12529 7355 12587 7361
rect 12894 7352 12900 7364
rect 12952 7392 12958 7404
rect 13449 7395 13507 7401
rect 13449 7392 13461 7395
rect 12952 7364 13461 7392
rect 12952 7352 12958 7364
rect 13449 7361 13461 7364
rect 13495 7361 13507 7395
rect 13449 7355 13507 7361
rect 14090 7324 14096 7336
rect 14003 7296 14096 7324
rect 14090 7284 14096 7296
rect 14148 7324 14154 7336
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 14148 7296 14657 7324
rect 14148 7284 14154 7296
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 14645 7287 14703 7293
rect 16368 7327 16426 7333
rect 16368 7293 16380 7327
rect 16414 7324 16426 7327
rect 16414 7296 16896 7324
rect 16414 7293 16426 7296
rect 16368 7287 16426 7293
rect 5077 7259 5135 7265
rect 5077 7225 5089 7259
rect 5123 7256 5135 7259
rect 5258 7256 5264 7268
rect 5123 7228 5264 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 5258 7216 5264 7228
rect 5316 7216 5322 7268
rect 16868 7197 16896 7296
rect 16853 7191 16911 7197
rect 16853 7157 16865 7191
rect 16899 7188 16911 7191
rect 17862 7188 17868 7200
rect 16899 7160 17868 7188
rect 16899 7157 16911 7160
rect 16853 7151 16911 7157
rect 17862 7148 17868 7160
rect 17920 7148 17926 7200
rect 1104 7098 17756 7120
rect 1104 7046 7288 7098
rect 7340 7046 7352 7098
rect 7404 7046 7416 7098
rect 7468 7046 7480 7098
rect 7532 7046 13595 7098
rect 13647 7046 13659 7098
rect 13711 7046 13723 7098
rect 13775 7046 13787 7098
rect 13839 7046 17756 7098
rect 1104 7024 17756 7046
rect 5258 6944 5264 6996
rect 5316 6984 5322 6996
rect 5583 6987 5641 6993
rect 5583 6984 5595 6987
rect 5316 6956 5595 6984
rect 5316 6944 5322 6956
rect 5583 6953 5595 6956
rect 5629 6953 5641 6987
rect 5583 6947 5641 6953
rect 13863 6987 13921 6993
rect 13863 6953 13875 6987
rect 13909 6984 13921 6987
rect 14090 6984 14096 6996
rect 13909 6956 14096 6984
rect 13909 6953 13921 6956
rect 13863 6947 13921 6953
rect 14090 6944 14096 6956
rect 14148 6944 14154 6996
rect 12894 6916 12900 6928
rect 12855 6888 12900 6916
rect 12894 6876 12900 6888
rect 12952 6876 12958 6928
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6848 5503 6851
rect 5534 6848 5540 6860
rect 5491 6820 5540 6848
rect 5491 6817 5503 6820
rect 5445 6811 5503 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 13722 6848 13728 6860
rect 13683 6820 13728 6848
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 1854 6780 1860 6792
rect 1815 6752 1860 6780
rect 1854 6740 1860 6752
rect 1912 6740 1918 6792
rect 2314 6780 2320 6792
rect 2275 6752 2320 6780
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 11882 6740 11888 6792
rect 11940 6780 11946 6792
rect 12253 6783 12311 6789
rect 12253 6780 12265 6783
rect 11940 6752 12265 6780
rect 11940 6740 11946 6752
rect 12253 6749 12265 6752
rect 12299 6749 12311 6783
rect 12253 6743 12311 6749
rect 1104 6554 17756 6576
rect 1104 6502 4135 6554
rect 4187 6502 4199 6554
rect 4251 6502 4263 6554
rect 4315 6502 4327 6554
rect 4379 6502 10441 6554
rect 10493 6502 10505 6554
rect 10557 6502 10569 6554
rect 10621 6502 10633 6554
rect 10685 6502 16748 6554
rect 16800 6502 16812 6554
rect 16864 6502 16876 6554
rect 16928 6502 16940 6554
rect 16992 6502 17756 6554
rect 1104 6480 17756 6502
rect 13722 6372 13728 6384
rect 9324 6344 13728 6372
rect 9324 6316 9352 6344
rect 13722 6332 13728 6344
rect 13780 6332 13786 6384
rect 1535 6307 1593 6313
rect 1535 6273 1547 6307
rect 1581 6304 1593 6307
rect 1854 6304 1860 6316
rect 1581 6276 1860 6304
rect 1581 6273 1593 6276
rect 1535 6267 1593 6273
rect 1854 6264 1860 6276
rect 1912 6304 1918 6316
rect 2225 6307 2283 6313
rect 2225 6304 2237 6307
rect 1912 6276 2237 6304
rect 1912 6264 1918 6276
rect 2225 6273 2237 6276
rect 2271 6273 2283 6307
rect 9306 6304 9312 6316
rect 9267 6276 9312 6304
rect 2225 6267 2283 6273
rect 9306 6264 9312 6276
rect 9364 6264 9370 6316
rect 11882 6264 11888 6316
rect 11940 6304 11946 6316
rect 12805 6307 12863 6313
rect 12805 6304 12817 6307
rect 11940 6276 12817 6304
rect 11940 6264 11946 6276
rect 12805 6273 12817 6276
rect 12851 6273 12863 6307
rect 12805 6267 12863 6273
rect 1448 6239 1506 6245
rect 1448 6205 1460 6239
rect 1494 6236 1506 6239
rect 1494 6208 1716 6236
rect 1494 6205 1506 6208
rect 1448 6199 1506 6205
rect 1688 6180 1716 6208
rect 1670 6128 1676 6180
rect 1728 6168 1734 6180
rect 1857 6171 1915 6177
rect 1857 6168 1869 6171
rect 1728 6140 1869 6168
rect 1728 6128 1734 6140
rect 1857 6137 1869 6140
rect 1903 6137 1915 6171
rect 9033 6171 9091 6177
rect 9033 6168 9045 6171
rect 1857 6131 1915 6137
rect 8772 6140 9045 6168
rect 5534 6100 5540 6112
rect 5447 6072 5540 6100
rect 5534 6060 5540 6072
rect 5592 6100 5598 6112
rect 6454 6100 6460 6112
rect 5592 6072 6460 6100
rect 5592 6060 5598 6072
rect 6454 6060 6460 6072
rect 6512 6060 6518 6112
rect 8772 6109 8800 6140
rect 9033 6137 9045 6140
rect 9079 6137 9091 6171
rect 9033 6131 9091 6137
rect 12253 6171 12311 6177
rect 12253 6137 12265 6171
rect 12299 6168 12311 6171
rect 12526 6168 12532 6180
rect 12299 6140 12532 6168
rect 12299 6137 12311 6140
rect 12253 6131 12311 6137
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 7929 6103 7987 6109
rect 7929 6069 7941 6103
rect 7975 6100 7987 6103
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 7975 6072 8769 6100
rect 7975 6069 7987 6072
rect 7929 6063 7987 6069
rect 8757 6069 8769 6072
rect 8803 6069 8815 6103
rect 11882 6100 11888 6112
rect 11843 6072 11888 6100
rect 8757 6063 8815 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 1104 6010 17756 6032
rect 1104 5958 7288 6010
rect 7340 5958 7352 6010
rect 7404 5958 7416 6010
rect 7468 5958 7480 6010
rect 7532 5958 13595 6010
rect 13647 5958 13659 6010
rect 13711 5958 13723 6010
rect 13775 5958 13787 6010
rect 13839 5958 17756 6010
rect 1104 5936 17756 5958
rect 12526 5856 12532 5908
rect 12584 5896 12590 5908
rect 13035 5899 13093 5905
rect 13035 5896 13047 5899
rect 12584 5868 13047 5896
rect 12584 5856 12590 5868
rect 13035 5865 13047 5868
rect 13081 5865 13093 5899
rect 13035 5859 13093 5865
rect 8757 5831 8815 5837
rect 8757 5797 8769 5831
rect 8803 5828 8815 5831
rect 9306 5828 9312 5840
rect 8803 5800 9312 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 6270 5760 6276 5772
rect 6231 5732 6276 5760
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 12897 5763 12955 5769
rect 12897 5729 12909 5763
rect 12943 5760 12955 5763
rect 12986 5760 12992 5772
rect 12943 5732 12992 5760
rect 12943 5729 12955 5732
rect 12897 5723 12955 5729
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 8110 5692 8116 5704
rect 8071 5664 8116 5692
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 10459 5695 10517 5701
rect 10459 5661 10471 5695
rect 10505 5692 10517 5695
rect 11422 5692 11428 5704
rect 10505 5664 11428 5692
rect 10505 5661 10517 5664
rect 10459 5655 10517 5661
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 11882 5692 11888 5704
rect 11843 5664 11888 5692
rect 11882 5652 11888 5664
rect 11940 5652 11946 5704
rect 6411 5559 6469 5565
rect 6411 5525 6423 5559
rect 6457 5556 6469 5559
rect 7006 5556 7012 5568
rect 6457 5528 7012 5556
rect 6457 5525 6469 5528
rect 6411 5519 6469 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 10226 5556 10232 5568
rect 10187 5528 10232 5556
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 1104 5466 17756 5488
rect 1104 5414 4135 5466
rect 4187 5414 4199 5466
rect 4251 5414 4263 5466
rect 4315 5414 4327 5466
rect 4379 5414 10441 5466
rect 10493 5414 10505 5466
rect 10557 5414 10569 5466
rect 10621 5414 10633 5466
rect 10685 5414 16748 5466
rect 16800 5414 16812 5466
rect 16864 5414 16876 5466
rect 16928 5414 16940 5466
rect 16992 5414 17756 5466
rect 1104 5392 17756 5414
rect 106 5312 112 5364
rect 164 5352 170 5364
rect 6270 5352 6276 5364
rect 164 5324 6276 5352
rect 164 5312 170 5324
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 7006 5352 7012 5364
rect 6967 5324 7012 5352
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 8168 5324 8217 5352
rect 8168 5312 8174 5324
rect 8205 5321 8217 5324
rect 8251 5321 8263 5355
rect 8205 5315 8263 5321
rect 9490 5312 9496 5364
rect 9548 5352 9554 5364
rect 9585 5355 9643 5361
rect 9585 5352 9597 5355
rect 9548 5324 9597 5352
rect 9548 5312 9554 5324
rect 9585 5321 9597 5324
rect 9631 5321 9643 5355
rect 11422 5352 11428 5364
rect 11383 5324 11428 5352
rect 9585 5315 9643 5321
rect 11422 5312 11428 5324
rect 11480 5312 11486 5364
rect 12986 5352 12992 5364
rect 12947 5324 12992 5352
rect 12986 5312 12992 5324
rect 13044 5312 13050 5364
rect 7024 5216 7052 5312
rect 7837 5287 7895 5293
rect 7837 5253 7849 5287
rect 7883 5284 7895 5287
rect 8128 5284 8156 5312
rect 7883 5256 8156 5284
rect 7883 5253 7895 5256
rect 7837 5247 7895 5253
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 7024 5188 7297 5216
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5148 9459 5151
rect 10556 5151 10614 5157
rect 9447 5120 10088 5148
rect 9447 5117 9459 5120
rect 9401 5111 9459 5117
rect 10060 5089 10088 5120
rect 10556 5117 10568 5151
rect 10602 5148 10614 5151
rect 10602 5120 11100 5148
rect 10602 5117 10614 5120
rect 10556 5111 10614 5117
rect 10045 5083 10103 5089
rect 10045 5049 10057 5083
rect 10091 5080 10103 5083
rect 10643 5083 10701 5089
rect 10643 5080 10655 5083
rect 10091 5052 10655 5080
rect 10091 5049 10103 5052
rect 10045 5043 10103 5049
rect 10643 5049 10655 5052
rect 10689 5049 10701 5083
rect 10643 5043 10701 5049
rect 6362 4972 6368 5024
rect 6420 5012 6426 5024
rect 10226 5012 10232 5024
rect 6420 4984 10232 5012
rect 6420 4972 6426 4984
rect 10226 4972 10232 4984
rect 10284 5012 10290 5024
rect 11072 5021 11100 5120
rect 10321 5015 10379 5021
rect 10321 5012 10333 5015
rect 10284 4984 10333 5012
rect 10284 4972 10290 4984
rect 10321 4981 10333 4984
rect 10367 4981 10379 5015
rect 10321 4975 10379 4981
rect 11057 5015 11115 5021
rect 11057 4981 11069 5015
rect 11103 5012 11115 5015
rect 11606 5012 11612 5024
rect 11103 4984 11612 5012
rect 11103 4981 11115 4984
rect 11057 4975 11115 4981
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 1104 4922 17756 4944
rect 1104 4870 7288 4922
rect 7340 4870 7352 4922
rect 7404 4870 7416 4922
rect 7468 4870 7480 4922
rect 7532 4870 13595 4922
rect 13647 4870 13659 4922
rect 13711 4870 13723 4922
rect 13775 4870 13787 4922
rect 13839 4870 17756 4922
rect 1104 4848 17756 4870
rect 7745 4743 7803 4749
rect 7745 4709 7757 4743
rect 7791 4740 7803 4743
rect 8018 4740 8024 4752
rect 7791 4712 8024 4740
rect 7791 4709 7803 4712
rect 7745 4703 7803 4709
rect 8018 4700 8024 4712
rect 8076 4700 8082 4752
rect 8110 4700 8116 4752
rect 8168 4740 8174 4752
rect 8389 4743 8447 4749
rect 8389 4740 8401 4743
rect 8168 4712 8401 4740
rect 8168 4700 8174 4712
rect 8389 4709 8401 4712
rect 8435 4709 8447 4743
rect 8389 4703 8447 4709
rect 12504 4675 12562 4681
rect 12504 4641 12516 4675
rect 12550 4672 12562 4675
rect 13262 4672 13268 4684
rect 12550 4644 13268 4672
rect 12550 4641 12562 4644
rect 12504 4635 12562 4641
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 9674 4604 9680 4616
rect 9635 4576 9680 4604
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 10689 4607 10747 4613
rect 10689 4573 10701 4607
rect 10735 4604 10747 4607
rect 10778 4604 10784 4616
rect 10735 4576 10784 4604
rect 10735 4573 10747 4576
rect 10689 4567 10747 4573
rect 10778 4564 10784 4576
rect 10836 4564 10842 4616
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 12342 4428 12348 4480
rect 12400 4468 12406 4480
rect 12575 4471 12633 4477
rect 12575 4468 12587 4471
rect 12400 4440 12587 4468
rect 12400 4428 12406 4440
rect 12575 4437 12587 4440
rect 12621 4437 12633 4471
rect 12575 4431 12633 4437
rect 1104 4378 17756 4400
rect 1104 4326 4135 4378
rect 4187 4326 4199 4378
rect 4251 4326 4263 4378
rect 4315 4326 4327 4378
rect 4379 4326 10441 4378
rect 10493 4326 10505 4378
rect 10557 4326 10569 4378
rect 10621 4326 10633 4378
rect 10685 4326 16748 4378
rect 16800 4326 16812 4378
rect 16864 4326 16876 4378
rect 16928 4326 16940 4378
rect 16992 4326 17756 4378
rect 1104 4304 17756 4326
rect 7650 4264 7656 4276
rect 7611 4236 7656 4264
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 9674 4196 9680 4208
rect 8680 4168 9680 4196
rect 1489 4131 1547 4137
rect 1489 4097 1501 4131
rect 1535 4128 1547 4131
rect 1578 4128 1584 4140
rect 1535 4100 1584 4128
rect 1535 4097 1547 4100
rect 1489 4091 1547 4097
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 2130 4128 2136 4140
rect 2091 4100 2136 4128
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 8680 4137 8708 4168
rect 9674 4156 9680 4168
rect 9732 4156 9738 4208
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 8527 4100 8677 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8665 4097 8677 4100
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 10689 4131 10747 4137
rect 10689 4128 10701 4131
rect 10551 4100 10701 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 10689 4097 10701 4100
rect 10735 4128 10747 4131
rect 10778 4128 10784 4140
rect 10735 4100 10784 4128
rect 10735 4097 10747 4100
rect 10689 4091 10747 4097
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 14918 4069 14924 4072
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4029 7527 4063
rect 14896 4063 14924 4069
rect 14896 4060 14908 4063
rect 14831 4032 14908 4060
rect 7469 4023 7527 4029
rect 14896 4029 14908 4032
rect 14976 4060 14982 4072
rect 15289 4063 15347 4069
rect 15289 4060 15301 4063
rect 14976 4032 15301 4060
rect 14896 4023 14924 4029
rect 7377 3927 7435 3933
rect 7377 3893 7389 3927
rect 7423 3924 7435 3927
rect 7484 3924 7512 4023
rect 14918 4020 14924 4023
rect 14976 4020 14982 4032
rect 15289 4029 15301 4032
rect 15335 4029 15347 4063
rect 15289 4023 15347 4029
rect 15908 4063 15966 4069
rect 15908 4029 15920 4063
rect 15954 4060 15966 4063
rect 15954 4032 16436 4060
rect 15954 4029 15966 4032
rect 15908 4023 15966 4029
rect 9306 3992 9312 4004
rect 9267 3964 9312 3992
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 11333 3995 11391 4001
rect 11333 3961 11345 3995
rect 11379 3992 11391 3995
rect 11606 3992 11612 4004
rect 11379 3964 11612 3992
rect 11379 3961 11391 3964
rect 11333 3955 11391 3961
rect 11606 3952 11612 3964
rect 11664 3952 11670 4004
rect 7650 3924 7656 3936
rect 7423 3896 7656 3924
rect 7423 3893 7435 3896
rect 7377 3887 7435 3893
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 8018 3924 8024 3936
rect 7979 3896 8024 3924
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 12434 3924 12440 3936
rect 12395 3896 12440 3924
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12989 3927 13047 3933
rect 12989 3893 13001 3927
rect 13035 3924 13047 3927
rect 13262 3924 13268 3936
rect 13035 3896 13268 3924
rect 13035 3893 13047 3896
rect 12989 3887 13047 3893
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 14967 3927 15025 3933
rect 14967 3893 14979 3927
rect 15013 3924 15025 3927
rect 15378 3924 15384 3936
rect 15013 3896 15384 3924
rect 15013 3893 15025 3896
rect 14967 3887 15025 3893
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 15654 3884 15660 3936
rect 15712 3924 15718 3936
rect 16408 3933 16436 4032
rect 15979 3927 16037 3933
rect 15979 3924 15991 3927
rect 15712 3896 15991 3924
rect 15712 3884 15718 3896
rect 15979 3893 15991 3896
rect 16025 3893 16037 3927
rect 15979 3887 16037 3893
rect 16393 3927 16451 3933
rect 16393 3893 16405 3927
rect 16439 3924 16451 3927
rect 16574 3924 16580 3936
rect 16439 3896 16580 3924
rect 16439 3893 16451 3896
rect 16393 3887 16451 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 1104 3834 17756 3856
rect 1104 3782 7288 3834
rect 7340 3782 7352 3834
rect 7404 3782 7416 3834
rect 7468 3782 7480 3834
rect 7532 3782 13595 3834
rect 13647 3782 13659 3834
rect 13711 3782 13723 3834
rect 13775 3782 13787 3834
rect 13839 3782 17756 3834
rect 1104 3760 17756 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 7239 3723 7297 3729
rect 7239 3689 7251 3723
rect 7285 3720 7297 3723
rect 8018 3720 8024 3732
rect 7285 3692 8024 3720
rect 7285 3689 7297 3692
rect 7239 3683 7297 3689
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 8251 3655 8309 3661
rect 8251 3652 8263 3655
rect 7708 3624 8263 3652
rect 7708 3612 7714 3624
rect 8251 3621 8263 3624
rect 8297 3621 8309 3655
rect 8251 3615 8309 3621
rect 9306 3612 9312 3664
rect 9364 3652 9370 3664
rect 10413 3655 10471 3661
rect 10413 3652 10425 3655
rect 9364 3624 10425 3652
rect 9364 3612 9370 3624
rect 10413 3621 10425 3624
rect 10459 3621 10471 3655
rect 15378 3652 15384 3664
rect 15339 3624 15384 3652
rect 10413 3615 10471 3621
rect 15378 3612 15384 3624
rect 15436 3612 15442 3664
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 8018 3544 8024 3596
rect 8076 3584 8082 3596
rect 8164 3587 8222 3593
rect 8164 3584 8176 3587
rect 8076 3556 8176 3584
rect 8076 3544 8082 3556
rect 8164 3553 8176 3556
rect 8210 3584 8222 3587
rect 9324 3584 9352 3612
rect 8210 3556 9352 3584
rect 13792 3587 13850 3593
rect 8210 3553 8222 3556
rect 8164 3547 8222 3553
rect 13792 3553 13804 3587
rect 13838 3584 13850 3587
rect 13906 3584 13912 3596
rect 13838 3556 13912 3584
rect 13838 3553 13850 3556
rect 13792 3547 13850 3553
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 7006 3516 7012 3528
rect 6967 3488 7012 3516
rect 7006 3476 7012 3488
rect 7064 3476 7070 3528
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9769 3519 9827 3525
rect 9769 3516 9781 3519
rect 9088 3488 9781 3516
rect 9088 3476 9094 3488
rect 9769 3485 9781 3488
rect 9815 3516 9827 3519
rect 10870 3516 10876 3528
rect 9815 3488 10876 3516
rect 9815 3485 9827 3488
rect 9769 3479 9827 3485
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 11330 3516 11336 3528
rect 11291 3488 11336 3516
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 11606 3516 11612 3528
rect 11567 3488 11612 3516
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 15746 3516 15752 3528
rect 15707 3488 15752 3516
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 13863 3383 13921 3389
rect 13863 3349 13875 3383
rect 13909 3380 13921 3383
rect 14182 3380 14188 3392
rect 13909 3352 14188 3380
rect 13909 3349 13921 3352
rect 13863 3343 13921 3349
rect 14182 3340 14188 3352
rect 14240 3340 14246 3392
rect 1104 3290 17756 3312
rect 1104 3238 4135 3290
rect 4187 3238 4199 3290
rect 4251 3238 4263 3290
rect 4315 3238 4327 3290
rect 4379 3238 10441 3290
rect 10493 3238 10505 3290
rect 10557 3238 10569 3290
rect 10621 3238 10633 3290
rect 10685 3238 16748 3290
rect 16800 3238 16812 3290
rect 16864 3238 16876 3290
rect 16928 3238 16940 3290
rect 16992 3238 17756 3290
rect 1104 3216 17756 3238
rect 106 3136 112 3188
rect 164 3176 170 3188
rect 1394 3176 1400 3188
rect 164 3148 1400 3176
rect 164 3136 170 3148
rect 1394 3136 1400 3148
rect 1452 3176 1458 3188
rect 1581 3179 1639 3185
rect 1581 3176 1593 3179
rect 1452 3148 1593 3176
rect 1452 3136 1458 3148
rect 1581 3145 1593 3148
rect 1627 3145 1639 3179
rect 8018 3176 8024 3188
rect 7979 3148 8024 3176
rect 1581 3139 1639 3145
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 9030 3176 9036 3188
rect 8991 3148 9036 3176
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 11330 3176 11336 3188
rect 11291 3148 11336 3176
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12434 3176 12440 3188
rect 12299 3148 12440 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 15378 3176 15384 3188
rect 15339 3148 15384 3176
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 15746 3136 15752 3188
rect 15804 3176 15810 3188
rect 16669 3179 16727 3185
rect 16669 3176 16681 3179
rect 15804 3148 16681 3176
rect 15804 3136 15810 3148
rect 16669 3145 16681 3148
rect 16715 3145 16727 3179
rect 16669 3139 16727 3145
rect 8665 3111 8723 3117
rect 8665 3077 8677 3111
rect 8711 3108 8723 3111
rect 8711 3080 12388 3108
rect 8711 3077 8723 3080
rect 8665 3071 8723 3077
rect 8180 2975 8238 2981
rect 8180 2941 8192 2975
rect 8226 2972 8238 2975
rect 8680 2972 8708 3071
rect 8226 2944 8708 2972
rect 9176 2975 9234 2981
rect 8226 2941 8238 2944
rect 8180 2935 8238 2941
rect 9176 2941 9188 2975
rect 9222 2972 9234 2975
rect 9222 2941 9235 2972
rect 9176 2935 9235 2941
rect 7006 2796 7012 2848
rect 7064 2836 7070 2848
rect 7193 2839 7251 2845
rect 7193 2836 7205 2839
rect 7064 2808 7205 2836
rect 7064 2796 7070 2808
rect 7193 2805 7205 2808
rect 7239 2836 7251 2839
rect 7742 2836 7748 2848
rect 7239 2808 7748 2836
rect 7239 2805 7251 2808
rect 7193 2799 7251 2805
rect 7742 2796 7748 2808
rect 7800 2796 7806 2848
rect 8251 2839 8309 2845
rect 8251 2805 8263 2839
rect 8297 2836 8309 2839
rect 8478 2836 8484 2848
rect 8297 2808 8484 2836
rect 8297 2805 8309 2808
rect 8251 2799 8309 2805
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 9207 2836 9235 2935
rect 9263 2907 9321 2913
rect 9263 2873 9275 2907
rect 9309 2904 9321 2907
rect 9953 2907 10011 2913
rect 9953 2904 9965 2907
rect 9309 2876 9965 2904
rect 9309 2873 9321 2876
rect 9263 2867 9321 2873
rect 9953 2873 9965 2876
rect 9999 2904 10011 2907
rect 10229 2907 10287 2913
rect 10229 2904 10241 2907
rect 9999 2876 10241 2904
rect 9999 2873 10011 2876
rect 9953 2867 10011 2873
rect 10229 2873 10241 2876
rect 10275 2873 10287 2907
rect 10870 2904 10876 2916
rect 10831 2876 10876 2904
rect 10229 2867 10287 2873
rect 10870 2864 10876 2876
rect 10928 2864 10934 2916
rect 12360 2904 12388 3080
rect 12452 3040 12480 3136
rect 12621 3043 12679 3049
rect 12621 3040 12633 3043
rect 12452 3012 12633 3040
rect 12621 3009 12633 3012
rect 12667 3009 12679 3043
rect 14182 3040 14188 3052
rect 14143 3012 14188 3040
rect 12621 3003 12679 3009
rect 14182 3000 14188 3012
rect 14240 3000 14246 3052
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3040 14887 3043
rect 15746 3040 15752 3052
rect 14875 3012 15752 3040
rect 14875 3009 14887 3012
rect 14829 3003 14887 3009
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 13265 2907 13323 2913
rect 13265 2904 13277 2907
rect 12360 2876 13277 2904
rect 13265 2873 13277 2876
rect 13311 2904 13323 2907
rect 16393 2907 16451 2913
rect 16393 2904 16405 2907
rect 13311 2876 16405 2904
rect 13311 2873 13323 2876
rect 13265 2867 13323 2873
rect 16393 2873 16405 2876
rect 16439 2873 16451 2907
rect 16393 2867 16451 2873
rect 9677 2839 9735 2845
rect 9677 2836 9689 2839
rect 9207 2808 9689 2836
rect 9677 2805 9689 2808
rect 9723 2836 9735 2839
rect 10318 2836 10324 2848
rect 9723 2808 10324 2836
rect 9723 2805 9735 2808
rect 9677 2799 9735 2805
rect 10318 2796 10324 2808
rect 10376 2796 10382 2848
rect 13817 2839 13875 2845
rect 13817 2805 13829 2839
rect 13863 2836 13875 2839
rect 13906 2836 13912 2848
rect 13863 2808 13912 2836
rect 13863 2805 13875 2808
rect 13817 2799 13875 2805
rect 13906 2796 13912 2808
rect 13964 2836 13970 2848
rect 14550 2836 14556 2848
rect 13964 2808 14556 2836
rect 13964 2796 13970 2808
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 1104 2746 17756 2768
rect 1104 2694 7288 2746
rect 7340 2694 7352 2746
rect 7404 2694 7416 2746
rect 7468 2694 7480 2746
rect 7532 2694 13595 2746
rect 13647 2694 13659 2746
rect 13711 2694 13723 2746
rect 13775 2694 13787 2746
rect 13839 2694 17756 2746
rect 1104 2672 17756 2694
rect 12342 2632 12348 2644
rect 12303 2604 12348 2632
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 14182 2632 14188 2644
rect 14143 2604 14188 2632
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 10870 2524 10876 2576
rect 10928 2564 10934 2576
rect 11425 2567 11483 2573
rect 11425 2564 11437 2567
rect 10928 2536 11437 2564
rect 10928 2524 10934 2536
rect 11425 2533 11437 2536
rect 11471 2533 11483 2567
rect 12360 2564 12388 2592
rect 12805 2567 12863 2573
rect 12805 2564 12817 2567
rect 12360 2536 12817 2564
rect 11425 2527 11483 2533
rect 12805 2533 12817 2536
rect 12851 2533 12863 2567
rect 12805 2527 12863 2533
rect 13446 2524 13452 2576
rect 13504 2564 13510 2576
rect 16301 2567 16359 2573
rect 16301 2564 16313 2567
rect 13504 2536 16313 2564
rect 13504 2524 13510 2536
rect 16301 2533 16313 2536
rect 16347 2533 16359 2567
rect 16301 2527 16359 2533
rect 8478 2456 8484 2508
rect 8536 2496 8542 2508
rect 8573 2499 8631 2505
rect 8573 2496 8585 2499
rect 8536 2468 8585 2496
rect 8536 2456 8542 2468
rect 8573 2465 8585 2468
rect 8619 2496 8631 2499
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8619 2468 9137 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9125 2459 9183 2465
rect 14420 2499 14478 2505
rect 14420 2465 14432 2499
rect 14466 2496 14478 2499
rect 14466 2468 14964 2496
rect 14466 2465 14478 2468
rect 14420 2459 14478 2465
rect 10597 2431 10655 2437
rect 10597 2397 10609 2431
rect 10643 2428 10655 2431
rect 10781 2431 10839 2437
rect 10781 2428 10793 2431
rect 10643 2400 10793 2428
rect 10643 2397 10655 2400
rect 10597 2391 10655 2397
rect 10781 2397 10793 2400
rect 10827 2428 10839 2431
rect 14507 2431 14565 2437
rect 14507 2428 14519 2431
rect 10827 2400 14519 2428
rect 10827 2397 10839 2400
rect 10781 2391 10839 2397
rect 14507 2397 14519 2400
rect 14553 2397 14565 2431
rect 14507 2391 14565 2397
rect 8757 2363 8815 2369
rect 8757 2329 8769 2363
rect 8803 2360 8815 2363
rect 9490 2360 9496 2372
rect 8803 2332 9496 2360
rect 8803 2329 8815 2332
rect 8757 2323 8815 2329
rect 9490 2320 9496 2332
rect 9548 2320 9554 2372
rect 11422 2320 11428 2372
rect 11480 2360 11486 2372
rect 13357 2363 13415 2369
rect 13357 2360 13369 2363
rect 11480 2332 13369 2360
rect 11480 2320 11486 2332
rect 13357 2329 13369 2332
rect 13403 2360 13415 2363
rect 13446 2360 13452 2372
rect 13403 2332 13452 2360
rect 13403 2329 13415 2332
rect 13357 2323 13415 2329
rect 13446 2320 13452 2332
rect 13504 2320 13510 2372
rect 14936 2369 14964 2468
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15654 2428 15660 2440
rect 15335 2400 15660 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15654 2388 15660 2400
rect 15712 2388 15718 2440
rect 14921 2363 14979 2369
rect 14921 2329 14933 2363
rect 14967 2360 14979 2363
rect 15378 2360 15384 2372
rect 14967 2332 15384 2360
rect 14967 2329 14979 2332
rect 14921 2323 14979 2329
rect 15378 2320 15384 2332
rect 15436 2320 15442 2372
rect 1104 2202 17756 2224
rect 1104 2150 4135 2202
rect 4187 2150 4199 2202
rect 4251 2150 4263 2202
rect 4315 2150 4327 2202
rect 4379 2150 10441 2202
rect 10493 2150 10505 2202
rect 10557 2150 10569 2202
rect 10621 2150 10633 2202
rect 10685 2150 16748 2202
rect 16800 2150 16812 2202
rect 16864 2150 16876 2202
rect 16928 2150 16940 2202
rect 16992 2150 17756 2202
rect 1104 2128 17756 2150
rect 11054 76 11060 128
rect 11112 116 11118 128
rect 11882 116 11888 128
rect 11112 88 11888 116
rect 11112 76 11118 88
rect 11882 76 11888 88
rect 11940 76 11946 128
<< via1 >>
rect 12532 20544 12584 20596
rect 13360 20544 13412 20596
rect 15292 19660 15344 19712
rect 16396 19660 16448 19712
rect 4135 18470 4187 18522
rect 4199 18470 4251 18522
rect 4263 18470 4315 18522
rect 4327 18470 4379 18522
rect 10441 18470 10493 18522
rect 10505 18470 10557 18522
rect 10569 18470 10621 18522
rect 10633 18470 10685 18522
rect 16748 18470 16800 18522
rect 16812 18470 16864 18522
rect 16876 18470 16928 18522
rect 16940 18470 16992 18522
rect 11428 18411 11480 18420
rect 11428 18377 11437 18411
rect 11437 18377 11471 18411
rect 11471 18377 11480 18411
rect 11428 18368 11480 18377
rect 2136 18164 2188 18216
rect 2688 18164 2740 18216
rect 4896 18164 4948 18216
rect 8484 18207 8536 18216
rect 8484 18173 8493 18207
rect 8493 18173 8527 18207
rect 8527 18173 8536 18207
rect 8484 18164 8536 18173
rect 11428 18164 11480 18216
rect 11612 18164 11664 18216
rect 8576 18096 8628 18148
rect 8668 18096 8720 18148
rect 18420 18096 18472 18148
rect 1400 18028 1452 18080
rect 2044 18028 2096 18080
rect 3976 18028 4028 18080
rect 5080 18028 5132 18080
rect 7932 18028 7984 18080
rect 9956 18071 10008 18080
rect 9956 18037 9965 18071
rect 9965 18037 9999 18071
rect 9999 18037 10008 18071
rect 9956 18028 10008 18037
rect 11520 18028 11572 18080
rect 14188 18028 14240 18080
rect 7288 17926 7340 17978
rect 7352 17926 7404 17978
rect 7416 17926 7468 17978
rect 7480 17926 7532 17978
rect 13595 17926 13647 17978
rect 13659 17926 13711 17978
rect 13723 17926 13775 17978
rect 13787 17926 13839 17978
rect 20 17824 72 17876
rect 6092 17824 6144 17876
rect 8116 17867 8168 17876
rect 8116 17833 8125 17867
rect 8125 17833 8159 17867
rect 8159 17833 8168 17867
rect 8116 17824 8168 17833
rect 10232 17867 10284 17876
rect 10232 17833 10241 17867
rect 10241 17833 10275 17867
rect 10275 17833 10284 17867
rect 10232 17824 10284 17833
rect 14372 17824 14424 17876
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 3240 17756 3292 17808
rect 4436 17756 4488 17808
rect 4896 17799 4948 17808
rect 4896 17765 4905 17799
rect 4905 17765 4939 17799
rect 4939 17765 4948 17799
rect 4896 17756 4948 17765
rect 11520 17799 11572 17808
rect 11520 17765 11529 17799
rect 11529 17765 11563 17799
rect 11563 17765 11572 17799
rect 11520 17756 11572 17765
rect 7932 17731 7984 17740
rect 7932 17697 7941 17731
rect 7941 17697 7975 17731
rect 7975 17697 7984 17731
rect 7932 17688 7984 17697
rect 10048 17731 10100 17740
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 12900 17688 12952 17740
rect 16304 17688 16356 17740
rect 6644 17620 6696 17672
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 15384 17663 15436 17672
rect 15384 17629 15393 17663
rect 15393 17629 15427 17663
rect 15427 17629 15436 17663
rect 15384 17620 15436 17629
rect 4436 17552 4488 17604
rect 112 17484 164 17536
rect 3884 17484 3936 17536
rect 16212 17484 16264 17536
rect 4135 17382 4187 17434
rect 4199 17382 4251 17434
rect 4263 17382 4315 17434
rect 4327 17382 4379 17434
rect 10441 17382 10493 17434
rect 10505 17382 10557 17434
rect 10569 17382 10621 17434
rect 10633 17382 10685 17434
rect 16748 17382 16800 17434
rect 16812 17382 16864 17434
rect 16876 17382 16928 17434
rect 16940 17382 16992 17434
rect 1400 17280 1452 17332
rect 3240 17323 3292 17332
rect 3240 17289 3249 17323
rect 3249 17289 3283 17323
rect 3283 17289 3292 17323
rect 3240 17280 3292 17289
rect 3976 17323 4028 17332
rect 3976 17289 3985 17323
rect 3985 17289 4019 17323
rect 4019 17289 4028 17323
rect 3976 17280 4028 17289
rect 7932 17280 7984 17332
rect 8576 17323 8628 17332
rect 8576 17289 8585 17323
rect 8585 17289 8619 17323
rect 8619 17289 8628 17323
rect 8576 17280 8628 17289
rect 9956 17280 10008 17332
rect 11520 17323 11572 17332
rect 4896 17144 4948 17196
rect 8484 17144 8536 17196
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 14188 17280 14240 17332
rect 16212 17323 16264 17332
rect 12164 17144 12216 17196
rect 16212 17289 16221 17323
rect 16221 17289 16255 17323
rect 16255 17289 16264 17323
rect 16212 17280 16264 17289
rect 17408 17280 17460 17332
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 6092 17076 6144 17128
rect 16212 17076 16264 17128
rect 2320 17008 2372 17060
rect 8208 17008 8260 17060
rect 8576 17008 8628 17060
rect 11888 17008 11940 17060
rect 13176 17051 13228 17060
rect 13176 17017 13185 17051
rect 13185 17017 13219 17051
rect 13219 17017 13228 17051
rect 13176 17008 13228 17017
rect 4436 16940 4488 16992
rect 6644 16983 6696 16992
rect 6644 16949 6653 16983
rect 6653 16949 6687 16983
rect 6687 16949 6696 16983
rect 6644 16940 6696 16949
rect 10048 16983 10100 16992
rect 10048 16949 10057 16983
rect 10057 16949 10091 16983
rect 10091 16949 10100 16983
rect 10048 16940 10100 16949
rect 10784 16940 10836 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 16304 16940 16356 16992
rect 7288 16838 7340 16890
rect 7352 16838 7404 16890
rect 7416 16838 7468 16890
rect 7480 16838 7532 16890
rect 13595 16838 13647 16890
rect 13659 16838 13711 16890
rect 13723 16838 13775 16890
rect 13787 16838 13839 16890
rect 4436 16736 4488 16788
rect 5448 16736 5500 16788
rect 6184 16779 6236 16788
rect 6184 16745 6193 16779
rect 6193 16745 6227 16779
rect 6227 16745 6236 16779
rect 6184 16736 6236 16745
rect 12164 16736 12216 16788
rect 13176 16779 13228 16788
rect 13176 16745 13185 16779
rect 13185 16745 13219 16779
rect 13219 16745 13228 16779
rect 13176 16736 13228 16745
rect 2044 16668 2096 16720
rect 11612 16711 11664 16720
rect 11612 16677 11621 16711
rect 11621 16677 11655 16711
rect 11655 16677 11664 16711
rect 11612 16668 11664 16677
rect 5080 16600 5132 16652
rect 6000 16643 6052 16652
rect 6000 16609 6009 16643
rect 6009 16609 6043 16643
rect 6043 16609 6052 16643
rect 6000 16600 6052 16609
rect 13636 16643 13688 16652
rect 13636 16609 13654 16643
rect 13654 16609 13688 16643
rect 18328 16736 18380 16788
rect 15384 16668 15436 16720
rect 13636 16600 13688 16609
rect 2228 16575 2280 16584
rect 2228 16541 2237 16575
rect 2237 16541 2271 16575
rect 2271 16541 2280 16575
rect 2228 16532 2280 16541
rect 8208 16532 8260 16584
rect 8484 16575 8536 16584
rect 8484 16541 8493 16575
rect 8493 16541 8527 16575
rect 8527 16541 8536 16575
rect 8484 16532 8536 16541
rect 10048 16575 10100 16584
rect 10048 16541 10057 16575
rect 10057 16541 10091 16575
rect 10091 16541 10100 16575
rect 10048 16532 10100 16541
rect 10324 16575 10376 16584
rect 10324 16541 10333 16575
rect 10333 16541 10367 16575
rect 10367 16541 10376 16575
rect 10324 16532 10376 16541
rect 11888 16575 11940 16584
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 11888 16532 11940 16541
rect 16304 16507 16356 16516
rect 16304 16473 16313 16507
rect 16313 16473 16347 16507
rect 16347 16473 16356 16507
rect 16304 16464 16356 16473
rect 4135 16294 4187 16346
rect 4199 16294 4251 16346
rect 4263 16294 4315 16346
rect 4327 16294 4379 16346
rect 10441 16294 10493 16346
rect 10505 16294 10557 16346
rect 10569 16294 10621 16346
rect 10633 16294 10685 16346
rect 16748 16294 16800 16346
rect 16812 16294 16864 16346
rect 16876 16294 16928 16346
rect 16940 16294 16992 16346
rect 2044 16192 2096 16244
rect 3884 16235 3936 16244
rect 3884 16201 3893 16235
rect 3893 16201 3927 16235
rect 3927 16201 3936 16235
rect 5080 16235 5132 16244
rect 3884 16192 3936 16201
rect 2136 16099 2188 16108
rect 2136 16065 2145 16099
rect 2145 16065 2179 16099
rect 2179 16065 2188 16099
rect 2136 16056 2188 16065
rect 5080 16201 5089 16235
rect 5089 16201 5123 16235
rect 5123 16201 5132 16235
rect 5080 16192 5132 16201
rect 6000 16192 6052 16244
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 6552 16056 6604 16108
rect 10324 16056 10376 16108
rect 8208 15988 8260 16040
rect 8944 15988 8996 16040
rect 2228 15920 2280 15972
rect 6736 15920 6788 15972
rect 11888 16192 11940 16244
rect 12900 16192 12952 16244
rect 13636 16235 13688 16244
rect 13636 16201 13645 16235
rect 13645 16201 13679 16235
rect 13679 16201 13688 16235
rect 13636 16192 13688 16201
rect 15108 16235 15160 16244
rect 15108 16201 15117 16235
rect 15117 16201 15151 16235
rect 15151 16201 15160 16235
rect 15108 16192 15160 16201
rect 15384 16192 15436 16244
rect 11612 16167 11664 16176
rect 11612 16133 11621 16167
rect 11621 16133 11655 16167
rect 11655 16133 11664 16167
rect 11612 16124 11664 16133
rect 16304 16167 16356 16176
rect 16304 16133 16313 16167
rect 16313 16133 16347 16167
rect 16347 16133 16356 16167
rect 16304 16124 16356 16133
rect 16120 16056 16172 16108
rect 8116 15852 8168 15904
rect 8944 15895 8996 15904
rect 8944 15861 8953 15895
rect 8953 15861 8987 15895
rect 8987 15861 8996 15895
rect 8944 15852 8996 15861
rect 9588 15852 9640 15904
rect 10048 15852 10100 15904
rect 10784 15852 10836 15904
rect 7288 15750 7340 15802
rect 7352 15750 7404 15802
rect 7416 15750 7468 15802
rect 7480 15750 7532 15802
rect 13595 15750 13647 15802
rect 13659 15750 13711 15802
rect 13723 15750 13775 15802
rect 13787 15750 13839 15802
rect 2136 15580 2188 15632
rect 6184 15580 6236 15632
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 6552 15487 6604 15496
rect 6552 15453 6561 15487
rect 6561 15453 6595 15487
rect 6595 15453 6604 15487
rect 6552 15444 6604 15453
rect 8116 15580 8168 15632
rect 8208 15580 8260 15632
rect 10324 15444 10376 15496
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 4135 15206 4187 15258
rect 4199 15206 4251 15258
rect 4263 15206 4315 15258
rect 4327 15206 4379 15258
rect 10441 15206 10493 15258
rect 10505 15206 10557 15258
rect 10569 15206 10621 15258
rect 10633 15206 10685 15258
rect 16748 15206 16800 15258
rect 16812 15206 16864 15258
rect 16876 15206 16928 15258
rect 16940 15206 16992 15258
rect 1768 15147 1820 15156
rect 1768 15113 1777 15147
rect 1777 15113 1811 15147
rect 1811 15113 1820 15147
rect 1768 15104 1820 15113
rect 6184 15147 6236 15156
rect 6184 15113 6193 15147
rect 6193 15113 6227 15147
rect 6227 15113 6236 15147
rect 6184 15104 6236 15113
rect 8116 15104 8168 15156
rect 10324 15104 10376 15156
rect 15844 15147 15896 15156
rect 15844 15113 15853 15147
rect 15853 15113 15887 15147
rect 15887 15113 15896 15147
rect 15844 15104 15896 15113
rect 1676 14968 1728 15020
rect 4436 14968 4488 15020
rect 6736 14968 6788 15020
rect 9588 15011 9640 15020
rect 9588 14977 9597 15011
rect 9597 14977 9631 15011
rect 9631 14977 9640 15011
rect 9588 14968 9640 14977
rect 2596 14875 2648 14884
rect 2596 14841 2605 14875
rect 2605 14841 2639 14875
rect 2639 14841 2648 14875
rect 2596 14832 2648 14841
rect 3608 14875 3660 14884
rect 3608 14841 3617 14875
rect 3617 14841 3651 14875
rect 3651 14841 3660 14875
rect 3608 14832 3660 14841
rect 5172 14875 5224 14884
rect 5172 14841 5181 14875
rect 5181 14841 5215 14875
rect 5215 14841 5224 14875
rect 5172 14832 5224 14841
rect 11060 14807 11112 14816
rect 11060 14773 11069 14807
rect 11069 14773 11103 14807
rect 11103 14773 11112 14807
rect 11060 14764 11112 14773
rect 16488 14764 16540 14816
rect 7288 14662 7340 14714
rect 7352 14662 7404 14714
rect 7416 14662 7468 14714
rect 7480 14662 7532 14714
rect 13595 14662 13647 14714
rect 13659 14662 13711 14714
rect 13723 14662 13775 14714
rect 13787 14662 13839 14714
rect 2596 14603 2648 14612
rect 2596 14569 2605 14603
rect 2605 14569 2639 14603
rect 2639 14569 2648 14603
rect 2596 14560 2648 14569
rect 5172 14560 5224 14612
rect 6644 14560 6696 14612
rect 2228 14535 2280 14544
rect 2228 14501 2237 14535
rect 2237 14501 2271 14535
rect 2271 14501 2280 14535
rect 2228 14492 2280 14501
rect 5632 14467 5684 14476
rect 5632 14433 5641 14467
rect 5641 14433 5675 14467
rect 5675 14433 5684 14467
rect 5632 14424 5684 14433
rect 7104 14424 7156 14476
rect 12440 14424 12492 14476
rect 2228 14356 2280 14408
rect 3976 14356 4028 14408
rect 2596 14288 2648 14340
rect 4135 14118 4187 14170
rect 4199 14118 4251 14170
rect 4263 14118 4315 14170
rect 4327 14118 4379 14170
rect 10441 14118 10493 14170
rect 10505 14118 10557 14170
rect 10569 14118 10621 14170
rect 10633 14118 10685 14170
rect 16748 14118 16800 14170
rect 16812 14118 16864 14170
rect 16876 14118 16928 14170
rect 16940 14118 16992 14170
rect 3976 14016 4028 14068
rect 7104 14059 7156 14068
rect 7104 14025 7113 14059
rect 7113 14025 7147 14059
rect 7147 14025 7156 14059
rect 7104 14016 7156 14025
rect 112 13948 164 14000
rect 5632 13991 5684 14000
rect 5632 13957 5641 13991
rect 5641 13957 5675 13991
rect 5675 13957 5684 13991
rect 5632 13948 5684 13957
rect 1124 13812 1176 13864
rect 2688 13923 2740 13932
rect 2688 13889 2697 13923
rect 2697 13889 2731 13923
rect 2731 13889 2740 13923
rect 2688 13880 2740 13889
rect 2964 13923 3016 13932
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 1676 13812 1728 13864
rect 8668 13880 8720 13932
rect 4988 13812 5040 13864
rect 2320 13744 2372 13796
rect 2228 13719 2280 13728
rect 2228 13685 2237 13719
rect 2237 13685 2271 13719
rect 2271 13685 2280 13719
rect 2228 13676 2280 13685
rect 7288 13574 7340 13626
rect 7352 13574 7404 13626
rect 7416 13574 7468 13626
rect 7480 13574 7532 13626
rect 13595 13574 13647 13626
rect 13659 13574 13711 13626
rect 13723 13574 13775 13626
rect 13787 13574 13839 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 3608 13472 3660 13524
rect 2044 13336 2096 13388
rect 2964 13336 3016 13388
rect 3976 13336 4028 13388
rect 16212 13336 16264 13388
rect 2044 13175 2096 13184
rect 2044 13141 2053 13175
rect 2053 13141 2087 13175
rect 2087 13141 2096 13175
rect 2044 13132 2096 13141
rect 2504 13132 2556 13184
rect 16304 13132 16356 13184
rect 4135 13030 4187 13082
rect 4199 13030 4251 13082
rect 4263 13030 4315 13082
rect 4327 13030 4379 13082
rect 10441 13030 10493 13082
rect 10505 13030 10557 13082
rect 10569 13030 10621 13082
rect 10633 13030 10685 13082
rect 16748 13030 16800 13082
rect 16812 13030 16864 13082
rect 16876 13030 16928 13082
rect 16940 13030 16992 13082
rect 2228 12928 2280 12980
rect 16212 12928 16264 12980
rect 2964 12860 3016 12912
rect 18420 12860 18472 12912
rect 1860 12767 1912 12776
rect 1860 12733 1869 12767
rect 1869 12733 1903 12767
rect 1903 12733 1912 12767
rect 1860 12724 1912 12733
rect 13176 12724 13228 12776
rect 16304 12767 16356 12776
rect 16304 12733 16313 12767
rect 16313 12733 16347 12767
rect 16347 12733 16356 12767
rect 16304 12724 16356 12733
rect 2780 12588 2832 12640
rect 3976 12588 4028 12640
rect 5264 12631 5316 12640
rect 5264 12597 5273 12631
rect 5273 12597 5307 12631
rect 5307 12597 5316 12631
rect 5264 12588 5316 12597
rect 5724 12631 5776 12640
rect 5724 12597 5733 12631
rect 5733 12597 5767 12631
rect 5767 12597 5776 12631
rect 5724 12588 5776 12597
rect 15108 12588 15160 12640
rect 15292 12631 15344 12640
rect 15292 12597 15301 12631
rect 15301 12597 15335 12631
rect 15335 12597 15344 12631
rect 15292 12588 15344 12597
rect 7288 12486 7340 12538
rect 7352 12486 7404 12538
rect 7416 12486 7468 12538
rect 7480 12486 7532 12538
rect 13595 12486 13647 12538
rect 13659 12486 13711 12538
rect 13723 12486 13775 12538
rect 13787 12486 13839 12538
rect 2964 12384 3016 12436
rect 5724 12384 5776 12436
rect 2044 12316 2096 12368
rect 15108 12316 15160 12368
rect 2504 12248 2556 12300
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 6276 12248 6328 12300
rect 3884 12180 3936 12232
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 112 12112 164 12164
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 4135 11942 4187 11994
rect 4199 11942 4251 11994
rect 4263 11942 4315 11994
rect 4327 11942 4379 11994
rect 10441 11942 10493 11994
rect 10505 11942 10557 11994
rect 10569 11942 10621 11994
rect 10633 11942 10685 11994
rect 16748 11942 16800 11994
rect 16812 11942 16864 11994
rect 16876 11942 16928 11994
rect 16940 11942 16992 11994
rect 2504 11883 2556 11892
rect 2504 11849 2513 11883
rect 2513 11849 2547 11883
rect 2547 11849 2556 11883
rect 2504 11840 2556 11849
rect 6276 11840 6328 11892
rect 14188 11883 14240 11892
rect 14188 11849 14197 11883
rect 14197 11849 14231 11883
rect 14231 11849 14240 11883
rect 14188 11840 14240 11849
rect 15108 11883 15160 11892
rect 15108 11849 15117 11883
rect 15117 11849 15151 11883
rect 15151 11849 15160 11883
rect 15108 11840 15160 11849
rect 15292 11840 15344 11892
rect 1584 11704 1636 11756
rect 3884 11747 3936 11756
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 3976 11704 4028 11756
rect 16212 11747 16264 11756
rect 16212 11713 16221 11747
rect 16221 11713 16255 11747
rect 16255 11713 16264 11747
rect 16212 11704 16264 11713
rect 14648 11636 14700 11688
rect 2320 11568 2372 11620
rect 5080 11543 5132 11552
rect 5080 11509 5089 11543
rect 5089 11509 5123 11543
rect 5123 11509 5132 11543
rect 5080 11500 5132 11509
rect 7288 11398 7340 11450
rect 7352 11398 7404 11450
rect 7416 11398 7468 11450
rect 7480 11398 7532 11450
rect 13595 11398 13647 11450
rect 13659 11398 13711 11450
rect 13723 11398 13775 11450
rect 13787 11398 13839 11450
rect 2320 11271 2372 11280
rect 2320 11237 2329 11271
rect 2329 11237 2363 11271
rect 2363 11237 2372 11271
rect 2320 11228 2372 11237
rect 15752 11271 15804 11280
rect 15752 11237 15761 11271
rect 15761 11237 15795 11271
rect 15795 11237 15804 11271
rect 15752 11228 15804 11237
rect 2136 11092 2188 11144
rect 16212 11135 16264 11144
rect 16212 11101 16221 11135
rect 16221 11101 16255 11135
rect 16255 11101 16264 11135
rect 16212 11092 16264 11101
rect 4135 10854 4187 10906
rect 4199 10854 4251 10906
rect 4263 10854 4315 10906
rect 4327 10854 4379 10906
rect 10441 10854 10493 10906
rect 10505 10854 10557 10906
rect 10569 10854 10621 10906
rect 10633 10854 10685 10906
rect 16748 10854 16800 10906
rect 16812 10854 16864 10906
rect 16876 10854 16928 10906
rect 16940 10854 16992 10906
rect 14648 10795 14700 10804
rect 14648 10761 14657 10795
rect 14657 10761 14691 10795
rect 14691 10761 14700 10795
rect 14648 10752 14700 10761
rect 15752 10684 15804 10736
rect 3976 10616 4028 10668
rect 5172 10591 5224 10600
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 15936 10616 15988 10668
rect 1676 10523 1728 10532
rect 1676 10489 1685 10523
rect 1685 10489 1719 10523
rect 1719 10489 1728 10523
rect 1676 10480 1728 10489
rect 2320 10523 2372 10532
rect 2320 10489 2329 10523
rect 2329 10489 2363 10523
rect 2363 10489 2372 10523
rect 2320 10480 2372 10489
rect 2136 10412 2188 10464
rect 3056 10412 3108 10464
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 7288 10310 7340 10362
rect 7352 10310 7404 10362
rect 7416 10310 7468 10362
rect 7480 10310 7532 10362
rect 13595 10310 13647 10362
rect 13659 10310 13711 10362
rect 13723 10310 13775 10362
rect 13787 10310 13839 10362
rect 1584 10208 1636 10260
rect 1676 10208 1728 10260
rect 3056 10208 3108 10260
rect 15568 10208 15620 10260
rect 112 10072 164 10124
rect 2504 10072 2556 10124
rect 14280 10072 14332 10124
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 15936 9979 15988 9988
rect 15936 9945 15945 9979
rect 15945 9945 15979 9979
rect 15979 9945 15988 9979
rect 15936 9936 15988 9945
rect 1952 9868 2004 9920
rect 4135 9766 4187 9818
rect 4199 9766 4251 9818
rect 4263 9766 4315 9818
rect 4327 9766 4379 9818
rect 10441 9766 10493 9818
rect 10505 9766 10557 9818
rect 10569 9766 10621 9818
rect 10633 9766 10685 9818
rect 16748 9766 16800 9818
rect 16812 9766 16864 9818
rect 16876 9766 16928 9818
rect 16940 9766 16992 9818
rect 15384 9707 15436 9716
rect 15384 9673 15393 9707
rect 15393 9673 15427 9707
rect 15427 9673 15436 9707
rect 15384 9664 15436 9673
rect 2412 9639 2464 9648
rect 2412 9605 2421 9639
rect 2421 9605 2455 9639
rect 2455 9605 2464 9639
rect 2412 9596 2464 9605
rect 1952 9528 2004 9580
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 15936 9528 15988 9537
rect 2688 9460 2740 9512
rect 2136 9435 2188 9444
rect 2136 9401 2145 9435
rect 2145 9401 2179 9435
rect 2179 9401 2188 9435
rect 2136 9392 2188 9401
rect 15568 9435 15620 9444
rect 15568 9401 15577 9435
rect 15577 9401 15611 9435
rect 15611 9401 15620 9435
rect 15568 9392 15620 9401
rect 2504 9324 2556 9376
rect 14280 9367 14332 9376
rect 14280 9333 14289 9367
rect 14289 9333 14323 9367
rect 14323 9333 14332 9367
rect 14280 9324 14332 9333
rect 7288 9222 7340 9274
rect 7352 9222 7404 9274
rect 7416 9222 7468 9274
rect 7480 9222 7532 9274
rect 13595 9222 13647 9274
rect 13659 9222 13711 9274
rect 13723 9222 13775 9274
rect 13787 9222 13839 9274
rect 1492 9120 1544 9172
rect 2504 9120 2556 9172
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 16028 8959 16080 8968
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 16304 8959 16356 8968
rect 16304 8925 16313 8959
rect 16313 8925 16347 8959
rect 16347 8925 16356 8959
rect 16304 8916 16356 8925
rect 15568 8891 15620 8900
rect 15568 8857 15577 8891
rect 15577 8857 15611 8891
rect 15611 8857 15620 8891
rect 15568 8848 15620 8857
rect 4135 8678 4187 8730
rect 4199 8678 4251 8730
rect 4263 8678 4315 8730
rect 4327 8678 4379 8730
rect 10441 8678 10493 8730
rect 10505 8678 10557 8730
rect 10569 8678 10621 8730
rect 10633 8678 10685 8730
rect 16748 8678 16800 8730
rect 16812 8678 16864 8730
rect 16876 8678 16928 8730
rect 16940 8678 16992 8730
rect 12532 8576 12584 8628
rect 16028 8619 16080 8628
rect 16028 8585 16037 8619
rect 16037 8585 16071 8619
rect 16071 8585 16080 8619
rect 16028 8576 16080 8585
rect 2504 8440 2556 8492
rect 2688 8483 2740 8492
rect 2688 8449 2697 8483
rect 2697 8449 2731 8483
rect 2731 8449 2740 8483
rect 2688 8440 2740 8449
rect 3976 8415 4028 8424
rect 3976 8381 3985 8415
rect 3985 8381 4019 8415
rect 4019 8381 4028 8415
rect 3976 8372 4028 8381
rect 17040 8576 17092 8628
rect 1768 8236 1820 8288
rect 13084 8279 13136 8288
rect 13084 8245 13093 8279
rect 13093 8245 13127 8279
rect 13127 8245 13136 8279
rect 13084 8236 13136 8245
rect 7288 8134 7340 8186
rect 7352 8134 7404 8186
rect 7416 8134 7468 8186
rect 7480 8134 7532 8186
rect 13595 8134 13647 8186
rect 13659 8134 13711 8186
rect 13723 8134 13775 8186
rect 13787 8134 13839 8186
rect 1768 8075 1820 8084
rect 1768 8041 1777 8075
rect 1777 8041 1811 8075
rect 1811 8041 1820 8075
rect 1768 8032 1820 8041
rect 13084 8032 13136 8084
rect 12900 7896 12952 7948
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 12072 7871 12124 7880
rect 12072 7837 12081 7871
rect 12081 7837 12115 7871
rect 12115 7837 12124 7871
rect 12072 7828 12124 7837
rect 16028 7871 16080 7880
rect 16028 7837 16037 7871
rect 16037 7837 16071 7871
rect 16071 7837 16080 7871
rect 16028 7828 16080 7837
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 4135 7590 4187 7642
rect 4199 7590 4251 7642
rect 4263 7590 4315 7642
rect 4327 7590 4379 7642
rect 10441 7590 10493 7642
rect 10505 7590 10557 7642
rect 10569 7590 10621 7642
rect 10633 7590 10685 7642
rect 16748 7590 16800 7642
rect 16812 7590 16864 7642
rect 16876 7590 16928 7642
rect 16940 7590 16992 7642
rect 12072 7488 12124 7540
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 2228 7352 2280 7404
rect 15200 7488 15252 7540
rect 16028 7531 16080 7540
rect 16028 7497 16037 7531
rect 16037 7497 16071 7531
rect 16071 7497 16080 7531
rect 16028 7488 16080 7497
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 14096 7284 14148 7293
rect 5264 7259 5316 7268
rect 5264 7225 5273 7259
rect 5273 7225 5307 7259
rect 5307 7225 5316 7259
rect 5264 7216 5316 7225
rect 17868 7148 17920 7200
rect 7288 7046 7340 7098
rect 7352 7046 7404 7098
rect 7416 7046 7468 7098
rect 7480 7046 7532 7098
rect 13595 7046 13647 7098
rect 13659 7046 13711 7098
rect 13723 7046 13775 7098
rect 13787 7046 13839 7098
rect 5264 6944 5316 6996
rect 14096 6944 14148 6996
rect 12900 6919 12952 6928
rect 12900 6885 12909 6919
rect 12909 6885 12943 6919
rect 12943 6885 12952 6919
rect 12900 6876 12952 6885
rect 5540 6808 5592 6860
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 1860 6783 1912 6792
rect 1860 6749 1869 6783
rect 1869 6749 1903 6783
rect 1903 6749 1912 6783
rect 1860 6740 1912 6749
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 11888 6740 11940 6792
rect 4135 6502 4187 6554
rect 4199 6502 4251 6554
rect 4263 6502 4315 6554
rect 4327 6502 4379 6554
rect 10441 6502 10493 6554
rect 10505 6502 10557 6554
rect 10569 6502 10621 6554
rect 10633 6502 10685 6554
rect 16748 6502 16800 6554
rect 16812 6502 16864 6554
rect 16876 6502 16928 6554
rect 16940 6502 16992 6554
rect 13728 6375 13780 6384
rect 13728 6341 13737 6375
rect 13737 6341 13771 6375
rect 13771 6341 13780 6375
rect 13728 6332 13780 6341
rect 1860 6264 1912 6316
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 11888 6264 11940 6316
rect 1676 6128 1728 6180
rect 5540 6103 5592 6112
rect 5540 6069 5549 6103
rect 5549 6069 5583 6103
rect 5583 6069 5592 6103
rect 5540 6060 5592 6069
rect 6460 6060 6512 6112
rect 12532 6171 12584 6180
rect 12532 6137 12541 6171
rect 12541 6137 12575 6171
rect 12575 6137 12584 6171
rect 12532 6128 12584 6137
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 11888 6060 11940 6069
rect 7288 5958 7340 6010
rect 7352 5958 7404 6010
rect 7416 5958 7468 6010
rect 7480 5958 7532 6010
rect 13595 5958 13647 6010
rect 13659 5958 13711 6010
rect 13723 5958 13775 6010
rect 13787 5958 13839 6010
rect 12532 5856 12584 5908
rect 9312 5788 9364 5840
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 6276 5720 6328 5729
rect 12992 5720 13044 5772
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 11428 5695 11480 5704
rect 11428 5661 11437 5695
rect 11437 5661 11471 5695
rect 11471 5661 11480 5695
rect 11428 5652 11480 5661
rect 11888 5695 11940 5704
rect 11888 5661 11897 5695
rect 11897 5661 11931 5695
rect 11931 5661 11940 5695
rect 11888 5652 11940 5661
rect 7012 5516 7064 5568
rect 10232 5559 10284 5568
rect 10232 5525 10241 5559
rect 10241 5525 10275 5559
rect 10275 5525 10284 5559
rect 10232 5516 10284 5525
rect 4135 5414 4187 5466
rect 4199 5414 4251 5466
rect 4263 5414 4315 5466
rect 4327 5414 4379 5466
rect 10441 5414 10493 5466
rect 10505 5414 10557 5466
rect 10569 5414 10621 5466
rect 10633 5414 10685 5466
rect 16748 5414 16800 5466
rect 16812 5414 16864 5466
rect 16876 5414 16928 5466
rect 16940 5414 16992 5466
rect 112 5312 164 5364
rect 6276 5355 6328 5364
rect 6276 5321 6285 5355
rect 6285 5321 6319 5355
rect 6319 5321 6328 5355
rect 6276 5312 6328 5321
rect 7012 5355 7064 5364
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 8116 5312 8168 5364
rect 9496 5312 9548 5364
rect 11428 5355 11480 5364
rect 11428 5321 11437 5355
rect 11437 5321 11471 5355
rect 11471 5321 11480 5355
rect 11428 5312 11480 5321
rect 12992 5355 13044 5364
rect 12992 5321 13001 5355
rect 13001 5321 13035 5355
rect 13035 5321 13044 5355
rect 12992 5312 13044 5321
rect 6368 4972 6420 5024
rect 10232 4972 10284 5024
rect 11612 4972 11664 5024
rect 7288 4870 7340 4922
rect 7352 4870 7404 4922
rect 7416 4870 7468 4922
rect 7480 4870 7532 4922
rect 13595 4870 13647 4922
rect 13659 4870 13711 4922
rect 13723 4870 13775 4922
rect 13787 4870 13839 4922
rect 8024 4700 8076 4752
rect 8116 4700 8168 4752
rect 13268 4632 13320 4684
rect 9680 4607 9732 4616
rect 9680 4573 9689 4607
rect 9689 4573 9723 4607
rect 9723 4573 9732 4607
rect 9680 4564 9732 4573
rect 10784 4564 10836 4616
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 12348 4428 12400 4480
rect 4135 4326 4187 4378
rect 4199 4326 4251 4378
rect 4263 4326 4315 4378
rect 4327 4326 4379 4378
rect 10441 4326 10493 4378
rect 10505 4326 10557 4378
rect 10569 4326 10621 4378
rect 10633 4326 10685 4378
rect 16748 4326 16800 4378
rect 16812 4326 16864 4378
rect 16876 4326 16928 4378
rect 16940 4326 16992 4378
rect 7656 4267 7708 4276
rect 7656 4233 7665 4267
rect 7665 4233 7699 4267
rect 7699 4233 7708 4267
rect 7656 4224 7708 4233
rect 1584 4088 1636 4140
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 9680 4156 9732 4208
rect 10784 4088 10836 4140
rect 14924 4063 14976 4072
rect 14924 4029 14942 4063
rect 14942 4029 14976 4063
rect 14924 4020 14976 4029
rect 9312 3995 9364 4004
rect 9312 3961 9321 3995
rect 9321 3961 9355 3995
rect 9355 3961 9364 3995
rect 9312 3952 9364 3961
rect 11612 3952 11664 4004
rect 7656 3884 7708 3936
rect 8024 3927 8076 3936
rect 8024 3893 8033 3927
rect 8033 3893 8067 3927
rect 8067 3893 8076 3927
rect 8024 3884 8076 3893
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 13268 3884 13320 3936
rect 15384 3884 15436 3936
rect 15660 3884 15712 3936
rect 16580 3884 16632 3936
rect 7288 3782 7340 3834
rect 7352 3782 7404 3834
rect 7416 3782 7468 3834
rect 7480 3782 7532 3834
rect 13595 3782 13647 3834
rect 13659 3782 13711 3834
rect 13723 3782 13775 3834
rect 13787 3782 13839 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 8024 3680 8076 3732
rect 7656 3612 7708 3664
rect 9312 3612 9364 3664
rect 15384 3655 15436 3664
rect 15384 3621 15393 3655
rect 15393 3621 15427 3655
rect 15427 3621 15436 3655
rect 15384 3612 15436 3621
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 8024 3544 8076 3596
rect 13912 3544 13964 3596
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7012 3476 7064 3485
rect 9036 3476 9088 3528
rect 10876 3476 10928 3528
rect 11336 3519 11388 3528
rect 11336 3485 11345 3519
rect 11345 3485 11379 3519
rect 11379 3485 11388 3519
rect 11336 3476 11388 3485
rect 11612 3519 11664 3528
rect 11612 3485 11621 3519
rect 11621 3485 11655 3519
rect 11655 3485 11664 3519
rect 11612 3476 11664 3485
rect 15752 3519 15804 3528
rect 15752 3485 15761 3519
rect 15761 3485 15795 3519
rect 15795 3485 15804 3519
rect 15752 3476 15804 3485
rect 14188 3340 14240 3392
rect 4135 3238 4187 3290
rect 4199 3238 4251 3290
rect 4263 3238 4315 3290
rect 4327 3238 4379 3290
rect 10441 3238 10493 3290
rect 10505 3238 10557 3290
rect 10569 3238 10621 3290
rect 10633 3238 10685 3290
rect 16748 3238 16800 3290
rect 16812 3238 16864 3290
rect 16876 3238 16928 3290
rect 16940 3238 16992 3290
rect 112 3136 164 3188
rect 1400 3136 1452 3188
rect 8024 3179 8076 3188
rect 8024 3145 8033 3179
rect 8033 3145 8067 3179
rect 8067 3145 8076 3179
rect 8024 3136 8076 3145
rect 9036 3179 9088 3188
rect 9036 3145 9045 3179
rect 9045 3145 9079 3179
rect 9079 3145 9088 3179
rect 9036 3136 9088 3145
rect 11336 3179 11388 3188
rect 11336 3145 11345 3179
rect 11345 3145 11379 3179
rect 11379 3145 11388 3179
rect 11336 3136 11388 3145
rect 12440 3136 12492 3188
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 15752 3136 15804 3188
rect 7012 2796 7064 2848
rect 7748 2796 7800 2848
rect 8484 2796 8536 2848
rect 10876 2907 10928 2916
rect 10876 2873 10885 2907
rect 10885 2873 10919 2907
rect 10919 2873 10928 2907
rect 10876 2864 10928 2873
rect 14188 3043 14240 3052
rect 14188 3009 14197 3043
rect 14197 3009 14231 3043
rect 14231 3009 14240 3043
rect 14188 3000 14240 3009
rect 15752 3043 15804 3052
rect 15752 3009 15761 3043
rect 15761 3009 15795 3043
rect 15795 3009 15804 3043
rect 15752 3000 15804 3009
rect 10324 2796 10376 2848
rect 13912 2796 13964 2848
rect 14556 2796 14608 2848
rect 7288 2694 7340 2746
rect 7352 2694 7404 2746
rect 7416 2694 7468 2746
rect 7480 2694 7532 2746
rect 13595 2694 13647 2746
rect 13659 2694 13711 2746
rect 13723 2694 13775 2746
rect 13787 2694 13839 2746
rect 12348 2635 12400 2644
rect 12348 2601 12357 2635
rect 12357 2601 12391 2635
rect 12391 2601 12400 2635
rect 12348 2592 12400 2601
rect 14188 2635 14240 2644
rect 14188 2601 14197 2635
rect 14197 2601 14231 2635
rect 14231 2601 14240 2635
rect 14188 2592 14240 2601
rect 10876 2524 10928 2576
rect 13452 2524 13504 2576
rect 8484 2456 8536 2508
rect 9496 2320 9548 2372
rect 11428 2320 11480 2372
rect 13452 2320 13504 2372
rect 15660 2431 15712 2440
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 15384 2320 15436 2372
rect 4135 2150 4187 2202
rect 4199 2150 4251 2202
rect 4263 2150 4315 2202
rect 4327 2150 4379 2202
rect 10441 2150 10493 2202
rect 10505 2150 10557 2202
rect 10569 2150 10621 2202
rect 10633 2150 10685 2202
rect 16748 2150 16800 2202
rect 16812 2150 16864 2202
rect 16876 2150 16928 2202
rect 16940 2150 16992 2202
rect 11060 76 11112 128
rect 11888 76 11940 128
<< metal2 >>
rect 478 20583 534 21063
rect 1398 20618 1454 21063
rect 2410 20618 2466 21063
rect 1398 20590 1716 20618
rect 1398 20583 1454 20590
rect 18 20496 74 20505
rect 18 20431 74 20440
rect 32 17882 60 20431
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 20 17876 72 17882
rect 20 17818 72 17824
rect 1412 17746 1440 18022
rect 1582 17912 1638 17921
rect 1582 17847 1638 17856
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 112 17536 164 17542
rect 112 17478 164 17484
rect 124 16289 152 17478
rect 1412 17338 1440 17682
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1490 16824 1546 16833
rect 1490 16759 1546 16768
rect 110 16280 166 16289
rect 110 16215 166 16224
rect 1122 14648 1178 14657
rect 1122 14583 1178 14592
rect 110 14104 166 14113
rect 110 14039 166 14048
rect 124 14006 152 14039
rect 112 14000 164 14006
rect 112 13942 164 13948
rect 1136 13870 1164 14583
rect 1124 13864 1176 13870
rect 1124 13806 1176 13812
rect 112 12164 164 12170
rect 112 12106 164 12112
rect 124 12073 152 12106
rect 110 12064 166 12073
rect 110 11999 166 12008
rect 112 10124 164 10130
rect 112 10066 164 10072
rect 124 9897 152 10066
rect 110 9888 166 9897
rect 110 9823 166 9832
rect 1504 9178 1532 16759
rect 1596 13530 1624 17847
rect 1688 17785 1716 20590
rect 2410 20590 2728 20618
rect 2410 20583 2466 20590
rect 2700 18222 2728 20590
rect 3422 20583 3478 21063
rect 4434 20583 4490 21063
rect 5446 20583 5502 21063
rect 6458 20618 6514 21063
rect 6196 20590 6514 20618
rect 2136 18216 2188 18222
rect 2136 18158 2188 18164
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 1674 17776 1730 17785
rect 1674 17711 1730 17720
rect 2056 16726 2084 18022
rect 2044 16720 2096 16726
rect 2044 16662 2096 16668
rect 2056 16250 2084 16662
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2148 16114 2176 18158
rect 3240 17808 3292 17814
rect 3240 17750 3292 17756
rect 3252 17338 3280 17750
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 2320 17060 2372 17066
rect 2320 17002 2372 17008
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2148 15638 2176 16050
rect 2240 15978 2268 16526
rect 2228 15972 2280 15978
rect 2228 15914 2280 15920
rect 2136 15632 2188 15638
rect 2136 15574 2188 15580
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1780 15162 1808 15438
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1688 13870 1716 14962
rect 2240 14550 2268 15914
rect 2228 14544 2280 14550
rect 2228 14486 2280 14492
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 2240 13734 2268 14350
rect 2332 13802 2360 17002
rect 3436 16561 3464 20583
rect 4109 18524 4405 18544
rect 4165 18522 4189 18524
rect 4245 18522 4269 18524
rect 4325 18522 4349 18524
rect 4187 18470 4189 18522
rect 4251 18470 4263 18522
rect 4325 18470 4327 18522
rect 4165 18468 4189 18470
rect 4245 18468 4269 18470
rect 4325 18468 4349 18470
rect 4109 18448 4405 18468
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3422 16552 3478 16561
rect 3422 16487 3478 16496
rect 3896 16250 3924 17478
rect 3988 17338 4016 18022
rect 4448 17814 4476 20583
rect 4986 18728 5042 18737
rect 4986 18663 5042 18672
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4908 17814 4936 18158
rect 4436 17808 4488 17814
rect 4436 17750 4488 17756
rect 4896 17808 4948 17814
rect 4896 17750 4948 17756
rect 4436 17604 4488 17610
rect 4436 17546 4488 17552
rect 4109 17436 4405 17456
rect 4165 17434 4189 17436
rect 4245 17434 4269 17436
rect 4325 17434 4349 17436
rect 4187 17382 4189 17434
rect 4251 17382 4263 17434
rect 4325 17382 4327 17434
rect 4165 17380 4189 17382
rect 4245 17380 4269 17382
rect 4325 17380 4349 17382
rect 4109 17360 4405 17380
rect 3976 17332 4028 17338
rect 3976 17274 4028 17280
rect 4448 16998 4476 17546
rect 4908 17202 4936 17750
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 4448 16794 4476 16934
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 4109 16348 4405 16368
rect 4165 16346 4189 16348
rect 4245 16346 4269 16348
rect 4325 16346 4349 16348
rect 4187 16294 4189 16346
rect 4251 16294 4263 16346
rect 4325 16294 4327 16346
rect 4165 16292 4189 16294
rect 4245 16292 4269 16294
rect 4325 16292 4349 16294
rect 4109 16272 4405 16292
rect 3884 16244 3936 16250
rect 3884 16186 3936 16192
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4109 15260 4405 15280
rect 4165 15258 4189 15260
rect 4245 15258 4269 15260
rect 4325 15258 4349 15260
rect 4187 15206 4189 15258
rect 4251 15206 4263 15258
rect 4325 15206 4327 15258
rect 4165 15204 4189 15206
rect 4245 15204 4269 15206
rect 4325 15204 4349 15206
rect 4109 15184 4405 15204
rect 4448 15026 4476 16050
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 2596 14884 2648 14890
rect 2596 14826 2648 14832
rect 3608 14884 3660 14890
rect 3608 14826 3660 14832
rect 2608 14618 2636 14826
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2608 14346 2636 14554
rect 2596 14340 2648 14346
rect 2596 14282 2648 14288
rect 2608 13920 2636 14282
rect 2688 13932 2740 13938
rect 2608 13892 2688 13920
rect 2688 13874 2740 13880
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2320 13796 2372 13802
rect 2320 13738 2372 13744
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2056 13190 2084 13330
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1596 11762 1624 12038
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1596 10266 1624 11698
rect 1676 10532 1728 10538
rect 1676 10474 1728 10480
rect 1688 10266 1716 10474
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1872 8401 1900 12718
rect 2056 12374 2084 13126
rect 2240 12986 2268 13670
rect 2976 13394 3004 13874
rect 3620 13530 3648 14826
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 14074 4016 14350
rect 4109 14172 4405 14192
rect 4165 14170 4189 14172
rect 4245 14170 4269 14172
rect 4325 14170 4349 14172
rect 4187 14118 4189 14170
rect 4251 14118 4263 14170
rect 4325 14118 4327 14170
rect 4165 14116 4189 14118
rect 4245 14116 4269 14118
rect 4325 14116 4349 14118
rect 4109 14096 4405 14116
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 5000 13870 5028 18663
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 5092 16658 5120 18022
rect 5460 16794 5488 20583
rect 6092 17876 6144 17882
rect 6092 17818 6144 17824
rect 6104 17134 6132 17818
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 6196 16794 6224 20590
rect 6458 20583 6514 20590
rect 7378 20618 7434 21063
rect 8390 20618 8446 21063
rect 7378 20590 7696 20618
rect 7378 20583 7434 20590
rect 7262 17980 7558 18000
rect 7318 17978 7342 17980
rect 7398 17978 7422 17980
rect 7478 17978 7502 17980
rect 7340 17926 7342 17978
rect 7404 17926 7416 17978
rect 7478 17926 7480 17978
rect 7318 17924 7342 17926
rect 7398 17924 7422 17926
rect 7478 17924 7502 17926
rect 7262 17904 7558 17924
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6656 16998 6684 17614
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 5092 16250 5120 16594
rect 6012 16250 6040 16594
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 6196 15162 6224 15574
rect 6564 15502 6592 16050
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 5172 14884 5224 14890
rect 5172 14826 5224 14832
rect 5184 14618 5212 14826
rect 6656 14618 6684 16934
rect 7262 16892 7558 16912
rect 7318 16890 7342 16892
rect 7398 16890 7422 16892
rect 7478 16890 7502 16892
rect 7340 16838 7342 16890
rect 7404 16838 7416 16890
rect 7478 16838 7480 16890
rect 7318 16836 7342 16838
rect 7398 16836 7422 16838
rect 7478 16836 7502 16838
rect 7262 16816 7558 16836
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 6748 15026 6776 15914
rect 7262 15804 7558 15824
rect 7318 15802 7342 15804
rect 7398 15802 7422 15804
rect 7478 15802 7502 15804
rect 7340 15750 7342 15802
rect 7404 15750 7416 15802
rect 7478 15750 7480 15802
rect 7318 15748 7342 15750
rect 7398 15748 7422 15750
rect 7478 15748 7502 15750
rect 7262 15728 7558 15748
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 7262 14716 7558 14736
rect 7318 14714 7342 14716
rect 7398 14714 7422 14716
rect 7478 14714 7502 14716
rect 7340 14662 7342 14714
rect 7404 14662 7416 14714
rect 7478 14662 7480 14714
rect 7318 14660 7342 14662
rect 7398 14660 7422 14662
rect 7478 14660 7502 14662
rect 7262 14640 7558 14660
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 5644 14006 5672 14418
rect 7116 14074 7144 14418
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 7262 13628 7558 13648
rect 7318 13626 7342 13628
rect 7398 13626 7422 13628
rect 7478 13626 7502 13628
rect 7340 13574 7342 13626
rect 7404 13574 7416 13626
rect 7478 13574 7480 13626
rect 7318 13572 7342 13574
rect 7398 13572 7422 13574
rect 7478 13572 7502 13574
rect 7262 13552 7558 13572
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 2516 12306 2544 13126
rect 2976 12918 3004 13330
rect 2964 12912 3016 12918
rect 2964 12854 3016 12860
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2516 11898 2544 12242
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 2332 11286 2360 11562
rect 2320 11280 2372 11286
rect 2320 11222 2372 11228
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2148 10470 2176 11086
rect 2320 10532 2372 10538
rect 2320 10474 2372 10480
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1964 9586 1992 9862
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 2148 9450 2176 10406
rect 2136 9444 2188 9450
rect 2136 9386 2188 9392
rect 1858 8392 1914 8401
rect 1858 8327 1914 8336
rect 1768 8288 1820 8294
rect 1768 8230 1820 8236
rect 1780 8090 1808 8230
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1780 7410 1808 8026
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1674 6352 1730 6361
rect 1872 6322 1900 6734
rect 1674 6287 1730 6296
rect 1860 6316 1912 6322
rect 1688 6186 1716 6287
rect 1860 6258 1912 6264
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 110 5672 166 5681
rect 110 5607 166 5616
rect 124 5370 152 5607
rect 112 5364 164 5370
rect 112 5306 164 5312
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1596 4146 1624 4422
rect 2148 4146 2176 9386
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2240 7410 2268 7822
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2332 6798 2360 10474
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2516 9674 2544 10066
rect 2424 9654 2544 9674
rect 2412 9648 2544 9654
rect 2464 9646 2544 9648
rect 2412 9590 2464 9596
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2516 9178 2544 9318
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2516 8498 2544 8910
rect 2700 8498 2728 9454
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2700 7886 2728 8434
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2792 5273 2820 12582
rect 2976 12442 3004 12854
rect 3988 12646 4016 13330
rect 4109 13084 4405 13104
rect 4165 13082 4189 13084
rect 4245 13082 4269 13084
rect 4325 13082 4349 13084
rect 4187 13030 4189 13082
rect 4251 13030 4263 13082
rect 4325 13030 4327 13082
rect 4165 13028 4189 13030
rect 4245 13028 4269 13030
rect 4325 13028 4349 13030
rect 4109 13008 4405 13028
rect 5262 12744 5318 12753
rect 5262 12679 5318 12688
rect 5276 12646 5304 12679
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5736 12442 5764 12582
rect 7262 12540 7558 12560
rect 7318 12538 7342 12540
rect 7398 12538 7422 12540
rect 7478 12538 7502 12540
rect 7340 12486 7342 12538
rect 7404 12486 7416 12538
rect 7478 12486 7480 12538
rect 7318 12484 7342 12486
rect 7398 12484 7422 12486
rect 7478 12484 7502 12486
rect 7262 12464 7558 12484
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 11762 3924 12174
rect 4109 11996 4405 12016
rect 4165 11994 4189 11996
rect 4245 11994 4269 11996
rect 4325 11994 4349 11996
rect 4187 11942 4189 11994
rect 4251 11942 4263 11994
rect 4325 11942 4327 11994
rect 4165 11940 4189 11942
rect 4245 11940 4269 11942
rect 4325 11940 4349 11942
rect 4109 11920 4405 11940
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3988 10674 4016 11698
rect 5092 11558 5120 12242
rect 6288 11898 6316 12242
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 7262 11452 7558 11472
rect 7318 11450 7342 11452
rect 7398 11450 7422 11452
rect 7478 11450 7502 11452
rect 7340 11398 7342 11450
rect 7404 11398 7416 11450
rect 7478 11398 7480 11450
rect 7318 11396 7342 11398
rect 7398 11396 7422 11398
rect 7478 11396 7502 11398
rect 7262 11376 7558 11396
rect 4109 10908 4405 10928
rect 4165 10906 4189 10908
rect 4245 10906 4269 10908
rect 4325 10906 4349 10908
rect 4187 10854 4189 10906
rect 4251 10854 4263 10906
rect 4325 10854 4327 10906
rect 4165 10852 4189 10854
rect 4245 10852 4269 10854
rect 4325 10852 4349 10854
rect 4109 10832 4405 10852
rect 5170 10704 5226 10713
rect 3976 10668 4028 10674
rect 5170 10639 5226 10648
rect 3976 10610 4028 10616
rect 5184 10606 5212 10639
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 3068 10266 3096 10406
rect 7262 10364 7558 10384
rect 7318 10362 7342 10364
rect 7398 10362 7422 10364
rect 7478 10362 7502 10364
rect 7340 10310 7342 10362
rect 7404 10310 7416 10362
rect 7478 10310 7480 10362
rect 7318 10308 7342 10310
rect 7398 10308 7422 10310
rect 7478 10308 7502 10310
rect 7262 10288 7558 10308
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 4109 9820 4405 9840
rect 4165 9818 4189 9820
rect 4245 9818 4269 9820
rect 4325 9818 4349 9820
rect 4187 9766 4189 9818
rect 4251 9766 4263 9818
rect 4325 9766 4327 9818
rect 4165 9764 4189 9766
rect 4245 9764 4269 9766
rect 4325 9764 4349 9766
rect 4109 9744 4405 9764
rect 7262 9276 7558 9296
rect 7318 9274 7342 9276
rect 7398 9274 7422 9276
rect 7478 9274 7502 9276
rect 7340 9222 7342 9274
rect 7404 9222 7416 9274
rect 7478 9222 7480 9274
rect 7318 9220 7342 9222
rect 7398 9220 7422 9222
rect 7478 9220 7502 9222
rect 7262 9200 7558 9220
rect 4109 8732 4405 8752
rect 4165 8730 4189 8732
rect 4245 8730 4269 8732
rect 4325 8730 4349 8732
rect 4187 8678 4189 8730
rect 4251 8678 4263 8730
rect 4325 8678 4327 8730
rect 4165 8676 4189 8678
rect 4245 8676 4269 8678
rect 4325 8676 4349 8678
rect 4109 8656 4405 8676
rect 3974 8528 4030 8537
rect 3974 8463 4030 8472
rect 3988 8430 4016 8463
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 7262 8188 7558 8208
rect 7318 8186 7342 8188
rect 7398 8186 7422 8188
rect 7478 8186 7502 8188
rect 7340 8134 7342 8186
rect 7404 8134 7416 8186
rect 7478 8134 7480 8186
rect 7318 8132 7342 8134
rect 7398 8132 7422 8134
rect 7478 8132 7502 8134
rect 7262 8112 7558 8132
rect 4109 7644 4405 7664
rect 4165 7642 4189 7644
rect 4245 7642 4269 7644
rect 4325 7642 4349 7644
rect 4187 7590 4189 7642
rect 4251 7590 4263 7642
rect 4325 7590 4327 7642
rect 4165 7588 4189 7590
rect 4245 7588 4269 7590
rect 4325 7588 4349 7590
rect 4109 7568 4405 7588
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5276 7002 5304 7210
rect 7262 7100 7558 7120
rect 7318 7098 7342 7100
rect 7398 7098 7422 7100
rect 7478 7098 7502 7100
rect 7340 7046 7342 7098
rect 7404 7046 7416 7098
rect 7478 7046 7480 7098
rect 7318 7044 7342 7046
rect 7398 7044 7422 7046
rect 7478 7044 7502 7046
rect 7262 7024 7558 7044
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 4109 6556 4405 6576
rect 4165 6554 4189 6556
rect 4245 6554 4269 6556
rect 4325 6554 4349 6556
rect 4187 6502 4189 6554
rect 4251 6502 4263 6554
rect 4325 6502 4327 6554
rect 4165 6500 4189 6502
rect 4245 6500 4269 6502
rect 4325 6500 4349 6502
rect 4109 6480 4405 6500
rect 5552 6118 5580 6802
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 4109 5468 4405 5488
rect 4165 5466 4189 5468
rect 4245 5466 4269 5468
rect 4325 5466 4349 5468
rect 4187 5414 4189 5466
rect 4251 5414 4263 5466
rect 4325 5414 4327 5466
rect 4165 5412 4189 5414
rect 4245 5412 4269 5414
rect 4325 5412 4349 5414
rect 4109 5392 4405 5412
rect 6288 5370 6316 5714
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 2778 5264 2834 5273
rect 2778 5199 2834 5208
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 4109 4380 4405 4400
rect 4165 4378 4189 4380
rect 4245 4378 4269 4380
rect 4325 4378 4349 4380
rect 4187 4326 4189 4378
rect 4251 4326 4263 4378
rect 4325 4326 4327 4378
rect 4165 4324 4189 4326
rect 4245 4324 4269 4326
rect 4325 4324 4349 4326
rect 4109 4304 4405 4324
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 1596 3738 1624 4082
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 110 3632 166 3641
rect 110 3567 166 3576
rect 1400 3596 1452 3602
rect 124 3194 152 3567
rect 1400 3538 1452 3544
rect 1412 3194 1440 3538
rect 4109 3292 4405 3312
rect 4165 3290 4189 3292
rect 4245 3290 4269 3292
rect 4325 3290 4349 3292
rect 4187 3238 4189 3290
rect 4251 3238 4263 3290
rect 4325 3238 4327 3290
rect 4165 3236 4189 3238
rect 4245 3236 4269 3238
rect 4325 3236 4349 3238
rect 4109 3216 4405 3236
rect 112 3188 164 3194
rect 112 3130 164 3136
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 6380 3097 6408 4966
rect 6366 3088 6422 3097
rect 6366 3023 6422 3032
rect 4109 2204 4405 2224
rect 4165 2202 4189 2204
rect 4245 2202 4269 2204
rect 4325 2202 4349 2204
rect 4187 2150 4189 2202
rect 4251 2150 4263 2202
rect 4325 2150 4327 2202
rect 4165 2148 4189 2150
rect 4245 2148 4269 2150
rect 4325 2148 4349 2150
rect 4109 2128 4405 2148
rect 570 0 626 480
rect 1766 0 1822 480
rect 3054 0 3110 480
rect 4342 0 4398 480
rect 5538 0 5594 480
rect 6472 82 6500 6054
rect 7262 6012 7558 6032
rect 7318 6010 7342 6012
rect 7398 6010 7422 6012
rect 7478 6010 7502 6012
rect 7340 5958 7342 6010
rect 7404 5958 7416 6010
rect 7478 5958 7480 6010
rect 7318 5956 7342 5958
rect 7398 5956 7422 5958
rect 7478 5956 7502 5958
rect 7262 5936 7558 5956
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7024 5370 7052 5510
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7262 4924 7558 4944
rect 7318 4922 7342 4924
rect 7398 4922 7422 4924
rect 7478 4922 7502 4924
rect 7340 4870 7342 4922
rect 7404 4870 7416 4922
rect 7478 4870 7480 4922
rect 7318 4868 7342 4870
rect 7398 4868 7422 4870
rect 7478 4868 7502 4870
rect 7262 4848 7558 4868
rect 7668 4282 7696 20590
rect 8128 20590 8446 20618
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 7944 17746 7972 18022
rect 8128 17882 8156 20590
rect 8390 20583 8446 20590
rect 9402 20618 9458 21063
rect 10414 20618 10470 21063
rect 9402 20590 9536 20618
rect 9402 20583 9458 20590
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 8116 17876 8168 17882
rect 8116 17818 8168 17824
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 7944 17338 7972 17682
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 8496 17202 8524 18158
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8668 18148 8720 18154
rect 8668 18090 8720 18096
rect 8588 17338 8616 18090
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 8220 16590 8248 17002
rect 8496 16590 8524 17138
rect 8588 17066 8616 17274
rect 8576 17060 8628 17066
rect 8576 17002 8628 17008
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8220 16046 8248 16526
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8128 15638 8156 15846
rect 8220 15638 8248 15982
rect 8116 15632 8168 15638
rect 8116 15574 8168 15580
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8128 15162 8156 15574
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8680 13938 8708 18090
rect 8944 16040 8996 16046
rect 8942 16008 8944 16017
rect 8996 16008 8998 16017
rect 8942 15943 8998 15952
rect 8956 15910 8984 15943
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9324 5846 9352 6258
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8128 5370 8156 5646
rect 9508 5370 9536 20590
rect 10244 20590 10470 20618
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9968 17338 9996 18022
rect 10244 17882 10272 20590
rect 10414 20583 10470 20590
rect 11426 20583 11482 21063
rect 12438 20583 12494 21063
rect 12532 20596 12584 20602
rect 10415 18524 10711 18544
rect 10471 18522 10495 18524
rect 10551 18522 10575 18524
rect 10631 18522 10655 18524
rect 10493 18470 10495 18522
rect 10557 18470 10569 18522
rect 10631 18470 10633 18522
rect 10471 18468 10495 18470
rect 10551 18468 10575 18470
rect 10631 18468 10655 18470
rect 10415 18448 10711 18468
rect 11440 18426 11468 20583
rect 11428 18420 11480 18426
rect 11428 18362 11480 18368
rect 11440 18222 11468 18362
rect 11428 18216 11480 18222
rect 11428 18158 11480 18164
rect 11612 18216 11664 18222
rect 11612 18158 11664 18164
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 11532 17814 11560 18022
rect 11520 17808 11572 17814
rect 11624 17785 11652 18158
rect 11520 17750 11572 17756
rect 11610 17776 11666 17785
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 10060 16998 10088 17682
rect 10415 17436 10711 17456
rect 10471 17434 10495 17436
rect 10551 17434 10575 17436
rect 10631 17434 10655 17436
rect 10493 17382 10495 17434
rect 10557 17382 10569 17434
rect 10631 17382 10633 17434
rect 10471 17380 10495 17382
rect 10551 17380 10575 17382
rect 10631 17380 10655 17382
rect 10415 17360 10711 17380
rect 11532 17338 11560 17750
rect 11610 17711 11666 17720
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 12176 17202 12204 17614
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 11888 17060 11940 17066
rect 11888 17002 11940 17008
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10060 15910 10088 16526
rect 10336 16114 10364 16526
rect 10415 16348 10711 16368
rect 10471 16346 10495 16348
rect 10551 16346 10575 16348
rect 10631 16346 10655 16348
rect 10493 16294 10495 16346
rect 10557 16294 10569 16346
rect 10631 16294 10633 16346
rect 10471 16292 10495 16294
rect 10551 16292 10575 16294
rect 10631 16292 10655 16294
rect 10415 16272 10711 16292
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10796 15910 10824 16934
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11624 16182 11652 16662
rect 11900 16590 11928 17002
rect 12176 16794 12204 17138
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11900 16250 11928 16526
rect 11888 16244 11940 16250
rect 11888 16186 11940 16192
rect 11612 16176 11664 16182
rect 11612 16118 11664 16124
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 9600 15026 9628 15846
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10336 15162 10364 15438
rect 10415 15260 10711 15280
rect 10471 15258 10495 15260
rect 10551 15258 10575 15260
rect 10631 15258 10655 15260
rect 10493 15206 10495 15258
rect 10557 15206 10569 15258
rect 10631 15206 10633 15258
rect 10471 15204 10495 15206
rect 10551 15204 10575 15206
rect 10631 15204 10655 15206
rect 10415 15184 10711 15204
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10415 14172 10711 14192
rect 10471 14170 10495 14172
rect 10551 14170 10575 14172
rect 10631 14170 10655 14172
rect 10493 14118 10495 14170
rect 10557 14118 10569 14170
rect 10631 14118 10633 14170
rect 10471 14116 10495 14118
rect 10551 14116 10575 14118
rect 10631 14116 10655 14118
rect 10415 14096 10711 14116
rect 10415 13084 10711 13104
rect 10471 13082 10495 13084
rect 10551 13082 10575 13084
rect 10631 13082 10655 13084
rect 10493 13030 10495 13082
rect 10557 13030 10569 13082
rect 10631 13030 10633 13082
rect 10471 13028 10495 13030
rect 10551 13028 10575 13030
rect 10631 13028 10655 13030
rect 10415 13008 10711 13028
rect 10415 11996 10711 12016
rect 10471 11994 10495 11996
rect 10551 11994 10575 11996
rect 10631 11994 10655 11996
rect 10493 11942 10495 11994
rect 10557 11942 10569 11994
rect 10631 11942 10633 11994
rect 10471 11940 10495 11942
rect 10551 11940 10575 11942
rect 10631 11940 10655 11942
rect 10415 11920 10711 11940
rect 10415 10908 10711 10928
rect 10471 10906 10495 10908
rect 10551 10906 10575 10908
rect 10631 10906 10655 10908
rect 10493 10854 10495 10906
rect 10557 10854 10569 10906
rect 10631 10854 10633 10906
rect 10471 10852 10495 10854
rect 10551 10852 10575 10854
rect 10631 10852 10655 10854
rect 10415 10832 10711 10852
rect 10415 9820 10711 9840
rect 10471 9818 10495 9820
rect 10551 9818 10575 9820
rect 10631 9818 10655 9820
rect 10493 9766 10495 9818
rect 10557 9766 10569 9818
rect 10631 9766 10633 9818
rect 10471 9764 10495 9766
rect 10551 9764 10575 9766
rect 10631 9764 10655 9766
rect 10415 9744 10711 9764
rect 10415 8732 10711 8752
rect 10471 8730 10495 8732
rect 10551 8730 10575 8732
rect 10631 8730 10655 8732
rect 10493 8678 10495 8730
rect 10557 8678 10569 8730
rect 10631 8678 10633 8730
rect 10471 8676 10495 8678
rect 10551 8676 10575 8678
rect 10631 8676 10655 8678
rect 10415 8656 10711 8676
rect 10415 7644 10711 7664
rect 10471 7642 10495 7644
rect 10551 7642 10575 7644
rect 10631 7642 10655 7644
rect 10493 7590 10495 7642
rect 10557 7590 10569 7642
rect 10631 7590 10633 7642
rect 10471 7588 10495 7590
rect 10551 7588 10575 7590
rect 10631 7588 10655 7590
rect 10415 7568 10711 7588
rect 10415 6556 10711 6576
rect 10471 6554 10495 6556
rect 10551 6554 10575 6556
rect 10631 6554 10655 6556
rect 10493 6502 10495 6554
rect 10557 6502 10569 6554
rect 10631 6502 10633 6554
rect 10471 6500 10495 6502
rect 10551 6500 10575 6502
rect 10631 6500 10655 6502
rect 10415 6480 10711 6500
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 8128 4758 8156 5306
rect 10244 5030 10272 5510
rect 10415 5468 10711 5488
rect 10471 5466 10495 5468
rect 10551 5466 10575 5468
rect 10631 5466 10655 5468
rect 10493 5414 10495 5466
rect 10557 5414 10569 5466
rect 10631 5414 10633 5466
rect 10471 5412 10495 5414
rect 10551 5412 10575 5414
rect 10631 5412 10655 5414
rect 10415 5392 10711 5412
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 8036 3942 8064 4694
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 9692 4214 9720 4558
rect 10415 4380 10711 4400
rect 10471 4378 10495 4380
rect 10551 4378 10575 4380
rect 10631 4378 10655 4380
rect 10493 4326 10495 4378
rect 10557 4326 10569 4378
rect 10631 4326 10633 4378
rect 10471 4324 10495 4326
rect 10551 4324 10575 4326
rect 10631 4324 10655 4326
rect 10415 4304 10711 4324
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 10796 4146 10824 4558
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7262 3836 7558 3856
rect 7318 3834 7342 3836
rect 7398 3834 7422 3836
rect 7478 3834 7502 3836
rect 7340 3782 7342 3834
rect 7404 3782 7416 3834
rect 7478 3782 7480 3834
rect 7318 3780 7342 3782
rect 7398 3780 7422 3782
rect 7478 3780 7502 3782
rect 7262 3760 7558 3780
rect 7668 3670 7696 3878
rect 8036 3738 8064 3878
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 9324 3670 9352 3946
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 9312 3664 9364 3670
rect 9312 3606 9364 3612
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 7024 2854 7052 3470
rect 8036 3194 8064 3538
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 9048 3194 9076 3470
rect 10415 3292 10711 3312
rect 10471 3290 10495 3292
rect 10551 3290 10575 3292
rect 10631 3290 10655 3292
rect 10493 3238 10495 3290
rect 10557 3238 10569 3290
rect 10631 3238 10633 3290
rect 10471 3236 10495 3238
rect 10551 3236 10575 3238
rect 10631 3236 10655 3238
rect 10415 3216 10711 3236
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 10888 2922 10916 3470
rect 10876 2916 10928 2922
rect 10876 2858 10928 2864
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 7262 2748 7558 2768
rect 7318 2746 7342 2748
rect 7398 2746 7422 2748
rect 7478 2746 7502 2748
rect 7340 2694 7342 2746
rect 7404 2694 7416 2746
rect 7478 2694 7480 2746
rect 7318 2692 7342 2694
rect 7398 2692 7422 2694
rect 7478 2692 7502 2694
rect 7262 2672 7558 2692
rect 6826 82 6882 480
rect 6472 54 6882 82
rect 7760 82 7788 2790
rect 8496 2514 8524 2790
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 9496 2372 9548 2378
rect 9496 2314 9548 2320
rect 8114 82 8170 480
rect 7760 54 8170 82
rect 6826 0 6882 54
rect 8114 0 8170 54
rect 9402 82 9458 480
rect 9508 82 9536 2314
rect 9402 54 9536 82
rect 10336 82 10364 2790
rect 10888 2582 10916 2858
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 10415 2204 10711 2224
rect 10471 2202 10495 2204
rect 10551 2202 10575 2204
rect 10631 2202 10655 2204
rect 10493 2150 10495 2202
rect 10557 2150 10569 2202
rect 10631 2150 10633 2202
rect 10471 2148 10495 2150
rect 10551 2148 10575 2150
rect 10631 2148 10655 2150
rect 10415 2128 10711 2148
rect 10598 82 10654 480
rect 11072 134 11100 14758
rect 12452 14482 12480 20583
rect 13358 20596 13414 21063
rect 13358 20583 13360 20596
rect 12532 20538 12584 20544
rect 13412 20583 13414 20596
rect 14370 20583 14426 21063
rect 15382 20618 15438 21063
rect 15212 20590 15438 20618
rect 13360 20538 13412 20544
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12544 8634 12572 20538
rect 13372 20507 13400 20538
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 13569 17980 13865 18000
rect 13625 17978 13649 17980
rect 13705 17978 13729 17980
rect 13785 17978 13809 17980
rect 13647 17926 13649 17978
rect 13711 17926 13723 17978
rect 13785 17926 13787 17978
rect 13625 17924 13649 17926
rect 13705 17924 13729 17926
rect 13785 17924 13809 17926
rect 13569 17904 13865 17924
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12912 16998 12940 17682
rect 14200 17338 14228 18022
rect 14384 17882 14412 20583
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 16250 12940 16934
rect 13188 16794 13216 17002
rect 13569 16892 13865 16912
rect 13625 16890 13649 16892
rect 13705 16890 13729 16892
rect 13785 16890 13809 16892
rect 13647 16838 13649 16890
rect 13711 16838 13723 16890
rect 13785 16838 13787 16890
rect 13625 16836 13649 16838
rect 13705 16836 13729 16838
rect 13785 16836 13809 16838
rect 13569 16816 13865 16836
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13174 16552 13230 16561
rect 13174 16487 13230 16496
rect 12900 16244 12952 16250
rect 12900 16186 12952 16192
rect 13188 12782 13216 16487
rect 13648 16250 13676 16594
rect 15120 16250 15148 17138
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 13569 15804 13865 15824
rect 13625 15802 13649 15804
rect 13705 15802 13729 15804
rect 13785 15802 13809 15804
rect 13647 15750 13649 15802
rect 13711 15750 13723 15802
rect 13785 15750 13787 15802
rect 13625 15748 13649 15750
rect 13705 15748 13729 15750
rect 13785 15748 13809 15750
rect 13569 15728 13865 15748
rect 13569 14716 13865 14736
rect 13625 14714 13649 14716
rect 13705 14714 13729 14716
rect 13785 14714 13809 14716
rect 13647 14662 13649 14714
rect 13711 14662 13723 14714
rect 13785 14662 13787 14714
rect 13625 14660 13649 14662
rect 13705 14660 13729 14662
rect 13785 14660 13809 14662
rect 13569 14640 13865 14660
rect 14922 13968 14978 13977
rect 14922 13903 14978 13912
rect 13569 13628 13865 13648
rect 13625 13626 13649 13628
rect 13705 13626 13729 13628
rect 13785 13626 13809 13628
rect 13647 13574 13649 13626
rect 13711 13574 13723 13626
rect 13785 13574 13787 13626
rect 13625 13572 13649 13574
rect 13705 13572 13729 13574
rect 13785 13572 13809 13574
rect 13569 13552 13865 13572
rect 14186 12880 14242 12889
rect 14186 12815 14242 12824
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13569 12540 13865 12560
rect 13625 12538 13649 12540
rect 13705 12538 13729 12540
rect 13785 12538 13809 12540
rect 13647 12486 13649 12538
rect 13711 12486 13723 12538
rect 13785 12486 13787 12538
rect 13625 12484 13649 12486
rect 13705 12484 13729 12486
rect 13785 12484 13809 12486
rect 13569 12464 13865 12484
rect 14200 11898 14228 12815
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 13569 11452 13865 11472
rect 13625 11450 13649 11452
rect 13705 11450 13729 11452
rect 13785 11450 13809 11452
rect 13647 11398 13649 11450
rect 13711 11398 13723 11450
rect 13785 11398 13787 11450
rect 13625 11396 13649 11398
rect 13705 11396 13729 11398
rect 13785 11396 13809 11398
rect 13569 11376 13865 11396
rect 14660 10810 14688 11630
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 13569 10364 13865 10384
rect 13625 10362 13649 10364
rect 13705 10362 13729 10364
rect 13785 10362 13809 10364
rect 13647 10310 13649 10362
rect 13711 10310 13723 10362
rect 13785 10310 13787 10362
rect 13625 10308 13649 10310
rect 13705 10308 13729 10310
rect 13785 10308 13809 10310
rect 13569 10288 13865 10308
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14292 9382 14320 10066
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 13569 9276 13865 9296
rect 13625 9274 13649 9276
rect 13705 9274 13729 9276
rect 13785 9274 13809 9276
rect 13647 9222 13649 9274
rect 13711 9222 13723 9274
rect 13785 9222 13787 9274
rect 13625 9220 13649 9222
rect 13705 9220 13729 9222
rect 13785 9220 13809 9222
rect 13569 9200 13865 9220
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 13096 8090 13124 8230
rect 13569 8188 13865 8208
rect 13625 8186 13649 8188
rect 13705 8186 13729 8188
rect 13785 8186 13809 8188
rect 13647 8134 13649 8186
rect 13711 8134 13723 8186
rect 13785 8134 13787 8186
rect 13625 8132 13649 8134
rect 13705 8132 13729 8134
rect 13785 8132 13809 8134
rect 13569 8112 13865 8132
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12084 7546 12112 7822
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12912 7410 12940 7890
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12912 6934 12940 7346
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 13569 7100 13865 7120
rect 13625 7098 13649 7100
rect 13705 7098 13729 7100
rect 13785 7098 13809 7100
rect 13647 7046 13649 7098
rect 13711 7046 13723 7098
rect 13785 7046 13787 7098
rect 13625 7044 13649 7046
rect 13705 7044 13729 7046
rect 13785 7044 13809 7046
rect 13569 7024 13865 7044
rect 14108 7002 14136 7278
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11900 6322 11928 6734
rect 13740 6390 13768 6802
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11900 6118 11928 6258
rect 12990 6216 13046 6225
rect 12532 6180 12584 6186
rect 12990 6151 13046 6160
rect 12532 6122 12584 6128
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11900 5710 11928 6054
rect 12544 5914 12572 6122
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 13004 5778 13032 6151
rect 13569 6012 13865 6032
rect 13625 6010 13649 6012
rect 13705 6010 13729 6012
rect 13785 6010 13809 6012
rect 13647 5958 13649 6010
rect 13711 5958 13723 6010
rect 13785 5958 13787 6010
rect 13625 5956 13649 5958
rect 13705 5956 13729 5958
rect 13785 5956 13809 5958
rect 13569 5936 13865 5956
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11440 5370 11468 5646
rect 13004 5370 13032 5714
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11624 4010 11652 4966
rect 13569 4924 13865 4944
rect 13625 4922 13649 4924
rect 13705 4922 13729 4924
rect 13785 4922 13809 4924
rect 13647 4870 13649 4922
rect 13711 4870 13723 4922
rect 13785 4870 13787 4922
rect 13625 4868 13649 4870
rect 13705 4868 13729 4870
rect 13785 4868 13809 4870
rect 13569 4848 13865 4868
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 11612 4004 11664 4010
rect 11612 3946 11664 3952
rect 11624 3534 11652 3946
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11348 3194 11376 3470
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11348 2360 11376 3130
rect 12360 2650 12388 4422
rect 13280 3942 13308 4626
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 12452 3194 12480 3878
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 11428 2372 11480 2378
rect 11348 2332 11428 2360
rect 11428 2314 11480 2320
rect 10336 54 10654 82
rect 11060 128 11112 134
rect 11060 70 11112 76
rect 11886 128 11942 480
rect 11886 76 11888 128
rect 11940 76 11942 128
rect 9402 0 9458 54
rect 10598 0 10654 54
rect 11886 0 11942 76
rect 13174 82 13230 480
rect 13280 82 13308 3878
rect 13569 3836 13865 3856
rect 13625 3834 13649 3836
rect 13705 3834 13729 3836
rect 13785 3834 13809 3836
rect 13647 3782 13649 3834
rect 13711 3782 13723 3834
rect 13785 3782 13787 3834
rect 13625 3780 13649 3782
rect 13705 3780 13729 3782
rect 13785 3780 13809 3782
rect 13569 3760 13865 3780
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13924 2854 13952 3538
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14200 3058 14228 3334
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13569 2748 13865 2768
rect 13625 2746 13649 2748
rect 13705 2746 13729 2748
rect 13785 2746 13809 2748
rect 13647 2694 13649 2746
rect 13711 2694 13723 2746
rect 13785 2694 13787 2746
rect 13625 2692 13649 2694
rect 13705 2692 13729 2694
rect 13785 2692 13809 2694
rect 13569 2672 13865 2692
rect 14200 2650 14228 2994
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13464 2378 13492 2518
rect 13452 2372 13504 2378
rect 13452 2314 13504 2320
rect 14292 1873 14320 9318
rect 14936 4078 14964 13903
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15120 12374 15148 12582
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15120 11898 15148 12310
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15212 7546 15240 20590
rect 15382 20583 15438 20590
rect 16394 20583 16450 21063
rect 17406 20583 17462 21063
rect 18418 20584 18474 21063
rect 18340 20583 18474 20584
rect 16408 19718 16436 20583
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 15304 12753 15332 19654
rect 16722 18524 17018 18544
rect 16778 18522 16802 18524
rect 16858 18522 16882 18524
rect 16938 18522 16962 18524
rect 16800 18470 16802 18522
rect 16864 18470 16876 18522
rect 16938 18470 16940 18522
rect 16778 18468 16802 18470
rect 16858 18468 16882 18470
rect 16938 18468 16962 18470
rect 16722 18448 17018 18468
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15396 16726 15424 17614
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16224 17338 16252 17478
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16224 17134 16252 17274
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16316 16998 16344 17682
rect 16722 17436 17018 17456
rect 16778 17434 16802 17436
rect 16858 17434 16882 17436
rect 16938 17434 16962 17436
rect 16800 17382 16802 17434
rect 16864 17382 16876 17434
rect 16938 17382 16940 17434
rect 16778 17380 16802 17382
rect 16858 17380 16882 17382
rect 16938 17380 16962 17382
rect 16722 17360 17018 17380
rect 17420 17338 17448 20583
rect 18340 20556 18460 20583
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 15384 16720 15436 16726
rect 15384 16662 15436 16668
rect 15396 16250 15424 16662
rect 16316 16522 16344 16934
rect 18340 16794 18368 20556
rect 18418 19680 18474 19689
rect 18418 19615 18474 19624
rect 18432 18154 18460 19615
rect 18420 18148 18472 18154
rect 18420 18090 18472 18096
rect 18418 17096 18474 17105
rect 18418 17031 18474 17040
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 16316 16182 16344 16458
rect 16722 16348 17018 16368
rect 16778 16346 16802 16348
rect 16858 16346 16882 16348
rect 16938 16346 16962 16348
rect 16800 16294 16802 16346
rect 16864 16294 16876 16346
rect 16938 16294 16940 16346
rect 16778 16292 16802 16294
rect 16858 16292 16882 16294
rect 16938 16292 16962 16294
rect 16722 16272 17018 16292
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16132 15502 16160 16050
rect 18432 16017 18460 17031
rect 18418 16008 18474 16017
rect 18418 15943 18474 15952
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 15856 15162 15884 15438
rect 16722 15260 17018 15280
rect 16778 15258 16802 15260
rect 16858 15258 16882 15260
rect 16938 15258 16962 15260
rect 16800 15206 16802 15258
rect 16864 15206 16876 15258
rect 16938 15206 16940 15258
rect 16778 15204 16802 15206
rect 16858 15204 16882 15206
rect 16938 15204 16962 15206
rect 16722 15184 17018 15204
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16224 12986 16252 13330
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 15290 12744 15346 12753
rect 15290 12679 15346 12688
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15304 11898 15332 12582
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15764 11286 15792 12174
rect 16224 11762 16252 12922
rect 16316 12782 16344 13126
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15764 10742 15792 11222
rect 16224 11150 16252 11698
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15580 10266 15608 10406
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15396 9722 15424 9998
rect 15948 9994 15976 10610
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15948 9586 15976 9930
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 15580 8906 15608 9386
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 16040 8634 16068 8910
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16316 7886 16344 8910
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16040 7546 16068 7822
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16500 4185 16528 14758
rect 16722 14172 17018 14192
rect 16778 14170 16802 14172
rect 16858 14170 16882 14172
rect 16938 14170 16962 14172
rect 16800 14118 16802 14170
rect 16864 14118 16876 14170
rect 16938 14118 16940 14170
rect 16778 14116 16802 14118
rect 16858 14116 16882 14118
rect 16938 14116 16962 14118
rect 16722 14096 17018 14116
rect 16722 13084 17018 13104
rect 16778 13082 16802 13084
rect 16858 13082 16882 13084
rect 16938 13082 16962 13084
rect 16800 13030 16802 13082
rect 16864 13030 16876 13082
rect 16938 13030 16940 13082
rect 16778 13028 16802 13030
rect 16858 13028 16882 13030
rect 16938 13028 16962 13030
rect 16722 13008 17018 13028
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 16722 11996 17018 12016
rect 16778 11994 16802 11996
rect 16858 11994 16882 11996
rect 16938 11994 16962 11996
rect 16800 11942 16802 11994
rect 16864 11942 16876 11994
rect 16938 11942 16940 11994
rect 16778 11940 16802 11942
rect 16858 11940 16882 11942
rect 16938 11940 16962 11942
rect 16722 11920 17018 11940
rect 18432 11801 18460 12854
rect 18418 11792 18474 11801
rect 18418 11727 18474 11736
rect 16722 10908 17018 10928
rect 16778 10906 16802 10908
rect 16858 10906 16882 10908
rect 16938 10906 16962 10908
rect 16800 10854 16802 10906
rect 16864 10854 16876 10906
rect 16938 10854 16940 10906
rect 16778 10852 16802 10854
rect 16858 10852 16882 10854
rect 16938 10852 16962 10854
rect 16722 10832 17018 10852
rect 16722 9820 17018 9840
rect 16778 9818 16802 9820
rect 16858 9818 16882 9820
rect 16938 9818 16962 9820
rect 16800 9766 16802 9818
rect 16864 9766 16876 9818
rect 16938 9766 16940 9818
rect 16778 9764 16802 9766
rect 16858 9764 16882 9766
rect 16938 9764 16962 9766
rect 16722 9744 17018 9764
rect 17038 8936 17094 8945
rect 17038 8871 17094 8880
rect 16722 8732 17018 8752
rect 16778 8730 16802 8732
rect 16858 8730 16882 8732
rect 16938 8730 16962 8732
rect 16800 8678 16802 8730
rect 16864 8678 16876 8730
rect 16938 8678 16940 8730
rect 16778 8676 16802 8678
rect 16858 8676 16882 8678
rect 16938 8676 16962 8678
rect 16722 8656 17018 8676
rect 17052 8634 17080 8871
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 16722 7644 17018 7664
rect 16778 7642 16802 7644
rect 16858 7642 16882 7644
rect 16938 7642 16962 7644
rect 16800 7590 16802 7642
rect 16864 7590 16876 7642
rect 16938 7590 16940 7642
rect 16778 7588 16802 7590
rect 16858 7588 16882 7590
rect 16938 7588 16962 7590
rect 16722 7568 17018 7588
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 16722 6556 17018 6576
rect 16778 6554 16802 6556
rect 16858 6554 16882 6556
rect 16938 6554 16962 6556
rect 16800 6502 16802 6554
rect 16864 6502 16876 6554
rect 16938 6502 16940 6554
rect 16778 6500 16802 6502
rect 16858 6500 16882 6502
rect 16938 6500 16962 6502
rect 16722 6480 17018 6500
rect 16722 5468 17018 5488
rect 16778 5466 16802 5468
rect 16858 5466 16882 5468
rect 16938 5466 16962 5468
rect 16800 5414 16802 5466
rect 16864 5414 16876 5466
rect 16938 5414 16940 5466
rect 16778 5412 16802 5414
rect 16858 5412 16882 5414
rect 16938 5412 16962 5414
rect 16722 5392 17018 5412
rect 16722 4380 17018 4400
rect 16778 4378 16802 4380
rect 16858 4378 16882 4380
rect 16938 4378 16962 4380
rect 16800 4326 16802 4378
rect 16864 4326 16876 4378
rect 16938 4326 16940 4378
rect 16778 4324 16802 4326
rect 16858 4324 16882 4326
rect 16938 4324 16962 4326
rect 16722 4304 17018 4324
rect 16486 4176 16542 4185
rect 16486 4111 16542 4120
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 15396 3670 15424 3878
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 15396 3194 15424 3606
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14278 1864 14334 1873
rect 14278 1799 14334 1808
rect 13174 54 13308 82
rect 14462 82 14518 480
rect 14568 82 14596 2790
rect 15672 2446 15700 3878
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15764 3194 15792 3470
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15764 3058 15792 3130
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 14462 54 14596 82
rect 15396 82 15424 2314
rect 15658 82 15714 480
rect 15396 54 15714 82
rect 16592 82 16620 3878
rect 16722 3292 17018 3312
rect 16778 3290 16802 3292
rect 16858 3290 16882 3292
rect 16938 3290 16962 3292
rect 16800 3238 16802 3290
rect 16864 3238 16876 3290
rect 16938 3238 16940 3290
rect 16778 3236 16802 3238
rect 16858 3236 16882 3238
rect 16938 3236 16962 3238
rect 16722 3216 17018 3236
rect 16722 2204 17018 2224
rect 16778 2202 16802 2204
rect 16858 2202 16882 2204
rect 16938 2202 16962 2204
rect 16800 2150 16802 2202
rect 16864 2150 16876 2202
rect 16938 2150 16940 2202
rect 16778 2148 16802 2150
rect 16858 2148 16882 2150
rect 16938 2148 16962 2150
rect 16722 2128 17018 2148
rect 16946 82 17002 480
rect 16592 54 17002 82
rect 17880 82 17908 7142
rect 18234 82 18290 480
rect 17880 54 18290 82
rect 13174 0 13230 54
rect 14462 0 14518 54
rect 15658 0 15714 54
rect 16946 0 17002 54
rect 18234 0 18290 54
<< via2 >>
rect 18 20440 74 20496
rect 1582 17856 1638 17912
rect 1490 16768 1546 16824
rect 110 16224 166 16280
rect 1122 14592 1178 14648
rect 110 14048 166 14104
rect 110 12008 166 12064
rect 110 9832 166 9888
rect 1674 17720 1730 17776
rect 4109 18522 4165 18524
rect 4189 18522 4245 18524
rect 4269 18522 4325 18524
rect 4349 18522 4405 18524
rect 4109 18470 4135 18522
rect 4135 18470 4165 18522
rect 4189 18470 4199 18522
rect 4199 18470 4245 18522
rect 4269 18470 4315 18522
rect 4315 18470 4325 18522
rect 4349 18470 4379 18522
rect 4379 18470 4405 18522
rect 4109 18468 4165 18470
rect 4189 18468 4245 18470
rect 4269 18468 4325 18470
rect 4349 18468 4405 18470
rect 3422 16496 3478 16552
rect 4986 18672 5042 18728
rect 4109 17434 4165 17436
rect 4189 17434 4245 17436
rect 4269 17434 4325 17436
rect 4349 17434 4405 17436
rect 4109 17382 4135 17434
rect 4135 17382 4165 17434
rect 4189 17382 4199 17434
rect 4199 17382 4245 17434
rect 4269 17382 4315 17434
rect 4315 17382 4325 17434
rect 4349 17382 4379 17434
rect 4379 17382 4405 17434
rect 4109 17380 4165 17382
rect 4189 17380 4245 17382
rect 4269 17380 4325 17382
rect 4349 17380 4405 17382
rect 4109 16346 4165 16348
rect 4189 16346 4245 16348
rect 4269 16346 4325 16348
rect 4349 16346 4405 16348
rect 4109 16294 4135 16346
rect 4135 16294 4165 16346
rect 4189 16294 4199 16346
rect 4199 16294 4245 16346
rect 4269 16294 4315 16346
rect 4315 16294 4325 16346
rect 4349 16294 4379 16346
rect 4379 16294 4405 16346
rect 4109 16292 4165 16294
rect 4189 16292 4245 16294
rect 4269 16292 4325 16294
rect 4349 16292 4405 16294
rect 4109 15258 4165 15260
rect 4189 15258 4245 15260
rect 4269 15258 4325 15260
rect 4349 15258 4405 15260
rect 4109 15206 4135 15258
rect 4135 15206 4165 15258
rect 4189 15206 4199 15258
rect 4199 15206 4245 15258
rect 4269 15206 4315 15258
rect 4315 15206 4325 15258
rect 4349 15206 4379 15258
rect 4379 15206 4405 15258
rect 4109 15204 4165 15206
rect 4189 15204 4245 15206
rect 4269 15204 4325 15206
rect 4349 15204 4405 15206
rect 4109 14170 4165 14172
rect 4189 14170 4245 14172
rect 4269 14170 4325 14172
rect 4349 14170 4405 14172
rect 4109 14118 4135 14170
rect 4135 14118 4165 14170
rect 4189 14118 4199 14170
rect 4199 14118 4245 14170
rect 4269 14118 4315 14170
rect 4315 14118 4325 14170
rect 4349 14118 4379 14170
rect 4379 14118 4405 14170
rect 4109 14116 4165 14118
rect 4189 14116 4245 14118
rect 4269 14116 4325 14118
rect 4349 14116 4405 14118
rect 7262 17978 7318 17980
rect 7342 17978 7398 17980
rect 7422 17978 7478 17980
rect 7502 17978 7558 17980
rect 7262 17926 7288 17978
rect 7288 17926 7318 17978
rect 7342 17926 7352 17978
rect 7352 17926 7398 17978
rect 7422 17926 7468 17978
rect 7468 17926 7478 17978
rect 7502 17926 7532 17978
rect 7532 17926 7558 17978
rect 7262 17924 7318 17926
rect 7342 17924 7398 17926
rect 7422 17924 7478 17926
rect 7502 17924 7558 17926
rect 7262 16890 7318 16892
rect 7342 16890 7398 16892
rect 7422 16890 7478 16892
rect 7502 16890 7558 16892
rect 7262 16838 7288 16890
rect 7288 16838 7318 16890
rect 7342 16838 7352 16890
rect 7352 16838 7398 16890
rect 7422 16838 7468 16890
rect 7468 16838 7478 16890
rect 7502 16838 7532 16890
rect 7532 16838 7558 16890
rect 7262 16836 7318 16838
rect 7342 16836 7398 16838
rect 7422 16836 7478 16838
rect 7502 16836 7558 16838
rect 7262 15802 7318 15804
rect 7342 15802 7398 15804
rect 7422 15802 7478 15804
rect 7502 15802 7558 15804
rect 7262 15750 7288 15802
rect 7288 15750 7318 15802
rect 7342 15750 7352 15802
rect 7352 15750 7398 15802
rect 7422 15750 7468 15802
rect 7468 15750 7478 15802
rect 7502 15750 7532 15802
rect 7532 15750 7558 15802
rect 7262 15748 7318 15750
rect 7342 15748 7398 15750
rect 7422 15748 7478 15750
rect 7502 15748 7558 15750
rect 7262 14714 7318 14716
rect 7342 14714 7398 14716
rect 7422 14714 7478 14716
rect 7502 14714 7558 14716
rect 7262 14662 7288 14714
rect 7288 14662 7318 14714
rect 7342 14662 7352 14714
rect 7352 14662 7398 14714
rect 7422 14662 7468 14714
rect 7468 14662 7478 14714
rect 7502 14662 7532 14714
rect 7532 14662 7558 14714
rect 7262 14660 7318 14662
rect 7342 14660 7398 14662
rect 7422 14660 7478 14662
rect 7502 14660 7558 14662
rect 7262 13626 7318 13628
rect 7342 13626 7398 13628
rect 7422 13626 7478 13628
rect 7502 13626 7558 13628
rect 7262 13574 7288 13626
rect 7288 13574 7318 13626
rect 7342 13574 7352 13626
rect 7352 13574 7398 13626
rect 7422 13574 7468 13626
rect 7468 13574 7478 13626
rect 7502 13574 7532 13626
rect 7532 13574 7558 13626
rect 7262 13572 7318 13574
rect 7342 13572 7398 13574
rect 7422 13572 7478 13574
rect 7502 13572 7558 13574
rect 1858 8336 1914 8392
rect 1674 6296 1730 6352
rect 110 5616 166 5672
rect 4109 13082 4165 13084
rect 4189 13082 4245 13084
rect 4269 13082 4325 13084
rect 4349 13082 4405 13084
rect 4109 13030 4135 13082
rect 4135 13030 4165 13082
rect 4189 13030 4199 13082
rect 4199 13030 4245 13082
rect 4269 13030 4315 13082
rect 4315 13030 4325 13082
rect 4349 13030 4379 13082
rect 4379 13030 4405 13082
rect 4109 13028 4165 13030
rect 4189 13028 4245 13030
rect 4269 13028 4325 13030
rect 4349 13028 4405 13030
rect 5262 12688 5318 12744
rect 7262 12538 7318 12540
rect 7342 12538 7398 12540
rect 7422 12538 7478 12540
rect 7502 12538 7558 12540
rect 7262 12486 7288 12538
rect 7288 12486 7318 12538
rect 7342 12486 7352 12538
rect 7352 12486 7398 12538
rect 7422 12486 7468 12538
rect 7468 12486 7478 12538
rect 7502 12486 7532 12538
rect 7532 12486 7558 12538
rect 7262 12484 7318 12486
rect 7342 12484 7398 12486
rect 7422 12484 7478 12486
rect 7502 12484 7558 12486
rect 4109 11994 4165 11996
rect 4189 11994 4245 11996
rect 4269 11994 4325 11996
rect 4349 11994 4405 11996
rect 4109 11942 4135 11994
rect 4135 11942 4165 11994
rect 4189 11942 4199 11994
rect 4199 11942 4245 11994
rect 4269 11942 4315 11994
rect 4315 11942 4325 11994
rect 4349 11942 4379 11994
rect 4379 11942 4405 11994
rect 4109 11940 4165 11942
rect 4189 11940 4245 11942
rect 4269 11940 4325 11942
rect 4349 11940 4405 11942
rect 7262 11450 7318 11452
rect 7342 11450 7398 11452
rect 7422 11450 7478 11452
rect 7502 11450 7558 11452
rect 7262 11398 7288 11450
rect 7288 11398 7318 11450
rect 7342 11398 7352 11450
rect 7352 11398 7398 11450
rect 7422 11398 7468 11450
rect 7468 11398 7478 11450
rect 7502 11398 7532 11450
rect 7532 11398 7558 11450
rect 7262 11396 7318 11398
rect 7342 11396 7398 11398
rect 7422 11396 7478 11398
rect 7502 11396 7558 11398
rect 4109 10906 4165 10908
rect 4189 10906 4245 10908
rect 4269 10906 4325 10908
rect 4349 10906 4405 10908
rect 4109 10854 4135 10906
rect 4135 10854 4165 10906
rect 4189 10854 4199 10906
rect 4199 10854 4245 10906
rect 4269 10854 4315 10906
rect 4315 10854 4325 10906
rect 4349 10854 4379 10906
rect 4379 10854 4405 10906
rect 4109 10852 4165 10854
rect 4189 10852 4245 10854
rect 4269 10852 4325 10854
rect 4349 10852 4405 10854
rect 5170 10648 5226 10704
rect 7262 10362 7318 10364
rect 7342 10362 7398 10364
rect 7422 10362 7478 10364
rect 7502 10362 7558 10364
rect 7262 10310 7288 10362
rect 7288 10310 7318 10362
rect 7342 10310 7352 10362
rect 7352 10310 7398 10362
rect 7422 10310 7468 10362
rect 7468 10310 7478 10362
rect 7502 10310 7532 10362
rect 7532 10310 7558 10362
rect 7262 10308 7318 10310
rect 7342 10308 7398 10310
rect 7422 10308 7478 10310
rect 7502 10308 7558 10310
rect 4109 9818 4165 9820
rect 4189 9818 4245 9820
rect 4269 9818 4325 9820
rect 4349 9818 4405 9820
rect 4109 9766 4135 9818
rect 4135 9766 4165 9818
rect 4189 9766 4199 9818
rect 4199 9766 4245 9818
rect 4269 9766 4315 9818
rect 4315 9766 4325 9818
rect 4349 9766 4379 9818
rect 4379 9766 4405 9818
rect 4109 9764 4165 9766
rect 4189 9764 4245 9766
rect 4269 9764 4325 9766
rect 4349 9764 4405 9766
rect 7262 9274 7318 9276
rect 7342 9274 7398 9276
rect 7422 9274 7478 9276
rect 7502 9274 7558 9276
rect 7262 9222 7288 9274
rect 7288 9222 7318 9274
rect 7342 9222 7352 9274
rect 7352 9222 7398 9274
rect 7422 9222 7468 9274
rect 7468 9222 7478 9274
rect 7502 9222 7532 9274
rect 7532 9222 7558 9274
rect 7262 9220 7318 9222
rect 7342 9220 7398 9222
rect 7422 9220 7478 9222
rect 7502 9220 7558 9222
rect 4109 8730 4165 8732
rect 4189 8730 4245 8732
rect 4269 8730 4325 8732
rect 4349 8730 4405 8732
rect 4109 8678 4135 8730
rect 4135 8678 4165 8730
rect 4189 8678 4199 8730
rect 4199 8678 4245 8730
rect 4269 8678 4315 8730
rect 4315 8678 4325 8730
rect 4349 8678 4379 8730
rect 4379 8678 4405 8730
rect 4109 8676 4165 8678
rect 4189 8676 4245 8678
rect 4269 8676 4325 8678
rect 4349 8676 4405 8678
rect 3974 8472 4030 8528
rect 7262 8186 7318 8188
rect 7342 8186 7398 8188
rect 7422 8186 7478 8188
rect 7502 8186 7558 8188
rect 7262 8134 7288 8186
rect 7288 8134 7318 8186
rect 7342 8134 7352 8186
rect 7352 8134 7398 8186
rect 7422 8134 7468 8186
rect 7468 8134 7478 8186
rect 7502 8134 7532 8186
rect 7532 8134 7558 8186
rect 7262 8132 7318 8134
rect 7342 8132 7398 8134
rect 7422 8132 7478 8134
rect 7502 8132 7558 8134
rect 4109 7642 4165 7644
rect 4189 7642 4245 7644
rect 4269 7642 4325 7644
rect 4349 7642 4405 7644
rect 4109 7590 4135 7642
rect 4135 7590 4165 7642
rect 4189 7590 4199 7642
rect 4199 7590 4245 7642
rect 4269 7590 4315 7642
rect 4315 7590 4325 7642
rect 4349 7590 4379 7642
rect 4379 7590 4405 7642
rect 4109 7588 4165 7590
rect 4189 7588 4245 7590
rect 4269 7588 4325 7590
rect 4349 7588 4405 7590
rect 7262 7098 7318 7100
rect 7342 7098 7398 7100
rect 7422 7098 7478 7100
rect 7502 7098 7558 7100
rect 7262 7046 7288 7098
rect 7288 7046 7318 7098
rect 7342 7046 7352 7098
rect 7352 7046 7398 7098
rect 7422 7046 7468 7098
rect 7468 7046 7478 7098
rect 7502 7046 7532 7098
rect 7532 7046 7558 7098
rect 7262 7044 7318 7046
rect 7342 7044 7398 7046
rect 7422 7044 7478 7046
rect 7502 7044 7558 7046
rect 4109 6554 4165 6556
rect 4189 6554 4245 6556
rect 4269 6554 4325 6556
rect 4349 6554 4405 6556
rect 4109 6502 4135 6554
rect 4135 6502 4165 6554
rect 4189 6502 4199 6554
rect 4199 6502 4245 6554
rect 4269 6502 4315 6554
rect 4315 6502 4325 6554
rect 4349 6502 4379 6554
rect 4379 6502 4405 6554
rect 4109 6500 4165 6502
rect 4189 6500 4245 6502
rect 4269 6500 4325 6502
rect 4349 6500 4405 6502
rect 4109 5466 4165 5468
rect 4189 5466 4245 5468
rect 4269 5466 4325 5468
rect 4349 5466 4405 5468
rect 4109 5414 4135 5466
rect 4135 5414 4165 5466
rect 4189 5414 4199 5466
rect 4199 5414 4245 5466
rect 4269 5414 4315 5466
rect 4315 5414 4325 5466
rect 4349 5414 4379 5466
rect 4379 5414 4405 5466
rect 4109 5412 4165 5414
rect 4189 5412 4245 5414
rect 4269 5412 4325 5414
rect 4349 5412 4405 5414
rect 2778 5208 2834 5264
rect 4109 4378 4165 4380
rect 4189 4378 4245 4380
rect 4269 4378 4325 4380
rect 4349 4378 4405 4380
rect 4109 4326 4135 4378
rect 4135 4326 4165 4378
rect 4189 4326 4199 4378
rect 4199 4326 4245 4378
rect 4269 4326 4315 4378
rect 4315 4326 4325 4378
rect 4349 4326 4379 4378
rect 4379 4326 4405 4378
rect 4109 4324 4165 4326
rect 4189 4324 4245 4326
rect 4269 4324 4325 4326
rect 4349 4324 4405 4326
rect 110 3576 166 3632
rect 4109 3290 4165 3292
rect 4189 3290 4245 3292
rect 4269 3290 4325 3292
rect 4349 3290 4405 3292
rect 4109 3238 4135 3290
rect 4135 3238 4165 3290
rect 4189 3238 4199 3290
rect 4199 3238 4245 3290
rect 4269 3238 4315 3290
rect 4315 3238 4325 3290
rect 4349 3238 4379 3290
rect 4379 3238 4405 3290
rect 4109 3236 4165 3238
rect 4189 3236 4245 3238
rect 4269 3236 4325 3238
rect 4349 3236 4405 3238
rect 6366 3032 6422 3088
rect 4109 2202 4165 2204
rect 4189 2202 4245 2204
rect 4269 2202 4325 2204
rect 4349 2202 4405 2204
rect 4109 2150 4135 2202
rect 4135 2150 4165 2202
rect 4189 2150 4199 2202
rect 4199 2150 4245 2202
rect 4269 2150 4315 2202
rect 4315 2150 4325 2202
rect 4349 2150 4379 2202
rect 4379 2150 4405 2202
rect 4109 2148 4165 2150
rect 4189 2148 4245 2150
rect 4269 2148 4325 2150
rect 4349 2148 4405 2150
rect 7262 6010 7318 6012
rect 7342 6010 7398 6012
rect 7422 6010 7478 6012
rect 7502 6010 7558 6012
rect 7262 5958 7288 6010
rect 7288 5958 7318 6010
rect 7342 5958 7352 6010
rect 7352 5958 7398 6010
rect 7422 5958 7468 6010
rect 7468 5958 7478 6010
rect 7502 5958 7532 6010
rect 7532 5958 7558 6010
rect 7262 5956 7318 5958
rect 7342 5956 7398 5958
rect 7422 5956 7478 5958
rect 7502 5956 7558 5958
rect 7262 4922 7318 4924
rect 7342 4922 7398 4924
rect 7422 4922 7478 4924
rect 7502 4922 7558 4924
rect 7262 4870 7288 4922
rect 7288 4870 7318 4922
rect 7342 4870 7352 4922
rect 7352 4870 7398 4922
rect 7422 4870 7468 4922
rect 7468 4870 7478 4922
rect 7502 4870 7532 4922
rect 7532 4870 7558 4922
rect 7262 4868 7318 4870
rect 7342 4868 7398 4870
rect 7422 4868 7478 4870
rect 7502 4868 7558 4870
rect 8942 15988 8944 16008
rect 8944 15988 8996 16008
rect 8996 15988 8998 16008
rect 8942 15952 8998 15988
rect 10415 18522 10471 18524
rect 10495 18522 10551 18524
rect 10575 18522 10631 18524
rect 10655 18522 10711 18524
rect 10415 18470 10441 18522
rect 10441 18470 10471 18522
rect 10495 18470 10505 18522
rect 10505 18470 10551 18522
rect 10575 18470 10621 18522
rect 10621 18470 10631 18522
rect 10655 18470 10685 18522
rect 10685 18470 10711 18522
rect 10415 18468 10471 18470
rect 10495 18468 10551 18470
rect 10575 18468 10631 18470
rect 10655 18468 10711 18470
rect 10415 17434 10471 17436
rect 10495 17434 10551 17436
rect 10575 17434 10631 17436
rect 10655 17434 10711 17436
rect 10415 17382 10441 17434
rect 10441 17382 10471 17434
rect 10495 17382 10505 17434
rect 10505 17382 10551 17434
rect 10575 17382 10621 17434
rect 10621 17382 10631 17434
rect 10655 17382 10685 17434
rect 10685 17382 10711 17434
rect 10415 17380 10471 17382
rect 10495 17380 10551 17382
rect 10575 17380 10631 17382
rect 10655 17380 10711 17382
rect 11610 17720 11666 17776
rect 10415 16346 10471 16348
rect 10495 16346 10551 16348
rect 10575 16346 10631 16348
rect 10655 16346 10711 16348
rect 10415 16294 10441 16346
rect 10441 16294 10471 16346
rect 10495 16294 10505 16346
rect 10505 16294 10551 16346
rect 10575 16294 10621 16346
rect 10621 16294 10631 16346
rect 10655 16294 10685 16346
rect 10685 16294 10711 16346
rect 10415 16292 10471 16294
rect 10495 16292 10551 16294
rect 10575 16292 10631 16294
rect 10655 16292 10711 16294
rect 10415 15258 10471 15260
rect 10495 15258 10551 15260
rect 10575 15258 10631 15260
rect 10655 15258 10711 15260
rect 10415 15206 10441 15258
rect 10441 15206 10471 15258
rect 10495 15206 10505 15258
rect 10505 15206 10551 15258
rect 10575 15206 10621 15258
rect 10621 15206 10631 15258
rect 10655 15206 10685 15258
rect 10685 15206 10711 15258
rect 10415 15204 10471 15206
rect 10495 15204 10551 15206
rect 10575 15204 10631 15206
rect 10655 15204 10711 15206
rect 10415 14170 10471 14172
rect 10495 14170 10551 14172
rect 10575 14170 10631 14172
rect 10655 14170 10711 14172
rect 10415 14118 10441 14170
rect 10441 14118 10471 14170
rect 10495 14118 10505 14170
rect 10505 14118 10551 14170
rect 10575 14118 10621 14170
rect 10621 14118 10631 14170
rect 10655 14118 10685 14170
rect 10685 14118 10711 14170
rect 10415 14116 10471 14118
rect 10495 14116 10551 14118
rect 10575 14116 10631 14118
rect 10655 14116 10711 14118
rect 10415 13082 10471 13084
rect 10495 13082 10551 13084
rect 10575 13082 10631 13084
rect 10655 13082 10711 13084
rect 10415 13030 10441 13082
rect 10441 13030 10471 13082
rect 10495 13030 10505 13082
rect 10505 13030 10551 13082
rect 10575 13030 10621 13082
rect 10621 13030 10631 13082
rect 10655 13030 10685 13082
rect 10685 13030 10711 13082
rect 10415 13028 10471 13030
rect 10495 13028 10551 13030
rect 10575 13028 10631 13030
rect 10655 13028 10711 13030
rect 10415 11994 10471 11996
rect 10495 11994 10551 11996
rect 10575 11994 10631 11996
rect 10655 11994 10711 11996
rect 10415 11942 10441 11994
rect 10441 11942 10471 11994
rect 10495 11942 10505 11994
rect 10505 11942 10551 11994
rect 10575 11942 10621 11994
rect 10621 11942 10631 11994
rect 10655 11942 10685 11994
rect 10685 11942 10711 11994
rect 10415 11940 10471 11942
rect 10495 11940 10551 11942
rect 10575 11940 10631 11942
rect 10655 11940 10711 11942
rect 10415 10906 10471 10908
rect 10495 10906 10551 10908
rect 10575 10906 10631 10908
rect 10655 10906 10711 10908
rect 10415 10854 10441 10906
rect 10441 10854 10471 10906
rect 10495 10854 10505 10906
rect 10505 10854 10551 10906
rect 10575 10854 10621 10906
rect 10621 10854 10631 10906
rect 10655 10854 10685 10906
rect 10685 10854 10711 10906
rect 10415 10852 10471 10854
rect 10495 10852 10551 10854
rect 10575 10852 10631 10854
rect 10655 10852 10711 10854
rect 10415 9818 10471 9820
rect 10495 9818 10551 9820
rect 10575 9818 10631 9820
rect 10655 9818 10711 9820
rect 10415 9766 10441 9818
rect 10441 9766 10471 9818
rect 10495 9766 10505 9818
rect 10505 9766 10551 9818
rect 10575 9766 10621 9818
rect 10621 9766 10631 9818
rect 10655 9766 10685 9818
rect 10685 9766 10711 9818
rect 10415 9764 10471 9766
rect 10495 9764 10551 9766
rect 10575 9764 10631 9766
rect 10655 9764 10711 9766
rect 10415 8730 10471 8732
rect 10495 8730 10551 8732
rect 10575 8730 10631 8732
rect 10655 8730 10711 8732
rect 10415 8678 10441 8730
rect 10441 8678 10471 8730
rect 10495 8678 10505 8730
rect 10505 8678 10551 8730
rect 10575 8678 10621 8730
rect 10621 8678 10631 8730
rect 10655 8678 10685 8730
rect 10685 8678 10711 8730
rect 10415 8676 10471 8678
rect 10495 8676 10551 8678
rect 10575 8676 10631 8678
rect 10655 8676 10711 8678
rect 10415 7642 10471 7644
rect 10495 7642 10551 7644
rect 10575 7642 10631 7644
rect 10655 7642 10711 7644
rect 10415 7590 10441 7642
rect 10441 7590 10471 7642
rect 10495 7590 10505 7642
rect 10505 7590 10551 7642
rect 10575 7590 10621 7642
rect 10621 7590 10631 7642
rect 10655 7590 10685 7642
rect 10685 7590 10711 7642
rect 10415 7588 10471 7590
rect 10495 7588 10551 7590
rect 10575 7588 10631 7590
rect 10655 7588 10711 7590
rect 10415 6554 10471 6556
rect 10495 6554 10551 6556
rect 10575 6554 10631 6556
rect 10655 6554 10711 6556
rect 10415 6502 10441 6554
rect 10441 6502 10471 6554
rect 10495 6502 10505 6554
rect 10505 6502 10551 6554
rect 10575 6502 10621 6554
rect 10621 6502 10631 6554
rect 10655 6502 10685 6554
rect 10685 6502 10711 6554
rect 10415 6500 10471 6502
rect 10495 6500 10551 6502
rect 10575 6500 10631 6502
rect 10655 6500 10711 6502
rect 10415 5466 10471 5468
rect 10495 5466 10551 5468
rect 10575 5466 10631 5468
rect 10655 5466 10711 5468
rect 10415 5414 10441 5466
rect 10441 5414 10471 5466
rect 10495 5414 10505 5466
rect 10505 5414 10551 5466
rect 10575 5414 10621 5466
rect 10621 5414 10631 5466
rect 10655 5414 10685 5466
rect 10685 5414 10711 5466
rect 10415 5412 10471 5414
rect 10495 5412 10551 5414
rect 10575 5412 10631 5414
rect 10655 5412 10711 5414
rect 10415 4378 10471 4380
rect 10495 4378 10551 4380
rect 10575 4378 10631 4380
rect 10655 4378 10711 4380
rect 10415 4326 10441 4378
rect 10441 4326 10471 4378
rect 10495 4326 10505 4378
rect 10505 4326 10551 4378
rect 10575 4326 10621 4378
rect 10621 4326 10631 4378
rect 10655 4326 10685 4378
rect 10685 4326 10711 4378
rect 10415 4324 10471 4326
rect 10495 4324 10551 4326
rect 10575 4324 10631 4326
rect 10655 4324 10711 4326
rect 7262 3834 7318 3836
rect 7342 3834 7398 3836
rect 7422 3834 7478 3836
rect 7502 3834 7558 3836
rect 7262 3782 7288 3834
rect 7288 3782 7318 3834
rect 7342 3782 7352 3834
rect 7352 3782 7398 3834
rect 7422 3782 7468 3834
rect 7468 3782 7478 3834
rect 7502 3782 7532 3834
rect 7532 3782 7558 3834
rect 7262 3780 7318 3782
rect 7342 3780 7398 3782
rect 7422 3780 7478 3782
rect 7502 3780 7558 3782
rect 10415 3290 10471 3292
rect 10495 3290 10551 3292
rect 10575 3290 10631 3292
rect 10655 3290 10711 3292
rect 10415 3238 10441 3290
rect 10441 3238 10471 3290
rect 10495 3238 10505 3290
rect 10505 3238 10551 3290
rect 10575 3238 10621 3290
rect 10621 3238 10631 3290
rect 10655 3238 10685 3290
rect 10685 3238 10711 3290
rect 10415 3236 10471 3238
rect 10495 3236 10551 3238
rect 10575 3236 10631 3238
rect 10655 3236 10711 3238
rect 7262 2746 7318 2748
rect 7342 2746 7398 2748
rect 7422 2746 7478 2748
rect 7502 2746 7558 2748
rect 7262 2694 7288 2746
rect 7288 2694 7318 2746
rect 7342 2694 7352 2746
rect 7352 2694 7398 2746
rect 7422 2694 7468 2746
rect 7468 2694 7478 2746
rect 7502 2694 7532 2746
rect 7532 2694 7558 2746
rect 7262 2692 7318 2694
rect 7342 2692 7398 2694
rect 7422 2692 7478 2694
rect 7502 2692 7558 2694
rect 10415 2202 10471 2204
rect 10495 2202 10551 2204
rect 10575 2202 10631 2204
rect 10655 2202 10711 2204
rect 10415 2150 10441 2202
rect 10441 2150 10471 2202
rect 10495 2150 10505 2202
rect 10505 2150 10551 2202
rect 10575 2150 10621 2202
rect 10621 2150 10631 2202
rect 10655 2150 10685 2202
rect 10685 2150 10711 2202
rect 10415 2148 10471 2150
rect 10495 2148 10551 2150
rect 10575 2148 10631 2150
rect 10655 2148 10711 2150
rect 13569 17978 13625 17980
rect 13649 17978 13705 17980
rect 13729 17978 13785 17980
rect 13809 17978 13865 17980
rect 13569 17926 13595 17978
rect 13595 17926 13625 17978
rect 13649 17926 13659 17978
rect 13659 17926 13705 17978
rect 13729 17926 13775 17978
rect 13775 17926 13785 17978
rect 13809 17926 13839 17978
rect 13839 17926 13865 17978
rect 13569 17924 13625 17926
rect 13649 17924 13705 17926
rect 13729 17924 13785 17926
rect 13809 17924 13865 17926
rect 13569 16890 13625 16892
rect 13649 16890 13705 16892
rect 13729 16890 13785 16892
rect 13809 16890 13865 16892
rect 13569 16838 13595 16890
rect 13595 16838 13625 16890
rect 13649 16838 13659 16890
rect 13659 16838 13705 16890
rect 13729 16838 13775 16890
rect 13775 16838 13785 16890
rect 13809 16838 13839 16890
rect 13839 16838 13865 16890
rect 13569 16836 13625 16838
rect 13649 16836 13705 16838
rect 13729 16836 13785 16838
rect 13809 16836 13865 16838
rect 13174 16496 13230 16552
rect 13569 15802 13625 15804
rect 13649 15802 13705 15804
rect 13729 15802 13785 15804
rect 13809 15802 13865 15804
rect 13569 15750 13595 15802
rect 13595 15750 13625 15802
rect 13649 15750 13659 15802
rect 13659 15750 13705 15802
rect 13729 15750 13775 15802
rect 13775 15750 13785 15802
rect 13809 15750 13839 15802
rect 13839 15750 13865 15802
rect 13569 15748 13625 15750
rect 13649 15748 13705 15750
rect 13729 15748 13785 15750
rect 13809 15748 13865 15750
rect 13569 14714 13625 14716
rect 13649 14714 13705 14716
rect 13729 14714 13785 14716
rect 13809 14714 13865 14716
rect 13569 14662 13595 14714
rect 13595 14662 13625 14714
rect 13649 14662 13659 14714
rect 13659 14662 13705 14714
rect 13729 14662 13775 14714
rect 13775 14662 13785 14714
rect 13809 14662 13839 14714
rect 13839 14662 13865 14714
rect 13569 14660 13625 14662
rect 13649 14660 13705 14662
rect 13729 14660 13785 14662
rect 13809 14660 13865 14662
rect 14922 13912 14978 13968
rect 13569 13626 13625 13628
rect 13649 13626 13705 13628
rect 13729 13626 13785 13628
rect 13809 13626 13865 13628
rect 13569 13574 13595 13626
rect 13595 13574 13625 13626
rect 13649 13574 13659 13626
rect 13659 13574 13705 13626
rect 13729 13574 13775 13626
rect 13775 13574 13785 13626
rect 13809 13574 13839 13626
rect 13839 13574 13865 13626
rect 13569 13572 13625 13574
rect 13649 13572 13705 13574
rect 13729 13572 13785 13574
rect 13809 13572 13865 13574
rect 14186 12824 14242 12880
rect 13569 12538 13625 12540
rect 13649 12538 13705 12540
rect 13729 12538 13785 12540
rect 13809 12538 13865 12540
rect 13569 12486 13595 12538
rect 13595 12486 13625 12538
rect 13649 12486 13659 12538
rect 13659 12486 13705 12538
rect 13729 12486 13775 12538
rect 13775 12486 13785 12538
rect 13809 12486 13839 12538
rect 13839 12486 13865 12538
rect 13569 12484 13625 12486
rect 13649 12484 13705 12486
rect 13729 12484 13785 12486
rect 13809 12484 13865 12486
rect 13569 11450 13625 11452
rect 13649 11450 13705 11452
rect 13729 11450 13785 11452
rect 13809 11450 13865 11452
rect 13569 11398 13595 11450
rect 13595 11398 13625 11450
rect 13649 11398 13659 11450
rect 13659 11398 13705 11450
rect 13729 11398 13775 11450
rect 13775 11398 13785 11450
rect 13809 11398 13839 11450
rect 13839 11398 13865 11450
rect 13569 11396 13625 11398
rect 13649 11396 13705 11398
rect 13729 11396 13785 11398
rect 13809 11396 13865 11398
rect 13569 10362 13625 10364
rect 13649 10362 13705 10364
rect 13729 10362 13785 10364
rect 13809 10362 13865 10364
rect 13569 10310 13595 10362
rect 13595 10310 13625 10362
rect 13649 10310 13659 10362
rect 13659 10310 13705 10362
rect 13729 10310 13775 10362
rect 13775 10310 13785 10362
rect 13809 10310 13839 10362
rect 13839 10310 13865 10362
rect 13569 10308 13625 10310
rect 13649 10308 13705 10310
rect 13729 10308 13785 10310
rect 13809 10308 13865 10310
rect 13569 9274 13625 9276
rect 13649 9274 13705 9276
rect 13729 9274 13785 9276
rect 13809 9274 13865 9276
rect 13569 9222 13595 9274
rect 13595 9222 13625 9274
rect 13649 9222 13659 9274
rect 13659 9222 13705 9274
rect 13729 9222 13775 9274
rect 13775 9222 13785 9274
rect 13809 9222 13839 9274
rect 13839 9222 13865 9274
rect 13569 9220 13625 9222
rect 13649 9220 13705 9222
rect 13729 9220 13785 9222
rect 13809 9220 13865 9222
rect 13569 8186 13625 8188
rect 13649 8186 13705 8188
rect 13729 8186 13785 8188
rect 13809 8186 13865 8188
rect 13569 8134 13595 8186
rect 13595 8134 13625 8186
rect 13649 8134 13659 8186
rect 13659 8134 13705 8186
rect 13729 8134 13775 8186
rect 13775 8134 13785 8186
rect 13809 8134 13839 8186
rect 13839 8134 13865 8186
rect 13569 8132 13625 8134
rect 13649 8132 13705 8134
rect 13729 8132 13785 8134
rect 13809 8132 13865 8134
rect 13569 7098 13625 7100
rect 13649 7098 13705 7100
rect 13729 7098 13785 7100
rect 13809 7098 13865 7100
rect 13569 7046 13595 7098
rect 13595 7046 13625 7098
rect 13649 7046 13659 7098
rect 13659 7046 13705 7098
rect 13729 7046 13775 7098
rect 13775 7046 13785 7098
rect 13809 7046 13839 7098
rect 13839 7046 13865 7098
rect 13569 7044 13625 7046
rect 13649 7044 13705 7046
rect 13729 7044 13785 7046
rect 13809 7044 13865 7046
rect 12990 6160 13046 6216
rect 13569 6010 13625 6012
rect 13649 6010 13705 6012
rect 13729 6010 13785 6012
rect 13809 6010 13865 6012
rect 13569 5958 13595 6010
rect 13595 5958 13625 6010
rect 13649 5958 13659 6010
rect 13659 5958 13705 6010
rect 13729 5958 13775 6010
rect 13775 5958 13785 6010
rect 13809 5958 13839 6010
rect 13839 5958 13865 6010
rect 13569 5956 13625 5958
rect 13649 5956 13705 5958
rect 13729 5956 13785 5958
rect 13809 5956 13865 5958
rect 13569 4922 13625 4924
rect 13649 4922 13705 4924
rect 13729 4922 13785 4924
rect 13809 4922 13865 4924
rect 13569 4870 13595 4922
rect 13595 4870 13625 4922
rect 13649 4870 13659 4922
rect 13659 4870 13705 4922
rect 13729 4870 13775 4922
rect 13775 4870 13785 4922
rect 13809 4870 13839 4922
rect 13839 4870 13865 4922
rect 13569 4868 13625 4870
rect 13649 4868 13705 4870
rect 13729 4868 13785 4870
rect 13809 4868 13865 4870
rect 13569 3834 13625 3836
rect 13649 3834 13705 3836
rect 13729 3834 13785 3836
rect 13809 3834 13865 3836
rect 13569 3782 13595 3834
rect 13595 3782 13625 3834
rect 13649 3782 13659 3834
rect 13659 3782 13705 3834
rect 13729 3782 13775 3834
rect 13775 3782 13785 3834
rect 13809 3782 13839 3834
rect 13839 3782 13865 3834
rect 13569 3780 13625 3782
rect 13649 3780 13705 3782
rect 13729 3780 13785 3782
rect 13809 3780 13865 3782
rect 13569 2746 13625 2748
rect 13649 2746 13705 2748
rect 13729 2746 13785 2748
rect 13809 2746 13865 2748
rect 13569 2694 13595 2746
rect 13595 2694 13625 2746
rect 13649 2694 13659 2746
rect 13659 2694 13705 2746
rect 13729 2694 13775 2746
rect 13775 2694 13785 2746
rect 13809 2694 13839 2746
rect 13839 2694 13865 2746
rect 13569 2692 13625 2694
rect 13649 2692 13705 2694
rect 13729 2692 13785 2694
rect 13809 2692 13865 2694
rect 16722 18522 16778 18524
rect 16802 18522 16858 18524
rect 16882 18522 16938 18524
rect 16962 18522 17018 18524
rect 16722 18470 16748 18522
rect 16748 18470 16778 18522
rect 16802 18470 16812 18522
rect 16812 18470 16858 18522
rect 16882 18470 16928 18522
rect 16928 18470 16938 18522
rect 16962 18470 16992 18522
rect 16992 18470 17018 18522
rect 16722 18468 16778 18470
rect 16802 18468 16858 18470
rect 16882 18468 16938 18470
rect 16962 18468 17018 18470
rect 16722 17434 16778 17436
rect 16802 17434 16858 17436
rect 16882 17434 16938 17436
rect 16962 17434 17018 17436
rect 16722 17382 16748 17434
rect 16748 17382 16778 17434
rect 16802 17382 16812 17434
rect 16812 17382 16858 17434
rect 16882 17382 16928 17434
rect 16928 17382 16938 17434
rect 16962 17382 16992 17434
rect 16992 17382 17018 17434
rect 16722 17380 16778 17382
rect 16802 17380 16858 17382
rect 16882 17380 16938 17382
rect 16962 17380 17018 17382
rect 18418 19624 18474 19680
rect 18418 17040 18474 17096
rect 16722 16346 16778 16348
rect 16802 16346 16858 16348
rect 16882 16346 16938 16348
rect 16962 16346 17018 16348
rect 16722 16294 16748 16346
rect 16748 16294 16778 16346
rect 16802 16294 16812 16346
rect 16812 16294 16858 16346
rect 16882 16294 16928 16346
rect 16928 16294 16938 16346
rect 16962 16294 16992 16346
rect 16992 16294 17018 16346
rect 16722 16292 16778 16294
rect 16802 16292 16858 16294
rect 16882 16292 16938 16294
rect 16962 16292 17018 16294
rect 18418 15952 18474 16008
rect 16722 15258 16778 15260
rect 16802 15258 16858 15260
rect 16882 15258 16938 15260
rect 16962 15258 17018 15260
rect 16722 15206 16748 15258
rect 16748 15206 16778 15258
rect 16802 15206 16812 15258
rect 16812 15206 16858 15258
rect 16882 15206 16928 15258
rect 16928 15206 16938 15258
rect 16962 15206 16992 15258
rect 16992 15206 17018 15258
rect 16722 15204 16778 15206
rect 16802 15204 16858 15206
rect 16882 15204 16938 15206
rect 16962 15204 17018 15206
rect 15290 12688 15346 12744
rect 16722 14170 16778 14172
rect 16802 14170 16858 14172
rect 16882 14170 16938 14172
rect 16962 14170 17018 14172
rect 16722 14118 16748 14170
rect 16748 14118 16778 14170
rect 16802 14118 16812 14170
rect 16812 14118 16858 14170
rect 16882 14118 16928 14170
rect 16928 14118 16938 14170
rect 16962 14118 16992 14170
rect 16992 14118 17018 14170
rect 16722 14116 16778 14118
rect 16802 14116 16858 14118
rect 16882 14116 16938 14118
rect 16962 14116 17018 14118
rect 16722 13082 16778 13084
rect 16802 13082 16858 13084
rect 16882 13082 16938 13084
rect 16962 13082 17018 13084
rect 16722 13030 16748 13082
rect 16748 13030 16778 13082
rect 16802 13030 16812 13082
rect 16812 13030 16858 13082
rect 16882 13030 16928 13082
rect 16928 13030 16938 13082
rect 16962 13030 16992 13082
rect 16992 13030 17018 13082
rect 16722 13028 16778 13030
rect 16802 13028 16858 13030
rect 16882 13028 16938 13030
rect 16962 13028 17018 13030
rect 16722 11994 16778 11996
rect 16802 11994 16858 11996
rect 16882 11994 16938 11996
rect 16962 11994 17018 11996
rect 16722 11942 16748 11994
rect 16748 11942 16778 11994
rect 16802 11942 16812 11994
rect 16812 11942 16858 11994
rect 16882 11942 16928 11994
rect 16928 11942 16938 11994
rect 16962 11942 16992 11994
rect 16992 11942 17018 11994
rect 16722 11940 16778 11942
rect 16802 11940 16858 11942
rect 16882 11940 16938 11942
rect 16962 11940 17018 11942
rect 18418 11736 18474 11792
rect 16722 10906 16778 10908
rect 16802 10906 16858 10908
rect 16882 10906 16938 10908
rect 16962 10906 17018 10908
rect 16722 10854 16748 10906
rect 16748 10854 16778 10906
rect 16802 10854 16812 10906
rect 16812 10854 16858 10906
rect 16882 10854 16928 10906
rect 16928 10854 16938 10906
rect 16962 10854 16992 10906
rect 16992 10854 17018 10906
rect 16722 10852 16778 10854
rect 16802 10852 16858 10854
rect 16882 10852 16938 10854
rect 16962 10852 17018 10854
rect 16722 9818 16778 9820
rect 16802 9818 16858 9820
rect 16882 9818 16938 9820
rect 16962 9818 17018 9820
rect 16722 9766 16748 9818
rect 16748 9766 16778 9818
rect 16802 9766 16812 9818
rect 16812 9766 16858 9818
rect 16882 9766 16928 9818
rect 16928 9766 16938 9818
rect 16962 9766 16992 9818
rect 16992 9766 17018 9818
rect 16722 9764 16778 9766
rect 16802 9764 16858 9766
rect 16882 9764 16938 9766
rect 16962 9764 17018 9766
rect 17038 8880 17094 8936
rect 16722 8730 16778 8732
rect 16802 8730 16858 8732
rect 16882 8730 16938 8732
rect 16962 8730 17018 8732
rect 16722 8678 16748 8730
rect 16748 8678 16778 8730
rect 16802 8678 16812 8730
rect 16812 8678 16858 8730
rect 16882 8678 16928 8730
rect 16928 8678 16938 8730
rect 16962 8678 16992 8730
rect 16992 8678 17018 8730
rect 16722 8676 16778 8678
rect 16802 8676 16858 8678
rect 16882 8676 16938 8678
rect 16962 8676 17018 8678
rect 16722 7642 16778 7644
rect 16802 7642 16858 7644
rect 16882 7642 16938 7644
rect 16962 7642 17018 7644
rect 16722 7590 16748 7642
rect 16748 7590 16778 7642
rect 16802 7590 16812 7642
rect 16812 7590 16858 7642
rect 16882 7590 16928 7642
rect 16928 7590 16938 7642
rect 16962 7590 16992 7642
rect 16992 7590 17018 7642
rect 16722 7588 16778 7590
rect 16802 7588 16858 7590
rect 16882 7588 16938 7590
rect 16962 7588 17018 7590
rect 16722 6554 16778 6556
rect 16802 6554 16858 6556
rect 16882 6554 16938 6556
rect 16962 6554 17018 6556
rect 16722 6502 16748 6554
rect 16748 6502 16778 6554
rect 16802 6502 16812 6554
rect 16812 6502 16858 6554
rect 16882 6502 16928 6554
rect 16928 6502 16938 6554
rect 16962 6502 16992 6554
rect 16992 6502 17018 6554
rect 16722 6500 16778 6502
rect 16802 6500 16858 6502
rect 16882 6500 16938 6502
rect 16962 6500 17018 6502
rect 16722 5466 16778 5468
rect 16802 5466 16858 5468
rect 16882 5466 16938 5468
rect 16962 5466 17018 5468
rect 16722 5414 16748 5466
rect 16748 5414 16778 5466
rect 16802 5414 16812 5466
rect 16812 5414 16858 5466
rect 16882 5414 16928 5466
rect 16928 5414 16938 5466
rect 16962 5414 16992 5466
rect 16992 5414 17018 5466
rect 16722 5412 16778 5414
rect 16802 5412 16858 5414
rect 16882 5412 16938 5414
rect 16962 5412 17018 5414
rect 16722 4378 16778 4380
rect 16802 4378 16858 4380
rect 16882 4378 16938 4380
rect 16962 4378 17018 4380
rect 16722 4326 16748 4378
rect 16748 4326 16778 4378
rect 16802 4326 16812 4378
rect 16812 4326 16858 4378
rect 16882 4326 16928 4378
rect 16928 4326 16938 4378
rect 16962 4326 16992 4378
rect 16992 4326 17018 4378
rect 16722 4324 16778 4326
rect 16802 4324 16858 4326
rect 16882 4324 16938 4326
rect 16962 4324 17018 4326
rect 16486 4120 16542 4176
rect 14278 1808 14334 1864
rect 16722 3290 16778 3292
rect 16802 3290 16858 3292
rect 16882 3290 16938 3292
rect 16962 3290 17018 3292
rect 16722 3238 16748 3290
rect 16748 3238 16778 3290
rect 16802 3238 16812 3290
rect 16812 3238 16858 3290
rect 16882 3238 16928 3290
rect 16928 3238 16938 3290
rect 16962 3238 16992 3290
rect 16992 3238 17018 3290
rect 16722 3236 16778 3238
rect 16802 3236 16858 3238
rect 16882 3236 16938 3238
rect 16962 3236 17018 3238
rect 16722 2202 16778 2204
rect 16802 2202 16858 2204
rect 16882 2202 16938 2204
rect 16962 2202 17018 2204
rect 16722 2150 16748 2202
rect 16748 2150 16778 2202
rect 16802 2150 16812 2202
rect 16812 2150 16858 2202
rect 16882 2150 16928 2202
rect 16928 2150 16938 2202
rect 16962 2150 16992 2202
rect 16992 2150 17018 2202
rect 16722 2148 16778 2150
rect 16802 2148 16858 2150
rect 16882 2148 16938 2150
rect 16962 2148 17018 2150
<< metal3 >>
rect 0 20496 480 20528
rect 0 20440 18 20496
rect 74 20440 480 20496
rect 0 20408 480 20440
rect 18439 19685 18919 19712
rect 18413 19682 18919 19685
rect 18332 19680 18919 19682
rect 18332 19624 18418 19680
rect 18474 19624 18919 19680
rect 18332 19622 18919 19624
rect 18413 19619 18919 19622
rect 18439 19592 18919 19619
rect 0 19320 480 19440
rect 62 18730 122 19320
rect 4981 18730 5047 18733
rect 62 18728 5047 18730
rect 62 18672 4986 18728
rect 5042 18672 5047 18728
rect 62 18670 5047 18672
rect 4981 18667 5047 18670
rect 4097 18528 4417 18529
rect 4097 18464 4105 18528
rect 4169 18464 4185 18528
rect 4249 18464 4265 18528
rect 4329 18464 4345 18528
rect 4409 18464 4417 18528
rect 4097 18463 4417 18464
rect 10403 18528 10723 18529
rect 10403 18464 10411 18528
rect 10475 18464 10491 18528
rect 10555 18464 10571 18528
rect 10635 18464 10651 18528
rect 10715 18464 10723 18528
rect 10403 18463 10723 18464
rect 16710 18528 17030 18529
rect 16710 18464 16718 18528
rect 16782 18464 16798 18528
rect 16862 18464 16878 18528
rect 16942 18464 16958 18528
rect 17022 18464 17030 18528
rect 16710 18463 17030 18464
rect 0 18232 480 18352
rect 62 17914 122 18232
rect 7250 17984 7570 17985
rect 7250 17920 7258 17984
rect 7322 17920 7338 17984
rect 7402 17920 7418 17984
rect 7482 17920 7498 17984
rect 7562 17920 7570 17984
rect 7250 17919 7570 17920
rect 13557 17984 13877 17985
rect 13557 17920 13565 17984
rect 13629 17920 13645 17984
rect 13709 17920 13725 17984
rect 13789 17920 13805 17984
rect 13869 17920 13877 17984
rect 13557 17919 13877 17920
rect 1577 17914 1643 17917
rect 62 17912 1643 17914
rect 62 17856 1582 17912
rect 1638 17856 1643 17912
rect 62 17854 1643 17856
rect 1577 17851 1643 17854
rect 1669 17778 1735 17781
rect 11605 17778 11671 17781
rect 1669 17776 11671 17778
rect 1669 17720 1674 17776
rect 1730 17720 11610 17776
rect 11666 17720 11671 17776
rect 1669 17718 11671 17720
rect 1669 17715 1735 17718
rect 11605 17715 11671 17718
rect 4097 17440 4417 17441
rect 0 17280 480 17400
rect 4097 17376 4105 17440
rect 4169 17376 4185 17440
rect 4249 17376 4265 17440
rect 4329 17376 4345 17440
rect 4409 17376 4417 17440
rect 4097 17375 4417 17376
rect 10403 17440 10723 17441
rect 10403 17376 10411 17440
rect 10475 17376 10491 17440
rect 10555 17376 10571 17440
rect 10635 17376 10651 17440
rect 10715 17376 10723 17440
rect 10403 17375 10723 17376
rect 16710 17440 17030 17441
rect 16710 17376 16718 17440
rect 16782 17376 16798 17440
rect 16862 17376 16878 17440
rect 16942 17376 16958 17440
rect 17022 17376 17030 17440
rect 16710 17375 17030 17376
rect 62 16826 122 17280
rect 18439 17101 18919 17128
rect 18413 17098 18919 17101
rect 18332 17096 18919 17098
rect 18332 17040 18418 17096
rect 18474 17040 18919 17096
rect 18332 17038 18919 17040
rect 18413 17035 18919 17038
rect 18439 17008 18919 17035
rect 7250 16896 7570 16897
rect 7250 16832 7258 16896
rect 7322 16832 7338 16896
rect 7402 16832 7418 16896
rect 7482 16832 7498 16896
rect 7562 16832 7570 16896
rect 7250 16831 7570 16832
rect 13557 16896 13877 16897
rect 13557 16832 13565 16896
rect 13629 16832 13645 16896
rect 13709 16832 13725 16896
rect 13789 16832 13805 16896
rect 13869 16832 13877 16896
rect 13557 16831 13877 16832
rect 1485 16826 1551 16829
rect 62 16824 1551 16826
rect 62 16768 1490 16824
rect 1546 16768 1551 16824
rect 62 16766 1551 16768
rect 1485 16763 1551 16766
rect 3417 16554 3483 16557
rect 13169 16554 13235 16557
rect 3417 16552 13235 16554
rect 3417 16496 3422 16552
rect 3478 16496 13174 16552
rect 13230 16496 13235 16552
rect 3417 16494 13235 16496
rect 3417 16491 3483 16494
rect 13169 16491 13235 16494
rect 4097 16352 4417 16353
rect 0 16280 480 16312
rect 4097 16288 4105 16352
rect 4169 16288 4185 16352
rect 4249 16288 4265 16352
rect 4329 16288 4345 16352
rect 4409 16288 4417 16352
rect 4097 16287 4417 16288
rect 10403 16352 10723 16353
rect 10403 16288 10411 16352
rect 10475 16288 10491 16352
rect 10555 16288 10571 16352
rect 10635 16288 10651 16352
rect 10715 16288 10723 16352
rect 10403 16287 10723 16288
rect 16710 16352 17030 16353
rect 16710 16288 16718 16352
rect 16782 16288 16798 16352
rect 16862 16288 16878 16352
rect 16942 16288 16958 16352
rect 17022 16288 17030 16352
rect 16710 16287 17030 16288
rect 0 16224 110 16280
rect 166 16224 480 16280
rect 0 16192 480 16224
rect 8937 16010 9003 16013
rect 18413 16010 18479 16013
rect 8937 16008 18479 16010
rect 8937 15952 8942 16008
rect 8998 15952 18418 16008
rect 18474 15952 18479 16008
rect 8937 15950 18479 15952
rect 8937 15947 9003 15950
rect 18413 15947 18479 15950
rect 7250 15808 7570 15809
rect 7250 15744 7258 15808
rect 7322 15744 7338 15808
rect 7402 15744 7418 15808
rect 7482 15744 7498 15808
rect 7562 15744 7570 15808
rect 7250 15743 7570 15744
rect 13557 15808 13877 15809
rect 13557 15744 13565 15808
rect 13629 15744 13645 15808
rect 13709 15744 13725 15808
rect 13789 15744 13805 15808
rect 13869 15744 13877 15808
rect 13557 15743 13877 15744
rect 4097 15264 4417 15265
rect 0 15104 480 15224
rect 4097 15200 4105 15264
rect 4169 15200 4185 15264
rect 4249 15200 4265 15264
rect 4329 15200 4345 15264
rect 4409 15200 4417 15264
rect 4097 15199 4417 15200
rect 10403 15264 10723 15265
rect 10403 15200 10411 15264
rect 10475 15200 10491 15264
rect 10555 15200 10571 15264
rect 10635 15200 10651 15264
rect 10715 15200 10723 15264
rect 10403 15199 10723 15200
rect 16710 15264 17030 15265
rect 16710 15200 16718 15264
rect 16782 15200 16798 15264
rect 16862 15200 16878 15264
rect 16942 15200 16958 15264
rect 17022 15200 17030 15264
rect 16710 15199 17030 15200
rect 62 14650 122 15104
rect 7250 14720 7570 14721
rect 7250 14656 7258 14720
rect 7322 14656 7338 14720
rect 7402 14656 7418 14720
rect 7482 14656 7498 14720
rect 7562 14656 7570 14720
rect 7250 14655 7570 14656
rect 13557 14720 13877 14721
rect 13557 14656 13565 14720
rect 13629 14656 13645 14720
rect 13709 14656 13725 14720
rect 13789 14656 13805 14720
rect 13869 14656 13877 14720
rect 13557 14655 13877 14656
rect 1117 14650 1183 14653
rect 62 14648 1183 14650
rect 62 14592 1122 14648
rect 1178 14592 1183 14648
rect 62 14590 1183 14592
rect 1117 14587 1183 14590
rect 18439 14288 18919 14408
rect 4097 14176 4417 14177
rect 0 14104 480 14136
rect 4097 14112 4105 14176
rect 4169 14112 4185 14176
rect 4249 14112 4265 14176
rect 4329 14112 4345 14176
rect 4409 14112 4417 14176
rect 4097 14111 4417 14112
rect 10403 14176 10723 14177
rect 10403 14112 10411 14176
rect 10475 14112 10491 14176
rect 10555 14112 10571 14176
rect 10635 14112 10651 14176
rect 10715 14112 10723 14176
rect 10403 14111 10723 14112
rect 16710 14176 17030 14177
rect 16710 14112 16718 14176
rect 16782 14112 16798 14176
rect 16862 14112 16878 14176
rect 16942 14112 16958 14176
rect 17022 14112 17030 14176
rect 16710 14111 17030 14112
rect 0 14048 110 14104
rect 166 14048 480 14104
rect 0 14016 480 14048
rect 14917 13970 14983 13973
rect 18462 13970 18522 14288
rect 14917 13968 18522 13970
rect 14917 13912 14922 13968
rect 14978 13912 18522 13968
rect 14917 13910 18522 13912
rect 14917 13907 14983 13910
rect 7250 13632 7570 13633
rect 7250 13568 7258 13632
rect 7322 13568 7338 13632
rect 7402 13568 7418 13632
rect 7482 13568 7498 13632
rect 7562 13568 7570 13632
rect 7250 13567 7570 13568
rect 13557 13632 13877 13633
rect 13557 13568 13565 13632
rect 13629 13568 13645 13632
rect 13709 13568 13725 13632
rect 13789 13568 13805 13632
rect 13869 13568 13877 13632
rect 13557 13567 13877 13568
rect 0 13064 480 13184
rect 4097 13088 4417 13089
rect 62 12882 122 13064
rect 4097 13024 4105 13088
rect 4169 13024 4185 13088
rect 4249 13024 4265 13088
rect 4329 13024 4345 13088
rect 4409 13024 4417 13088
rect 4097 13023 4417 13024
rect 10403 13088 10723 13089
rect 10403 13024 10411 13088
rect 10475 13024 10491 13088
rect 10555 13024 10571 13088
rect 10635 13024 10651 13088
rect 10715 13024 10723 13088
rect 10403 13023 10723 13024
rect 16710 13088 17030 13089
rect 16710 13024 16718 13088
rect 16782 13024 16798 13088
rect 16862 13024 16878 13088
rect 16942 13024 16958 13088
rect 17022 13024 17030 13088
rect 16710 13023 17030 13024
rect 14181 12882 14247 12885
rect 62 12880 14247 12882
rect 62 12824 14186 12880
rect 14242 12824 14247 12880
rect 62 12822 14247 12824
rect 14181 12819 14247 12822
rect 5257 12746 5323 12749
rect 15285 12746 15351 12749
rect 5257 12744 15351 12746
rect 5257 12688 5262 12744
rect 5318 12688 15290 12744
rect 15346 12688 15351 12744
rect 5257 12686 15351 12688
rect 5257 12683 5323 12686
rect 15285 12683 15351 12686
rect 7250 12544 7570 12545
rect 7250 12480 7258 12544
rect 7322 12480 7338 12544
rect 7402 12480 7418 12544
rect 7482 12480 7498 12544
rect 7562 12480 7570 12544
rect 7250 12479 7570 12480
rect 13557 12544 13877 12545
rect 13557 12480 13565 12544
rect 13629 12480 13645 12544
rect 13709 12480 13725 12544
rect 13789 12480 13805 12544
rect 13869 12480 13877 12544
rect 13557 12479 13877 12480
rect 0 12064 480 12096
rect 0 12008 110 12064
rect 166 12008 480 12064
rect 0 11976 480 12008
rect 4097 12000 4417 12001
rect 4097 11936 4105 12000
rect 4169 11936 4185 12000
rect 4249 11936 4265 12000
rect 4329 11936 4345 12000
rect 4409 11936 4417 12000
rect 4097 11935 4417 11936
rect 10403 12000 10723 12001
rect 10403 11936 10411 12000
rect 10475 11936 10491 12000
rect 10555 11936 10571 12000
rect 10635 11936 10651 12000
rect 10715 11936 10723 12000
rect 10403 11935 10723 11936
rect 16710 12000 17030 12001
rect 16710 11936 16718 12000
rect 16782 11936 16798 12000
rect 16862 11936 16878 12000
rect 16942 11936 16958 12000
rect 17022 11936 17030 12000
rect 16710 11935 17030 11936
rect 18439 11797 18919 11824
rect 18413 11794 18919 11797
rect 18332 11792 18919 11794
rect 18332 11736 18418 11792
rect 18474 11736 18919 11792
rect 18332 11734 18919 11736
rect 18413 11731 18919 11734
rect 18439 11704 18919 11731
rect 7250 11456 7570 11457
rect 7250 11392 7258 11456
rect 7322 11392 7338 11456
rect 7402 11392 7418 11456
rect 7482 11392 7498 11456
rect 7562 11392 7570 11456
rect 7250 11391 7570 11392
rect 13557 11456 13877 11457
rect 13557 11392 13565 11456
rect 13629 11392 13645 11456
rect 13709 11392 13725 11456
rect 13789 11392 13805 11456
rect 13869 11392 13877 11456
rect 13557 11391 13877 11392
rect 0 10888 480 11008
rect 4097 10912 4417 10913
rect 62 10706 122 10888
rect 4097 10848 4105 10912
rect 4169 10848 4185 10912
rect 4249 10848 4265 10912
rect 4329 10848 4345 10912
rect 4409 10848 4417 10912
rect 4097 10847 4417 10848
rect 10403 10912 10723 10913
rect 10403 10848 10411 10912
rect 10475 10848 10491 10912
rect 10555 10848 10571 10912
rect 10635 10848 10651 10912
rect 10715 10848 10723 10912
rect 10403 10847 10723 10848
rect 16710 10912 17030 10913
rect 16710 10848 16718 10912
rect 16782 10848 16798 10912
rect 16862 10848 16878 10912
rect 16942 10848 16958 10912
rect 17022 10848 17030 10912
rect 16710 10847 17030 10848
rect 5165 10706 5231 10709
rect 62 10704 5231 10706
rect 62 10648 5170 10704
rect 5226 10648 5231 10704
rect 62 10646 5231 10648
rect 5165 10643 5231 10646
rect 7250 10368 7570 10369
rect 7250 10304 7258 10368
rect 7322 10304 7338 10368
rect 7402 10304 7418 10368
rect 7482 10304 7498 10368
rect 7562 10304 7570 10368
rect 7250 10303 7570 10304
rect 13557 10368 13877 10369
rect 13557 10304 13565 10368
rect 13629 10304 13645 10368
rect 13709 10304 13725 10368
rect 13789 10304 13805 10368
rect 13869 10304 13877 10368
rect 13557 10303 13877 10304
rect 0 9888 480 9920
rect 0 9832 110 9888
rect 166 9832 480 9888
rect 0 9800 480 9832
rect 4097 9824 4417 9825
rect 4097 9760 4105 9824
rect 4169 9760 4185 9824
rect 4249 9760 4265 9824
rect 4329 9760 4345 9824
rect 4409 9760 4417 9824
rect 4097 9759 4417 9760
rect 10403 9824 10723 9825
rect 10403 9760 10411 9824
rect 10475 9760 10491 9824
rect 10555 9760 10571 9824
rect 10635 9760 10651 9824
rect 10715 9760 10723 9824
rect 10403 9759 10723 9760
rect 16710 9824 17030 9825
rect 16710 9760 16718 9824
rect 16782 9760 16798 9824
rect 16862 9760 16878 9824
rect 16942 9760 16958 9824
rect 17022 9760 17030 9824
rect 16710 9759 17030 9760
rect 7250 9280 7570 9281
rect 7250 9216 7258 9280
rect 7322 9216 7338 9280
rect 7402 9216 7418 9280
rect 7482 9216 7498 9280
rect 7562 9216 7570 9280
rect 7250 9215 7570 9216
rect 13557 9280 13877 9281
rect 13557 9216 13565 9280
rect 13629 9216 13645 9280
rect 13709 9216 13725 9280
rect 13789 9216 13805 9280
rect 13869 9216 13877 9280
rect 13557 9215 13877 9216
rect 18439 9120 18919 9240
rect 0 8848 480 8968
rect 17033 8938 17099 8941
rect 18462 8938 18522 9120
rect 17033 8936 18522 8938
rect 17033 8880 17038 8936
rect 17094 8880 18522 8936
rect 17033 8878 18522 8880
rect 17033 8875 17099 8878
rect 62 8530 122 8848
rect 4097 8736 4417 8737
rect 4097 8672 4105 8736
rect 4169 8672 4185 8736
rect 4249 8672 4265 8736
rect 4329 8672 4345 8736
rect 4409 8672 4417 8736
rect 4097 8671 4417 8672
rect 10403 8736 10723 8737
rect 10403 8672 10411 8736
rect 10475 8672 10491 8736
rect 10555 8672 10571 8736
rect 10635 8672 10651 8736
rect 10715 8672 10723 8736
rect 10403 8671 10723 8672
rect 16710 8736 17030 8737
rect 16710 8672 16718 8736
rect 16782 8672 16798 8736
rect 16862 8672 16878 8736
rect 16942 8672 16958 8736
rect 17022 8672 17030 8736
rect 16710 8671 17030 8672
rect 3969 8530 4035 8533
rect 62 8528 4035 8530
rect 62 8472 3974 8528
rect 4030 8472 4035 8528
rect 62 8470 4035 8472
rect 3969 8467 4035 8470
rect 1853 8394 1919 8397
rect 62 8392 1919 8394
rect 62 8336 1858 8392
rect 1914 8336 1919 8392
rect 62 8334 1919 8336
rect 62 7880 122 8334
rect 1853 8331 1919 8334
rect 7250 8192 7570 8193
rect 7250 8128 7258 8192
rect 7322 8128 7338 8192
rect 7402 8128 7418 8192
rect 7482 8128 7498 8192
rect 7562 8128 7570 8192
rect 7250 8127 7570 8128
rect 13557 8192 13877 8193
rect 13557 8128 13565 8192
rect 13629 8128 13645 8192
rect 13709 8128 13725 8192
rect 13789 8128 13805 8192
rect 13869 8128 13877 8192
rect 13557 8127 13877 8128
rect 0 7760 480 7880
rect 4097 7648 4417 7649
rect 4097 7584 4105 7648
rect 4169 7584 4185 7648
rect 4249 7584 4265 7648
rect 4329 7584 4345 7648
rect 4409 7584 4417 7648
rect 4097 7583 4417 7584
rect 10403 7648 10723 7649
rect 10403 7584 10411 7648
rect 10475 7584 10491 7648
rect 10555 7584 10571 7648
rect 10635 7584 10651 7648
rect 10715 7584 10723 7648
rect 10403 7583 10723 7584
rect 16710 7648 17030 7649
rect 16710 7584 16718 7648
rect 16782 7584 16798 7648
rect 16862 7584 16878 7648
rect 16942 7584 16958 7648
rect 17022 7584 17030 7648
rect 16710 7583 17030 7584
rect 7250 7104 7570 7105
rect 7250 7040 7258 7104
rect 7322 7040 7338 7104
rect 7402 7040 7418 7104
rect 7482 7040 7498 7104
rect 7562 7040 7570 7104
rect 7250 7039 7570 7040
rect 13557 7104 13877 7105
rect 13557 7040 13565 7104
rect 13629 7040 13645 7104
rect 13709 7040 13725 7104
rect 13789 7040 13805 7104
rect 13869 7040 13877 7104
rect 13557 7039 13877 7040
rect 0 6672 480 6792
rect 62 6354 122 6672
rect 4097 6560 4417 6561
rect 4097 6496 4105 6560
rect 4169 6496 4185 6560
rect 4249 6496 4265 6560
rect 4329 6496 4345 6560
rect 4409 6496 4417 6560
rect 4097 6495 4417 6496
rect 10403 6560 10723 6561
rect 10403 6496 10411 6560
rect 10475 6496 10491 6560
rect 10555 6496 10571 6560
rect 10635 6496 10651 6560
rect 10715 6496 10723 6560
rect 10403 6495 10723 6496
rect 16710 6560 17030 6561
rect 16710 6496 16718 6560
rect 16782 6496 16798 6560
rect 16862 6496 16878 6560
rect 16942 6496 16958 6560
rect 17022 6496 17030 6560
rect 16710 6495 17030 6496
rect 18439 6400 18919 6520
rect 1669 6354 1735 6357
rect 62 6352 1735 6354
rect 62 6296 1674 6352
rect 1730 6296 1735 6352
rect 62 6294 1735 6296
rect 1669 6291 1735 6294
rect 12985 6218 13051 6221
rect 18462 6218 18522 6400
rect 12985 6216 18522 6218
rect 12985 6160 12990 6216
rect 13046 6160 18522 6216
rect 12985 6158 18522 6160
rect 12985 6155 13051 6158
rect 7250 6016 7570 6017
rect 7250 5952 7258 6016
rect 7322 5952 7338 6016
rect 7402 5952 7418 6016
rect 7482 5952 7498 6016
rect 7562 5952 7570 6016
rect 7250 5951 7570 5952
rect 13557 6016 13877 6017
rect 13557 5952 13565 6016
rect 13629 5952 13645 6016
rect 13709 5952 13725 6016
rect 13789 5952 13805 6016
rect 13869 5952 13877 6016
rect 13557 5951 13877 5952
rect 0 5672 480 5704
rect 0 5616 110 5672
rect 166 5616 480 5672
rect 0 5584 480 5616
rect 4097 5472 4417 5473
rect 4097 5408 4105 5472
rect 4169 5408 4185 5472
rect 4249 5408 4265 5472
rect 4329 5408 4345 5472
rect 4409 5408 4417 5472
rect 4097 5407 4417 5408
rect 10403 5472 10723 5473
rect 10403 5408 10411 5472
rect 10475 5408 10491 5472
rect 10555 5408 10571 5472
rect 10635 5408 10651 5472
rect 10715 5408 10723 5472
rect 10403 5407 10723 5408
rect 16710 5472 17030 5473
rect 16710 5408 16718 5472
rect 16782 5408 16798 5472
rect 16862 5408 16878 5472
rect 16942 5408 16958 5472
rect 17022 5408 17030 5472
rect 16710 5407 17030 5408
rect 2773 5266 2839 5269
rect 62 5264 2839 5266
rect 62 5208 2778 5264
rect 2834 5208 2839 5264
rect 62 5206 2839 5208
rect 62 4752 122 5206
rect 2773 5203 2839 5206
rect 7250 4928 7570 4929
rect 7250 4864 7258 4928
rect 7322 4864 7338 4928
rect 7402 4864 7418 4928
rect 7482 4864 7498 4928
rect 7562 4864 7570 4928
rect 7250 4863 7570 4864
rect 13557 4928 13877 4929
rect 13557 4864 13565 4928
rect 13629 4864 13645 4928
rect 13709 4864 13725 4928
rect 13789 4864 13805 4928
rect 13869 4864 13877 4928
rect 13557 4863 13877 4864
rect 0 4632 480 4752
rect 4097 4384 4417 4385
rect 4097 4320 4105 4384
rect 4169 4320 4185 4384
rect 4249 4320 4265 4384
rect 4329 4320 4345 4384
rect 4409 4320 4417 4384
rect 4097 4319 4417 4320
rect 10403 4384 10723 4385
rect 10403 4320 10411 4384
rect 10475 4320 10491 4384
rect 10555 4320 10571 4384
rect 10635 4320 10651 4384
rect 10715 4320 10723 4384
rect 10403 4319 10723 4320
rect 16710 4384 17030 4385
rect 16710 4320 16718 4384
rect 16782 4320 16798 4384
rect 16862 4320 16878 4384
rect 16942 4320 16958 4384
rect 17022 4320 17030 4384
rect 16710 4319 17030 4320
rect 16481 4178 16547 4181
rect 16481 4176 18522 4178
rect 16481 4120 16486 4176
rect 16542 4120 18522 4176
rect 16481 4118 18522 4120
rect 16481 4115 16547 4118
rect 18462 3936 18522 4118
rect 7250 3840 7570 3841
rect 7250 3776 7258 3840
rect 7322 3776 7338 3840
rect 7402 3776 7418 3840
rect 7482 3776 7498 3840
rect 7562 3776 7570 3840
rect 7250 3775 7570 3776
rect 13557 3840 13877 3841
rect 13557 3776 13565 3840
rect 13629 3776 13645 3840
rect 13709 3776 13725 3840
rect 13789 3776 13805 3840
rect 13869 3776 13877 3840
rect 18439 3816 18919 3936
rect 13557 3775 13877 3776
rect 0 3632 480 3664
rect 0 3576 110 3632
rect 166 3576 480 3632
rect 0 3544 480 3576
rect 4097 3296 4417 3297
rect 4097 3232 4105 3296
rect 4169 3232 4185 3296
rect 4249 3232 4265 3296
rect 4329 3232 4345 3296
rect 4409 3232 4417 3296
rect 4097 3231 4417 3232
rect 10403 3296 10723 3297
rect 10403 3232 10411 3296
rect 10475 3232 10491 3296
rect 10555 3232 10571 3296
rect 10635 3232 10651 3296
rect 10715 3232 10723 3296
rect 10403 3231 10723 3232
rect 16710 3296 17030 3297
rect 16710 3232 16718 3296
rect 16782 3232 16798 3296
rect 16862 3232 16878 3296
rect 16942 3232 16958 3296
rect 17022 3232 17030 3296
rect 16710 3231 17030 3232
rect 6361 3090 6427 3093
rect 62 3088 6427 3090
rect 62 3032 6366 3088
rect 6422 3032 6427 3088
rect 62 3030 6427 3032
rect 62 2576 122 3030
rect 6361 3027 6427 3030
rect 7250 2752 7570 2753
rect 7250 2688 7258 2752
rect 7322 2688 7338 2752
rect 7402 2688 7418 2752
rect 7482 2688 7498 2752
rect 7562 2688 7570 2752
rect 7250 2687 7570 2688
rect 13557 2752 13877 2753
rect 13557 2688 13565 2752
rect 13629 2688 13645 2752
rect 13709 2688 13725 2752
rect 13789 2688 13805 2752
rect 13869 2688 13877 2752
rect 13557 2687 13877 2688
rect 0 2456 480 2576
rect 4097 2208 4417 2209
rect 4097 2144 4105 2208
rect 4169 2144 4185 2208
rect 4249 2144 4265 2208
rect 4329 2144 4345 2208
rect 4409 2144 4417 2208
rect 4097 2143 4417 2144
rect 10403 2208 10723 2209
rect 10403 2144 10411 2208
rect 10475 2144 10491 2208
rect 10555 2144 10571 2208
rect 10635 2144 10651 2208
rect 10715 2144 10723 2208
rect 10403 2143 10723 2144
rect 16710 2208 17030 2209
rect 16710 2144 16718 2208
rect 16782 2144 16798 2208
rect 16862 2144 16878 2208
rect 16942 2144 16958 2208
rect 17022 2144 17030 2208
rect 16710 2143 17030 2144
rect 14273 1866 14339 1869
rect 14273 1864 18522 1866
rect 14273 1808 14278 1864
rect 14334 1808 18522 1864
rect 14273 1806 18522 1808
rect 14273 1803 14339 1806
rect 0 1368 480 1488
rect 18462 1352 18522 1806
rect 18439 1232 18919 1352
rect 0 416 480 536
<< via3 >>
rect 4105 18524 4169 18528
rect 4105 18468 4109 18524
rect 4109 18468 4165 18524
rect 4165 18468 4169 18524
rect 4105 18464 4169 18468
rect 4185 18524 4249 18528
rect 4185 18468 4189 18524
rect 4189 18468 4245 18524
rect 4245 18468 4249 18524
rect 4185 18464 4249 18468
rect 4265 18524 4329 18528
rect 4265 18468 4269 18524
rect 4269 18468 4325 18524
rect 4325 18468 4329 18524
rect 4265 18464 4329 18468
rect 4345 18524 4409 18528
rect 4345 18468 4349 18524
rect 4349 18468 4405 18524
rect 4405 18468 4409 18524
rect 4345 18464 4409 18468
rect 10411 18524 10475 18528
rect 10411 18468 10415 18524
rect 10415 18468 10471 18524
rect 10471 18468 10475 18524
rect 10411 18464 10475 18468
rect 10491 18524 10555 18528
rect 10491 18468 10495 18524
rect 10495 18468 10551 18524
rect 10551 18468 10555 18524
rect 10491 18464 10555 18468
rect 10571 18524 10635 18528
rect 10571 18468 10575 18524
rect 10575 18468 10631 18524
rect 10631 18468 10635 18524
rect 10571 18464 10635 18468
rect 10651 18524 10715 18528
rect 10651 18468 10655 18524
rect 10655 18468 10711 18524
rect 10711 18468 10715 18524
rect 10651 18464 10715 18468
rect 16718 18524 16782 18528
rect 16718 18468 16722 18524
rect 16722 18468 16778 18524
rect 16778 18468 16782 18524
rect 16718 18464 16782 18468
rect 16798 18524 16862 18528
rect 16798 18468 16802 18524
rect 16802 18468 16858 18524
rect 16858 18468 16862 18524
rect 16798 18464 16862 18468
rect 16878 18524 16942 18528
rect 16878 18468 16882 18524
rect 16882 18468 16938 18524
rect 16938 18468 16942 18524
rect 16878 18464 16942 18468
rect 16958 18524 17022 18528
rect 16958 18468 16962 18524
rect 16962 18468 17018 18524
rect 17018 18468 17022 18524
rect 16958 18464 17022 18468
rect 7258 17980 7322 17984
rect 7258 17924 7262 17980
rect 7262 17924 7318 17980
rect 7318 17924 7322 17980
rect 7258 17920 7322 17924
rect 7338 17980 7402 17984
rect 7338 17924 7342 17980
rect 7342 17924 7398 17980
rect 7398 17924 7402 17980
rect 7338 17920 7402 17924
rect 7418 17980 7482 17984
rect 7418 17924 7422 17980
rect 7422 17924 7478 17980
rect 7478 17924 7482 17980
rect 7418 17920 7482 17924
rect 7498 17980 7562 17984
rect 7498 17924 7502 17980
rect 7502 17924 7558 17980
rect 7558 17924 7562 17980
rect 7498 17920 7562 17924
rect 13565 17980 13629 17984
rect 13565 17924 13569 17980
rect 13569 17924 13625 17980
rect 13625 17924 13629 17980
rect 13565 17920 13629 17924
rect 13645 17980 13709 17984
rect 13645 17924 13649 17980
rect 13649 17924 13705 17980
rect 13705 17924 13709 17980
rect 13645 17920 13709 17924
rect 13725 17980 13789 17984
rect 13725 17924 13729 17980
rect 13729 17924 13785 17980
rect 13785 17924 13789 17980
rect 13725 17920 13789 17924
rect 13805 17980 13869 17984
rect 13805 17924 13809 17980
rect 13809 17924 13865 17980
rect 13865 17924 13869 17980
rect 13805 17920 13869 17924
rect 4105 17436 4169 17440
rect 4105 17380 4109 17436
rect 4109 17380 4165 17436
rect 4165 17380 4169 17436
rect 4105 17376 4169 17380
rect 4185 17436 4249 17440
rect 4185 17380 4189 17436
rect 4189 17380 4245 17436
rect 4245 17380 4249 17436
rect 4185 17376 4249 17380
rect 4265 17436 4329 17440
rect 4265 17380 4269 17436
rect 4269 17380 4325 17436
rect 4325 17380 4329 17436
rect 4265 17376 4329 17380
rect 4345 17436 4409 17440
rect 4345 17380 4349 17436
rect 4349 17380 4405 17436
rect 4405 17380 4409 17436
rect 4345 17376 4409 17380
rect 10411 17436 10475 17440
rect 10411 17380 10415 17436
rect 10415 17380 10471 17436
rect 10471 17380 10475 17436
rect 10411 17376 10475 17380
rect 10491 17436 10555 17440
rect 10491 17380 10495 17436
rect 10495 17380 10551 17436
rect 10551 17380 10555 17436
rect 10491 17376 10555 17380
rect 10571 17436 10635 17440
rect 10571 17380 10575 17436
rect 10575 17380 10631 17436
rect 10631 17380 10635 17436
rect 10571 17376 10635 17380
rect 10651 17436 10715 17440
rect 10651 17380 10655 17436
rect 10655 17380 10711 17436
rect 10711 17380 10715 17436
rect 10651 17376 10715 17380
rect 16718 17436 16782 17440
rect 16718 17380 16722 17436
rect 16722 17380 16778 17436
rect 16778 17380 16782 17436
rect 16718 17376 16782 17380
rect 16798 17436 16862 17440
rect 16798 17380 16802 17436
rect 16802 17380 16858 17436
rect 16858 17380 16862 17436
rect 16798 17376 16862 17380
rect 16878 17436 16942 17440
rect 16878 17380 16882 17436
rect 16882 17380 16938 17436
rect 16938 17380 16942 17436
rect 16878 17376 16942 17380
rect 16958 17436 17022 17440
rect 16958 17380 16962 17436
rect 16962 17380 17018 17436
rect 17018 17380 17022 17436
rect 16958 17376 17022 17380
rect 7258 16892 7322 16896
rect 7258 16836 7262 16892
rect 7262 16836 7318 16892
rect 7318 16836 7322 16892
rect 7258 16832 7322 16836
rect 7338 16892 7402 16896
rect 7338 16836 7342 16892
rect 7342 16836 7398 16892
rect 7398 16836 7402 16892
rect 7338 16832 7402 16836
rect 7418 16892 7482 16896
rect 7418 16836 7422 16892
rect 7422 16836 7478 16892
rect 7478 16836 7482 16892
rect 7418 16832 7482 16836
rect 7498 16892 7562 16896
rect 7498 16836 7502 16892
rect 7502 16836 7558 16892
rect 7558 16836 7562 16892
rect 7498 16832 7562 16836
rect 13565 16892 13629 16896
rect 13565 16836 13569 16892
rect 13569 16836 13625 16892
rect 13625 16836 13629 16892
rect 13565 16832 13629 16836
rect 13645 16892 13709 16896
rect 13645 16836 13649 16892
rect 13649 16836 13705 16892
rect 13705 16836 13709 16892
rect 13645 16832 13709 16836
rect 13725 16892 13789 16896
rect 13725 16836 13729 16892
rect 13729 16836 13785 16892
rect 13785 16836 13789 16892
rect 13725 16832 13789 16836
rect 13805 16892 13869 16896
rect 13805 16836 13809 16892
rect 13809 16836 13865 16892
rect 13865 16836 13869 16892
rect 13805 16832 13869 16836
rect 4105 16348 4169 16352
rect 4105 16292 4109 16348
rect 4109 16292 4165 16348
rect 4165 16292 4169 16348
rect 4105 16288 4169 16292
rect 4185 16348 4249 16352
rect 4185 16292 4189 16348
rect 4189 16292 4245 16348
rect 4245 16292 4249 16348
rect 4185 16288 4249 16292
rect 4265 16348 4329 16352
rect 4265 16292 4269 16348
rect 4269 16292 4325 16348
rect 4325 16292 4329 16348
rect 4265 16288 4329 16292
rect 4345 16348 4409 16352
rect 4345 16292 4349 16348
rect 4349 16292 4405 16348
rect 4405 16292 4409 16348
rect 4345 16288 4409 16292
rect 10411 16348 10475 16352
rect 10411 16292 10415 16348
rect 10415 16292 10471 16348
rect 10471 16292 10475 16348
rect 10411 16288 10475 16292
rect 10491 16348 10555 16352
rect 10491 16292 10495 16348
rect 10495 16292 10551 16348
rect 10551 16292 10555 16348
rect 10491 16288 10555 16292
rect 10571 16348 10635 16352
rect 10571 16292 10575 16348
rect 10575 16292 10631 16348
rect 10631 16292 10635 16348
rect 10571 16288 10635 16292
rect 10651 16348 10715 16352
rect 10651 16292 10655 16348
rect 10655 16292 10711 16348
rect 10711 16292 10715 16348
rect 10651 16288 10715 16292
rect 16718 16348 16782 16352
rect 16718 16292 16722 16348
rect 16722 16292 16778 16348
rect 16778 16292 16782 16348
rect 16718 16288 16782 16292
rect 16798 16348 16862 16352
rect 16798 16292 16802 16348
rect 16802 16292 16858 16348
rect 16858 16292 16862 16348
rect 16798 16288 16862 16292
rect 16878 16348 16942 16352
rect 16878 16292 16882 16348
rect 16882 16292 16938 16348
rect 16938 16292 16942 16348
rect 16878 16288 16942 16292
rect 16958 16348 17022 16352
rect 16958 16292 16962 16348
rect 16962 16292 17018 16348
rect 17018 16292 17022 16348
rect 16958 16288 17022 16292
rect 7258 15804 7322 15808
rect 7258 15748 7262 15804
rect 7262 15748 7318 15804
rect 7318 15748 7322 15804
rect 7258 15744 7322 15748
rect 7338 15804 7402 15808
rect 7338 15748 7342 15804
rect 7342 15748 7398 15804
rect 7398 15748 7402 15804
rect 7338 15744 7402 15748
rect 7418 15804 7482 15808
rect 7418 15748 7422 15804
rect 7422 15748 7478 15804
rect 7478 15748 7482 15804
rect 7418 15744 7482 15748
rect 7498 15804 7562 15808
rect 7498 15748 7502 15804
rect 7502 15748 7558 15804
rect 7558 15748 7562 15804
rect 7498 15744 7562 15748
rect 13565 15804 13629 15808
rect 13565 15748 13569 15804
rect 13569 15748 13625 15804
rect 13625 15748 13629 15804
rect 13565 15744 13629 15748
rect 13645 15804 13709 15808
rect 13645 15748 13649 15804
rect 13649 15748 13705 15804
rect 13705 15748 13709 15804
rect 13645 15744 13709 15748
rect 13725 15804 13789 15808
rect 13725 15748 13729 15804
rect 13729 15748 13785 15804
rect 13785 15748 13789 15804
rect 13725 15744 13789 15748
rect 13805 15804 13869 15808
rect 13805 15748 13809 15804
rect 13809 15748 13865 15804
rect 13865 15748 13869 15804
rect 13805 15744 13869 15748
rect 4105 15260 4169 15264
rect 4105 15204 4109 15260
rect 4109 15204 4165 15260
rect 4165 15204 4169 15260
rect 4105 15200 4169 15204
rect 4185 15260 4249 15264
rect 4185 15204 4189 15260
rect 4189 15204 4245 15260
rect 4245 15204 4249 15260
rect 4185 15200 4249 15204
rect 4265 15260 4329 15264
rect 4265 15204 4269 15260
rect 4269 15204 4325 15260
rect 4325 15204 4329 15260
rect 4265 15200 4329 15204
rect 4345 15260 4409 15264
rect 4345 15204 4349 15260
rect 4349 15204 4405 15260
rect 4405 15204 4409 15260
rect 4345 15200 4409 15204
rect 10411 15260 10475 15264
rect 10411 15204 10415 15260
rect 10415 15204 10471 15260
rect 10471 15204 10475 15260
rect 10411 15200 10475 15204
rect 10491 15260 10555 15264
rect 10491 15204 10495 15260
rect 10495 15204 10551 15260
rect 10551 15204 10555 15260
rect 10491 15200 10555 15204
rect 10571 15260 10635 15264
rect 10571 15204 10575 15260
rect 10575 15204 10631 15260
rect 10631 15204 10635 15260
rect 10571 15200 10635 15204
rect 10651 15260 10715 15264
rect 10651 15204 10655 15260
rect 10655 15204 10711 15260
rect 10711 15204 10715 15260
rect 10651 15200 10715 15204
rect 16718 15260 16782 15264
rect 16718 15204 16722 15260
rect 16722 15204 16778 15260
rect 16778 15204 16782 15260
rect 16718 15200 16782 15204
rect 16798 15260 16862 15264
rect 16798 15204 16802 15260
rect 16802 15204 16858 15260
rect 16858 15204 16862 15260
rect 16798 15200 16862 15204
rect 16878 15260 16942 15264
rect 16878 15204 16882 15260
rect 16882 15204 16938 15260
rect 16938 15204 16942 15260
rect 16878 15200 16942 15204
rect 16958 15260 17022 15264
rect 16958 15204 16962 15260
rect 16962 15204 17018 15260
rect 17018 15204 17022 15260
rect 16958 15200 17022 15204
rect 7258 14716 7322 14720
rect 7258 14660 7262 14716
rect 7262 14660 7318 14716
rect 7318 14660 7322 14716
rect 7258 14656 7322 14660
rect 7338 14716 7402 14720
rect 7338 14660 7342 14716
rect 7342 14660 7398 14716
rect 7398 14660 7402 14716
rect 7338 14656 7402 14660
rect 7418 14716 7482 14720
rect 7418 14660 7422 14716
rect 7422 14660 7478 14716
rect 7478 14660 7482 14716
rect 7418 14656 7482 14660
rect 7498 14716 7562 14720
rect 7498 14660 7502 14716
rect 7502 14660 7558 14716
rect 7558 14660 7562 14716
rect 7498 14656 7562 14660
rect 13565 14716 13629 14720
rect 13565 14660 13569 14716
rect 13569 14660 13625 14716
rect 13625 14660 13629 14716
rect 13565 14656 13629 14660
rect 13645 14716 13709 14720
rect 13645 14660 13649 14716
rect 13649 14660 13705 14716
rect 13705 14660 13709 14716
rect 13645 14656 13709 14660
rect 13725 14716 13789 14720
rect 13725 14660 13729 14716
rect 13729 14660 13785 14716
rect 13785 14660 13789 14716
rect 13725 14656 13789 14660
rect 13805 14716 13869 14720
rect 13805 14660 13809 14716
rect 13809 14660 13865 14716
rect 13865 14660 13869 14716
rect 13805 14656 13869 14660
rect 4105 14172 4169 14176
rect 4105 14116 4109 14172
rect 4109 14116 4165 14172
rect 4165 14116 4169 14172
rect 4105 14112 4169 14116
rect 4185 14172 4249 14176
rect 4185 14116 4189 14172
rect 4189 14116 4245 14172
rect 4245 14116 4249 14172
rect 4185 14112 4249 14116
rect 4265 14172 4329 14176
rect 4265 14116 4269 14172
rect 4269 14116 4325 14172
rect 4325 14116 4329 14172
rect 4265 14112 4329 14116
rect 4345 14172 4409 14176
rect 4345 14116 4349 14172
rect 4349 14116 4405 14172
rect 4405 14116 4409 14172
rect 4345 14112 4409 14116
rect 10411 14172 10475 14176
rect 10411 14116 10415 14172
rect 10415 14116 10471 14172
rect 10471 14116 10475 14172
rect 10411 14112 10475 14116
rect 10491 14172 10555 14176
rect 10491 14116 10495 14172
rect 10495 14116 10551 14172
rect 10551 14116 10555 14172
rect 10491 14112 10555 14116
rect 10571 14172 10635 14176
rect 10571 14116 10575 14172
rect 10575 14116 10631 14172
rect 10631 14116 10635 14172
rect 10571 14112 10635 14116
rect 10651 14172 10715 14176
rect 10651 14116 10655 14172
rect 10655 14116 10711 14172
rect 10711 14116 10715 14172
rect 10651 14112 10715 14116
rect 16718 14172 16782 14176
rect 16718 14116 16722 14172
rect 16722 14116 16778 14172
rect 16778 14116 16782 14172
rect 16718 14112 16782 14116
rect 16798 14172 16862 14176
rect 16798 14116 16802 14172
rect 16802 14116 16858 14172
rect 16858 14116 16862 14172
rect 16798 14112 16862 14116
rect 16878 14172 16942 14176
rect 16878 14116 16882 14172
rect 16882 14116 16938 14172
rect 16938 14116 16942 14172
rect 16878 14112 16942 14116
rect 16958 14172 17022 14176
rect 16958 14116 16962 14172
rect 16962 14116 17018 14172
rect 17018 14116 17022 14172
rect 16958 14112 17022 14116
rect 7258 13628 7322 13632
rect 7258 13572 7262 13628
rect 7262 13572 7318 13628
rect 7318 13572 7322 13628
rect 7258 13568 7322 13572
rect 7338 13628 7402 13632
rect 7338 13572 7342 13628
rect 7342 13572 7398 13628
rect 7398 13572 7402 13628
rect 7338 13568 7402 13572
rect 7418 13628 7482 13632
rect 7418 13572 7422 13628
rect 7422 13572 7478 13628
rect 7478 13572 7482 13628
rect 7418 13568 7482 13572
rect 7498 13628 7562 13632
rect 7498 13572 7502 13628
rect 7502 13572 7558 13628
rect 7558 13572 7562 13628
rect 7498 13568 7562 13572
rect 13565 13628 13629 13632
rect 13565 13572 13569 13628
rect 13569 13572 13625 13628
rect 13625 13572 13629 13628
rect 13565 13568 13629 13572
rect 13645 13628 13709 13632
rect 13645 13572 13649 13628
rect 13649 13572 13705 13628
rect 13705 13572 13709 13628
rect 13645 13568 13709 13572
rect 13725 13628 13789 13632
rect 13725 13572 13729 13628
rect 13729 13572 13785 13628
rect 13785 13572 13789 13628
rect 13725 13568 13789 13572
rect 13805 13628 13869 13632
rect 13805 13572 13809 13628
rect 13809 13572 13865 13628
rect 13865 13572 13869 13628
rect 13805 13568 13869 13572
rect 4105 13084 4169 13088
rect 4105 13028 4109 13084
rect 4109 13028 4165 13084
rect 4165 13028 4169 13084
rect 4105 13024 4169 13028
rect 4185 13084 4249 13088
rect 4185 13028 4189 13084
rect 4189 13028 4245 13084
rect 4245 13028 4249 13084
rect 4185 13024 4249 13028
rect 4265 13084 4329 13088
rect 4265 13028 4269 13084
rect 4269 13028 4325 13084
rect 4325 13028 4329 13084
rect 4265 13024 4329 13028
rect 4345 13084 4409 13088
rect 4345 13028 4349 13084
rect 4349 13028 4405 13084
rect 4405 13028 4409 13084
rect 4345 13024 4409 13028
rect 10411 13084 10475 13088
rect 10411 13028 10415 13084
rect 10415 13028 10471 13084
rect 10471 13028 10475 13084
rect 10411 13024 10475 13028
rect 10491 13084 10555 13088
rect 10491 13028 10495 13084
rect 10495 13028 10551 13084
rect 10551 13028 10555 13084
rect 10491 13024 10555 13028
rect 10571 13084 10635 13088
rect 10571 13028 10575 13084
rect 10575 13028 10631 13084
rect 10631 13028 10635 13084
rect 10571 13024 10635 13028
rect 10651 13084 10715 13088
rect 10651 13028 10655 13084
rect 10655 13028 10711 13084
rect 10711 13028 10715 13084
rect 10651 13024 10715 13028
rect 16718 13084 16782 13088
rect 16718 13028 16722 13084
rect 16722 13028 16778 13084
rect 16778 13028 16782 13084
rect 16718 13024 16782 13028
rect 16798 13084 16862 13088
rect 16798 13028 16802 13084
rect 16802 13028 16858 13084
rect 16858 13028 16862 13084
rect 16798 13024 16862 13028
rect 16878 13084 16942 13088
rect 16878 13028 16882 13084
rect 16882 13028 16938 13084
rect 16938 13028 16942 13084
rect 16878 13024 16942 13028
rect 16958 13084 17022 13088
rect 16958 13028 16962 13084
rect 16962 13028 17018 13084
rect 17018 13028 17022 13084
rect 16958 13024 17022 13028
rect 7258 12540 7322 12544
rect 7258 12484 7262 12540
rect 7262 12484 7318 12540
rect 7318 12484 7322 12540
rect 7258 12480 7322 12484
rect 7338 12540 7402 12544
rect 7338 12484 7342 12540
rect 7342 12484 7398 12540
rect 7398 12484 7402 12540
rect 7338 12480 7402 12484
rect 7418 12540 7482 12544
rect 7418 12484 7422 12540
rect 7422 12484 7478 12540
rect 7478 12484 7482 12540
rect 7418 12480 7482 12484
rect 7498 12540 7562 12544
rect 7498 12484 7502 12540
rect 7502 12484 7558 12540
rect 7558 12484 7562 12540
rect 7498 12480 7562 12484
rect 13565 12540 13629 12544
rect 13565 12484 13569 12540
rect 13569 12484 13625 12540
rect 13625 12484 13629 12540
rect 13565 12480 13629 12484
rect 13645 12540 13709 12544
rect 13645 12484 13649 12540
rect 13649 12484 13705 12540
rect 13705 12484 13709 12540
rect 13645 12480 13709 12484
rect 13725 12540 13789 12544
rect 13725 12484 13729 12540
rect 13729 12484 13785 12540
rect 13785 12484 13789 12540
rect 13725 12480 13789 12484
rect 13805 12540 13869 12544
rect 13805 12484 13809 12540
rect 13809 12484 13865 12540
rect 13865 12484 13869 12540
rect 13805 12480 13869 12484
rect 4105 11996 4169 12000
rect 4105 11940 4109 11996
rect 4109 11940 4165 11996
rect 4165 11940 4169 11996
rect 4105 11936 4169 11940
rect 4185 11996 4249 12000
rect 4185 11940 4189 11996
rect 4189 11940 4245 11996
rect 4245 11940 4249 11996
rect 4185 11936 4249 11940
rect 4265 11996 4329 12000
rect 4265 11940 4269 11996
rect 4269 11940 4325 11996
rect 4325 11940 4329 11996
rect 4265 11936 4329 11940
rect 4345 11996 4409 12000
rect 4345 11940 4349 11996
rect 4349 11940 4405 11996
rect 4405 11940 4409 11996
rect 4345 11936 4409 11940
rect 10411 11996 10475 12000
rect 10411 11940 10415 11996
rect 10415 11940 10471 11996
rect 10471 11940 10475 11996
rect 10411 11936 10475 11940
rect 10491 11996 10555 12000
rect 10491 11940 10495 11996
rect 10495 11940 10551 11996
rect 10551 11940 10555 11996
rect 10491 11936 10555 11940
rect 10571 11996 10635 12000
rect 10571 11940 10575 11996
rect 10575 11940 10631 11996
rect 10631 11940 10635 11996
rect 10571 11936 10635 11940
rect 10651 11996 10715 12000
rect 10651 11940 10655 11996
rect 10655 11940 10711 11996
rect 10711 11940 10715 11996
rect 10651 11936 10715 11940
rect 16718 11996 16782 12000
rect 16718 11940 16722 11996
rect 16722 11940 16778 11996
rect 16778 11940 16782 11996
rect 16718 11936 16782 11940
rect 16798 11996 16862 12000
rect 16798 11940 16802 11996
rect 16802 11940 16858 11996
rect 16858 11940 16862 11996
rect 16798 11936 16862 11940
rect 16878 11996 16942 12000
rect 16878 11940 16882 11996
rect 16882 11940 16938 11996
rect 16938 11940 16942 11996
rect 16878 11936 16942 11940
rect 16958 11996 17022 12000
rect 16958 11940 16962 11996
rect 16962 11940 17018 11996
rect 17018 11940 17022 11996
rect 16958 11936 17022 11940
rect 7258 11452 7322 11456
rect 7258 11396 7262 11452
rect 7262 11396 7318 11452
rect 7318 11396 7322 11452
rect 7258 11392 7322 11396
rect 7338 11452 7402 11456
rect 7338 11396 7342 11452
rect 7342 11396 7398 11452
rect 7398 11396 7402 11452
rect 7338 11392 7402 11396
rect 7418 11452 7482 11456
rect 7418 11396 7422 11452
rect 7422 11396 7478 11452
rect 7478 11396 7482 11452
rect 7418 11392 7482 11396
rect 7498 11452 7562 11456
rect 7498 11396 7502 11452
rect 7502 11396 7558 11452
rect 7558 11396 7562 11452
rect 7498 11392 7562 11396
rect 13565 11452 13629 11456
rect 13565 11396 13569 11452
rect 13569 11396 13625 11452
rect 13625 11396 13629 11452
rect 13565 11392 13629 11396
rect 13645 11452 13709 11456
rect 13645 11396 13649 11452
rect 13649 11396 13705 11452
rect 13705 11396 13709 11452
rect 13645 11392 13709 11396
rect 13725 11452 13789 11456
rect 13725 11396 13729 11452
rect 13729 11396 13785 11452
rect 13785 11396 13789 11452
rect 13725 11392 13789 11396
rect 13805 11452 13869 11456
rect 13805 11396 13809 11452
rect 13809 11396 13865 11452
rect 13865 11396 13869 11452
rect 13805 11392 13869 11396
rect 4105 10908 4169 10912
rect 4105 10852 4109 10908
rect 4109 10852 4165 10908
rect 4165 10852 4169 10908
rect 4105 10848 4169 10852
rect 4185 10908 4249 10912
rect 4185 10852 4189 10908
rect 4189 10852 4245 10908
rect 4245 10852 4249 10908
rect 4185 10848 4249 10852
rect 4265 10908 4329 10912
rect 4265 10852 4269 10908
rect 4269 10852 4325 10908
rect 4325 10852 4329 10908
rect 4265 10848 4329 10852
rect 4345 10908 4409 10912
rect 4345 10852 4349 10908
rect 4349 10852 4405 10908
rect 4405 10852 4409 10908
rect 4345 10848 4409 10852
rect 10411 10908 10475 10912
rect 10411 10852 10415 10908
rect 10415 10852 10471 10908
rect 10471 10852 10475 10908
rect 10411 10848 10475 10852
rect 10491 10908 10555 10912
rect 10491 10852 10495 10908
rect 10495 10852 10551 10908
rect 10551 10852 10555 10908
rect 10491 10848 10555 10852
rect 10571 10908 10635 10912
rect 10571 10852 10575 10908
rect 10575 10852 10631 10908
rect 10631 10852 10635 10908
rect 10571 10848 10635 10852
rect 10651 10908 10715 10912
rect 10651 10852 10655 10908
rect 10655 10852 10711 10908
rect 10711 10852 10715 10908
rect 10651 10848 10715 10852
rect 16718 10908 16782 10912
rect 16718 10852 16722 10908
rect 16722 10852 16778 10908
rect 16778 10852 16782 10908
rect 16718 10848 16782 10852
rect 16798 10908 16862 10912
rect 16798 10852 16802 10908
rect 16802 10852 16858 10908
rect 16858 10852 16862 10908
rect 16798 10848 16862 10852
rect 16878 10908 16942 10912
rect 16878 10852 16882 10908
rect 16882 10852 16938 10908
rect 16938 10852 16942 10908
rect 16878 10848 16942 10852
rect 16958 10908 17022 10912
rect 16958 10852 16962 10908
rect 16962 10852 17018 10908
rect 17018 10852 17022 10908
rect 16958 10848 17022 10852
rect 7258 10364 7322 10368
rect 7258 10308 7262 10364
rect 7262 10308 7318 10364
rect 7318 10308 7322 10364
rect 7258 10304 7322 10308
rect 7338 10364 7402 10368
rect 7338 10308 7342 10364
rect 7342 10308 7398 10364
rect 7398 10308 7402 10364
rect 7338 10304 7402 10308
rect 7418 10364 7482 10368
rect 7418 10308 7422 10364
rect 7422 10308 7478 10364
rect 7478 10308 7482 10364
rect 7418 10304 7482 10308
rect 7498 10364 7562 10368
rect 7498 10308 7502 10364
rect 7502 10308 7558 10364
rect 7558 10308 7562 10364
rect 7498 10304 7562 10308
rect 13565 10364 13629 10368
rect 13565 10308 13569 10364
rect 13569 10308 13625 10364
rect 13625 10308 13629 10364
rect 13565 10304 13629 10308
rect 13645 10364 13709 10368
rect 13645 10308 13649 10364
rect 13649 10308 13705 10364
rect 13705 10308 13709 10364
rect 13645 10304 13709 10308
rect 13725 10364 13789 10368
rect 13725 10308 13729 10364
rect 13729 10308 13785 10364
rect 13785 10308 13789 10364
rect 13725 10304 13789 10308
rect 13805 10364 13869 10368
rect 13805 10308 13809 10364
rect 13809 10308 13865 10364
rect 13865 10308 13869 10364
rect 13805 10304 13869 10308
rect 4105 9820 4169 9824
rect 4105 9764 4109 9820
rect 4109 9764 4165 9820
rect 4165 9764 4169 9820
rect 4105 9760 4169 9764
rect 4185 9820 4249 9824
rect 4185 9764 4189 9820
rect 4189 9764 4245 9820
rect 4245 9764 4249 9820
rect 4185 9760 4249 9764
rect 4265 9820 4329 9824
rect 4265 9764 4269 9820
rect 4269 9764 4325 9820
rect 4325 9764 4329 9820
rect 4265 9760 4329 9764
rect 4345 9820 4409 9824
rect 4345 9764 4349 9820
rect 4349 9764 4405 9820
rect 4405 9764 4409 9820
rect 4345 9760 4409 9764
rect 10411 9820 10475 9824
rect 10411 9764 10415 9820
rect 10415 9764 10471 9820
rect 10471 9764 10475 9820
rect 10411 9760 10475 9764
rect 10491 9820 10555 9824
rect 10491 9764 10495 9820
rect 10495 9764 10551 9820
rect 10551 9764 10555 9820
rect 10491 9760 10555 9764
rect 10571 9820 10635 9824
rect 10571 9764 10575 9820
rect 10575 9764 10631 9820
rect 10631 9764 10635 9820
rect 10571 9760 10635 9764
rect 10651 9820 10715 9824
rect 10651 9764 10655 9820
rect 10655 9764 10711 9820
rect 10711 9764 10715 9820
rect 10651 9760 10715 9764
rect 16718 9820 16782 9824
rect 16718 9764 16722 9820
rect 16722 9764 16778 9820
rect 16778 9764 16782 9820
rect 16718 9760 16782 9764
rect 16798 9820 16862 9824
rect 16798 9764 16802 9820
rect 16802 9764 16858 9820
rect 16858 9764 16862 9820
rect 16798 9760 16862 9764
rect 16878 9820 16942 9824
rect 16878 9764 16882 9820
rect 16882 9764 16938 9820
rect 16938 9764 16942 9820
rect 16878 9760 16942 9764
rect 16958 9820 17022 9824
rect 16958 9764 16962 9820
rect 16962 9764 17018 9820
rect 17018 9764 17022 9820
rect 16958 9760 17022 9764
rect 7258 9276 7322 9280
rect 7258 9220 7262 9276
rect 7262 9220 7318 9276
rect 7318 9220 7322 9276
rect 7258 9216 7322 9220
rect 7338 9276 7402 9280
rect 7338 9220 7342 9276
rect 7342 9220 7398 9276
rect 7398 9220 7402 9276
rect 7338 9216 7402 9220
rect 7418 9276 7482 9280
rect 7418 9220 7422 9276
rect 7422 9220 7478 9276
rect 7478 9220 7482 9276
rect 7418 9216 7482 9220
rect 7498 9276 7562 9280
rect 7498 9220 7502 9276
rect 7502 9220 7558 9276
rect 7558 9220 7562 9276
rect 7498 9216 7562 9220
rect 13565 9276 13629 9280
rect 13565 9220 13569 9276
rect 13569 9220 13625 9276
rect 13625 9220 13629 9276
rect 13565 9216 13629 9220
rect 13645 9276 13709 9280
rect 13645 9220 13649 9276
rect 13649 9220 13705 9276
rect 13705 9220 13709 9276
rect 13645 9216 13709 9220
rect 13725 9276 13789 9280
rect 13725 9220 13729 9276
rect 13729 9220 13785 9276
rect 13785 9220 13789 9276
rect 13725 9216 13789 9220
rect 13805 9276 13869 9280
rect 13805 9220 13809 9276
rect 13809 9220 13865 9276
rect 13865 9220 13869 9276
rect 13805 9216 13869 9220
rect 4105 8732 4169 8736
rect 4105 8676 4109 8732
rect 4109 8676 4165 8732
rect 4165 8676 4169 8732
rect 4105 8672 4169 8676
rect 4185 8732 4249 8736
rect 4185 8676 4189 8732
rect 4189 8676 4245 8732
rect 4245 8676 4249 8732
rect 4185 8672 4249 8676
rect 4265 8732 4329 8736
rect 4265 8676 4269 8732
rect 4269 8676 4325 8732
rect 4325 8676 4329 8732
rect 4265 8672 4329 8676
rect 4345 8732 4409 8736
rect 4345 8676 4349 8732
rect 4349 8676 4405 8732
rect 4405 8676 4409 8732
rect 4345 8672 4409 8676
rect 10411 8732 10475 8736
rect 10411 8676 10415 8732
rect 10415 8676 10471 8732
rect 10471 8676 10475 8732
rect 10411 8672 10475 8676
rect 10491 8732 10555 8736
rect 10491 8676 10495 8732
rect 10495 8676 10551 8732
rect 10551 8676 10555 8732
rect 10491 8672 10555 8676
rect 10571 8732 10635 8736
rect 10571 8676 10575 8732
rect 10575 8676 10631 8732
rect 10631 8676 10635 8732
rect 10571 8672 10635 8676
rect 10651 8732 10715 8736
rect 10651 8676 10655 8732
rect 10655 8676 10711 8732
rect 10711 8676 10715 8732
rect 10651 8672 10715 8676
rect 16718 8732 16782 8736
rect 16718 8676 16722 8732
rect 16722 8676 16778 8732
rect 16778 8676 16782 8732
rect 16718 8672 16782 8676
rect 16798 8732 16862 8736
rect 16798 8676 16802 8732
rect 16802 8676 16858 8732
rect 16858 8676 16862 8732
rect 16798 8672 16862 8676
rect 16878 8732 16942 8736
rect 16878 8676 16882 8732
rect 16882 8676 16938 8732
rect 16938 8676 16942 8732
rect 16878 8672 16942 8676
rect 16958 8732 17022 8736
rect 16958 8676 16962 8732
rect 16962 8676 17018 8732
rect 17018 8676 17022 8732
rect 16958 8672 17022 8676
rect 7258 8188 7322 8192
rect 7258 8132 7262 8188
rect 7262 8132 7318 8188
rect 7318 8132 7322 8188
rect 7258 8128 7322 8132
rect 7338 8188 7402 8192
rect 7338 8132 7342 8188
rect 7342 8132 7398 8188
rect 7398 8132 7402 8188
rect 7338 8128 7402 8132
rect 7418 8188 7482 8192
rect 7418 8132 7422 8188
rect 7422 8132 7478 8188
rect 7478 8132 7482 8188
rect 7418 8128 7482 8132
rect 7498 8188 7562 8192
rect 7498 8132 7502 8188
rect 7502 8132 7558 8188
rect 7558 8132 7562 8188
rect 7498 8128 7562 8132
rect 13565 8188 13629 8192
rect 13565 8132 13569 8188
rect 13569 8132 13625 8188
rect 13625 8132 13629 8188
rect 13565 8128 13629 8132
rect 13645 8188 13709 8192
rect 13645 8132 13649 8188
rect 13649 8132 13705 8188
rect 13705 8132 13709 8188
rect 13645 8128 13709 8132
rect 13725 8188 13789 8192
rect 13725 8132 13729 8188
rect 13729 8132 13785 8188
rect 13785 8132 13789 8188
rect 13725 8128 13789 8132
rect 13805 8188 13869 8192
rect 13805 8132 13809 8188
rect 13809 8132 13865 8188
rect 13865 8132 13869 8188
rect 13805 8128 13869 8132
rect 4105 7644 4169 7648
rect 4105 7588 4109 7644
rect 4109 7588 4165 7644
rect 4165 7588 4169 7644
rect 4105 7584 4169 7588
rect 4185 7644 4249 7648
rect 4185 7588 4189 7644
rect 4189 7588 4245 7644
rect 4245 7588 4249 7644
rect 4185 7584 4249 7588
rect 4265 7644 4329 7648
rect 4265 7588 4269 7644
rect 4269 7588 4325 7644
rect 4325 7588 4329 7644
rect 4265 7584 4329 7588
rect 4345 7644 4409 7648
rect 4345 7588 4349 7644
rect 4349 7588 4405 7644
rect 4405 7588 4409 7644
rect 4345 7584 4409 7588
rect 10411 7644 10475 7648
rect 10411 7588 10415 7644
rect 10415 7588 10471 7644
rect 10471 7588 10475 7644
rect 10411 7584 10475 7588
rect 10491 7644 10555 7648
rect 10491 7588 10495 7644
rect 10495 7588 10551 7644
rect 10551 7588 10555 7644
rect 10491 7584 10555 7588
rect 10571 7644 10635 7648
rect 10571 7588 10575 7644
rect 10575 7588 10631 7644
rect 10631 7588 10635 7644
rect 10571 7584 10635 7588
rect 10651 7644 10715 7648
rect 10651 7588 10655 7644
rect 10655 7588 10711 7644
rect 10711 7588 10715 7644
rect 10651 7584 10715 7588
rect 16718 7644 16782 7648
rect 16718 7588 16722 7644
rect 16722 7588 16778 7644
rect 16778 7588 16782 7644
rect 16718 7584 16782 7588
rect 16798 7644 16862 7648
rect 16798 7588 16802 7644
rect 16802 7588 16858 7644
rect 16858 7588 16862 7644
rect 16798 7584 16862 7588
rect 16878 7644 16942 7648
rect 16878 7588 16882 7644
rect 16882 7588 16938 7644
rect 16938 7588 16942 7644
rect 16878 7584 16942 7588
rect 16958 7644 17022 7648
rect 16958 7588 16962 7644
rect 16962 7588 17018 7644
rect 17018 7588 17022 7644
rect 16958 7584 17022 7588
rect 7258 7100 7322 7104
rect 7258 7044 7262 7100
rect 7262 7044 7318 7100
rect 7318 7044 7322 7100
rect 7258 7040 7322 7044
rect 7338 7100 7402 7104
rect 7338 7044 7342 7100
rect 7342 7044 7398 7100
rect 7398 7044 7402 7100
rect 7338 7040 7402 7044
rect 7418 7100 7482 7104
rect 7418 7044 7422 7100
rect 7422 7044 7478 7100
rect 7478 7044 7482 7100
rect 7418 7040 7482 7044
rect 7498 7100 7562 7104
rect 7498 7044 7502 7100
rect 7502 7044 7558 7100
rect 7558 7044 7562 7100
rect 7498 7040 7562 7044
rect 13565 7100 13629 7104
rect 13565 7044 13569 7100
rect 13569 7044 13625 7100
rect 13625 7044 13629 7100
rect 13565 7040 13629 7044
rect 13645 7100 13709 7104
rect 13645 7044 13649 7100
rect 13649 7044 13705 7100
rect 13705 7044 13709 7100
rect 13645 7040 13709 7044
rect 13725 7100 13789 7104
rect 13725 7044 13729 7100
rect 13729 7044 13785 7100
rect 13785 7044 13789 7100
rect 13725 7040 13789 7044
rect 13805 7100 13869 7104
rect 13805 7044 13809 7100
rect 13809 7044 13865 7100
rect 13865 7044 13869 7100
rect 13805 7040 13869 7044
rect 4105 6556 4169 6560
rect 4105 6500 4109 6556
rect 4109 6500 4165 6556
rect 4165 6500 4169 6556
rect 4105 6496 4169 6500
rect 4185 6556 4249 6560
rect 4185 6500 4189 6556
rect 4189 6500 4245 6556
rect 4245 6500 4249 6556
rect 4185 6496 4249 6500
rect 4265 6556 4329 6560
rect 4265 6500 4269 6556
rect 4269 6500 4325 6556
rect 4325 6500 4329 6556
rect 4265 6496 4329 6500
rect 4345 6556 4409 6560
rect 4345 6500 4349 6556
rect 4349 6500 4405 6556
rect 4405 6500 4409 6556
rect 4345 6496 4409 6500
rect 10411 6556 10475 6560
rect 10411 6500 10415 6556
rect 10415 6500 10471 6556
rect 10471 6500 10475 6556
rect 10411 6496 10475 6500
rect 10491 6556 10555 6560
rect 10491 6500 10495 6556
rect 10495 6500 10551 6556
rect 10551 6500 10555 6556
rect 10491 6496 10555 6500
rect 10571 6556 10635 6560
rect 10571 6500 10575 6556
rect 10575 6500 10631 6556
rect 10631 6500 10635 6556
rect 10571 6496 10635 6500
rect 10651 6556 10715 6560
rect 10651 6500 10655 6556
rect 10655 6500 10711 6556
rect 10711 6500 10715 6556
rect 10651 6496 10715 6500
rect 16718 6556 16782 6560
rect 16718 6500 16722 6556
rect 16722 6500 16778 6556
rect 16778 6500 16782 6556
rect 16718 6496 16782 6500
rect 16798 6556 16862 6560
rect 16798 6500 16802 6556
rect 16802 6500 16858 6556
rect 16858 6500 16862 6556
rect 16798 6496 16862 6500
rect 16878 6556 16942 6560
rect 16878 6500 16882 6556
rect 16882 6500 16938 6556
rect 16938 6500 16942 6556
rect 16878 6496 16942 6500
rect 16958 6556 17022 6560
rect 16958 6500 16962 6556
rect 16962 6500 17018 6556
rect 17018 6500 17022 6556
rect 16958 6496 17022 6500
rect 7258 6012 7322 6016
rect 7258 5956 7262 6012
rect 7262 5956 7318 6012
rect 7318 5956 7322 6012
rect 7258 5952 7322 5956
rect 7338 6012 7402 6016
rect 7338 5956 7342 6012
rect 7342 5956 7398 6012
rect 7398 5956 7402 6012
rect 7338 5952 7402 5956
rect 7418 6012 7482 6016
rect 7418 5956 7422 6012
rect 7422 5956 7478 6012
rect 7478 5956 7482 6012
rect 7418 5952 7482 5956
rect 7498 6012 7562 6016
rect 7498 5956 7502 6012
rect 7502 5956 7558 6012
rect 7558 5956 7562 6012
rect 7498 5952 7562 5956
rect 13565 6012 13629 6016
rect 13565 5956 13569 6012
rect 13569 5956 13625 6012
rect 13625 5956 13629 6012
rect 13565 5952 13629 5956
rect 13645 6012 13709 6016
rect 13645 5956 13649 6012
rect 13649 5956 13705 6012
rect 13705 5956 13709 6012
rect 13645 5952 13709 5956
rect 13725 6012 13789 6016
rect 13725 5956 13729 6012
rect 13729 5956 13785 6012
rect 13785 5956 13789 6012
rect 13725 5952 13789 5956
rect 13805 6012 13869 6016
rect 13805 5956 13809 6012
rect 13809 5956 13865 6012
rect 13865 5956 13869 6012
rect 13805 5952 13869 5956
rect 4105 5468 4169 5472
rect 4105 5412 4109 5468
rect 4109 5412 4165 5468
rect 4165 5412 4169 5468
rect 4105 5408 4169 5412
rect 4185 5468 4249 5472
rect 4185 5412 4189 5468
rect 4189 5412 4245 5468
rect 4245 5412 4249 5468
rect 4185 5408 4249 5412
rect 4265 5468 4329 5472
rect 4265 5412 4269 5468
rect 4269 5412 4325 5468
rect 4325 5412 4329 5468
rect 4265 5408 4329 5412
rect 4345 5468 4409 5472
rect 4345 5412 4349 5468
rect 4349 5412 4405 5468
rect 4405 5412 4409 5468
rect 4345 5408 4409 5412
rect 10411 5468 10475 5472
rect 10411 5412 10415 5468
rect 10415 5412 10471 5468
rect 10471 5412 10475 5468
rect 10411 5408 10475 5412
rect 10491 5468 10555 5472
rect 10491 5412 10495 5468
rect 10495 5412 10551 5468
rect 10551 5412 10555 5468
rect 10491 5408 10555 5412
rect 10571 5468 10635 5472
rect 10571 5412 10575 5468
rect 10575 5412 10631 5468
rect 10631 5412 10635 5468
rect 10571 5408 10635 5412
rect 10651 5468 10715 5472
rect 10651 5412 10655 5468
rect 10655 5412 10711 5468
rect 10711 5412 10715 5468
rect 10651 5408 10715 5412
rect 16718 5468 16782 5472
rect 16718 5412 16722 5468
rect 16722 5412 16778 5468
rect 16778 5412 16782 5468
rect 16718 5408 16782 5412
rect 16798 5468 16862 5472
rect 16798 5412 16802 5468
rect 16802 5412 16858 5468
rect 16858 5412 16862 5468
rect 16798 5408 16862 5412
rect 16878 5468 16942 5472
rect 16878 5412 16882 5468
rect 16882 5412 16938 5468
rect 16938 5412 16942 5468
rect 16878 5408 16942 5412
rect 16958 5468 17022 5472
rect 16958 5412 16962 5468
rect 16962 5412 17018 5468
rect 17018 5412 17022 5468
rect 16958 5408 17022 5412
rect 7258 4924 7322 4928
rect 7258 4868 7262 4924
rect 7262 4868 7318 4924
rect 7318 4868 7322 4924
rect 7258 4864 7322 4868
rect 7338 4924 7402 4928
rect 7338 4868 7342 4924
rect 7342 4868 7398 4924
rect 7398 4868 7402 4924
rect 7338 4864 7402 4868
rect 7418 4924 7482 4928
rect 7418 4868 7422 4924
rect 7422 4868 7478 4924
rect 7478 4868 7482 4924
rect 7418 4864 7482 4868
rect 7498 4924 7562 4928
rect 7498 4868 7502 4924
rect 7502 4868 7558 4924
rect 7558 4868 7562 4924
rect 7498 4864 7562 4868
rect 13565 4924 13629 4928
rect 13565 4868 13569 4924
rect 13569 4868 13625 4924
rect 13625 4868 13629 4924
rect 13565 4864 13629 4868
rect 13645 4924 13709 4928
rect 13645 4868 13649 4924
rect 13649 4868 13705 4924
rect 13705 4868 13709 4924
rect 13645 4864 13709 4868
rect 13725 4924 13789 4928
rect 13725 4868 13729 4924
rect 13729 4868 13785 4924
rect 13785 4868 13789 4924
rect 13725 4864 13789 4868
rect 13805 4924 13869 4928
rect 13805 4868 13809 4924
rect 13809 4868 13865 4924
rect 13865 4868 13869 4924
rect 13805 4864 13869 4868
rect 4105 4380 4169 4384
rect 4105 4324 4109 4380
rect 4109 4324 4165 4380
rect 4165 4324 4169 4380
rect 4105 4320 4169 4324
rect 4185 4380 4249 4384
rect 4185 4324 4189 4380
rect 4189 4324 4245 4380
rect 4245 4324 4249 4380
rect 4185 4320 4249 4324
rect 4265 4380 4329 4384
rect 4265 4324 4269 4380
rect 4269 4324 4325 4380
rect 4325 4324 4329 4380
rect 4265 4320 4329 4324
rect 4345 4380 4409 4384
rect 4345 4324 4349 4380
rect 4349 4324 4405 4380
rect 4405 4324 4409 4380
rect 4345 4320 4409 4324
rect 10411 4380 10475 4384
rect 10411 4324 10415 4380
rect 10415 4324 10471 4380
rect 10471 4324 10475 4380
rect 10411 4320 10475 4324
rect 10491 4380 10555 4384
rect 10491 4324 10495 4380
rect 10495 4324 10551 4380
rect 10551 4324 10555 4380
rect 10491 4320 10555 4324
rect 10571 4380 10635 4384
rect 10571 4324 10575 4380
rect 10575 4324 10631 4380
rect 10631 4324 10635 4380
rect 10571 4320 10635 4324
rect 10651 4380 10715 4384
rect 10651 4324 10655 4380
rect 10655 4324 10711 4380
rect 10711 4324 10715 4380
rect 10651 4320 10715 4324
rect 16718 4380 16782 4384
rect 16718 4324 16722 4380
rect 16722 4324 16778 4380
rect 16778 4324 16782 4380
rect 16718 4320 16782 4324
rect 16798 4380 16862 4384
rect 16798 4324 16802 4380
rect 16802 4324 16858 4380
rect 16858 4324 16862 4380
rect 16798 4320 16862 4324
rect 16878 4380 16942 4384
rect 16878 4324 16882 4380
rect 16882 4324 16938 4380
rect 16938 4324 16942 4380
rect 16878 4320 16942 4324
rect 16958 4380 17022 4384
rect 16958 4324 16962 4380
rect 16962 4324 17018 4380
rect 17018 4324 17022 4380
rect 16958 4320 17022 4324
rect 7258 3836 7322 3840
rect 7258 3780 7262 3836
rect 7262 3780 7318 3836
rect 7318 3780 7322 3836
rect 7258 3776 7322 3780
rect 7338 3836 7402 3840
rect 7338 3780 7342 3836
rect 7342 3780 7398 3836
rect 7398 3780 7402 3836
rect 7338 3776 7402 3780
rect 7418 3836 7482 3840
rect 7418 3780 7422 3836
rect 7422 3780 7478 3836
rect 7478 3780 7482 3836
rect 7418 3776 7482 3780
rect 7498 3836 7562 3840
rect 7498 3780 7502 3836
rect 7502 3780 7558 3836
rect 7558 3780 7562 3836
rect 7498 3776 7562 3780
rect 13565 3836 13629 3840
rect 13565 3780 13569 3836
rect 13569 3780 13625 3836
rect 13625 3780 13629 3836
rect 13565 3776 13629 3780
rect 13645 3836 13709 3840
rect 13645 3780 13649 3836
rect 13649 3780 13705 3836
rect 13705 3780 13709 3836
rect 13645 3776 13709 3780
rect 13725 3836 13789 3840
rect 13725 3780 13729 3836
rect 13729 3780 13785 3836
rect 13785 3780 13789 3836
rect 13725 3776 13789 3780
rect 13805 3836 13869 3840
rect 13805 3780 13809 3836
rect 13809 3780 13865 3836
rect 13865 3780 13869 3836
rect 13805 3776 13869 3780
rect 4105 3292 4169 3296
rect 4105 3236 4109 3292
rect 4109 3236 4165 3292
rect 4165 3236 4169 3292
rect 4105 3232 4169 3236
rect 4185 3292 4249 3296
rect 4185 3236 4189 3292
rect 4189 3236 4245 3292
rect 4245 3236 4249 3292
rect 4185 3232 4249 3236
rect 4265 3292 4329 3296
rect 4265 3236 4269 3292
rect 4269 3236 4325 3292
rect 4325 3236 4329 3292
rect 4265 3232 4329 3236
rect 4345 3292 4409 3296
rect 4345 3236 4349 3292
rect 4349 3236 4405 3292
rect 4405 3236 4409 3292
rect 4345 3232 4409 3236
rect 10411 3292 10475 3296
rect 10411 3236 10415 3292
rect 10415 3236 10471 3292
rect 10471 3236 10475 3292
rect 10411 3232 10475 3236
rect 10491 3292 10555 3296
rect 10491 3236 10495 3292
rect 10495 3236 10551 3292
rect 10551 3236 10555 3292
rect 10491 3232 10555 3236
rect 10571 3292 10635 3296
rect 10571 3236 10575 3292
rect 10575 3236 10631 3292
rect 10631 3236 10635 3292
rect 10571 3232 10635 3236
rect 10651 3292 10715 3296
rect 10651 3236 10655 3292
rect 10655 3236 10711 3292
rect 10711 3236 10715 3292
rect 10651 3232 10715 3236
rect 16718 3292 16782 3296
rect 16718 3236 16722 3292
rect 16722 3236 16778 3292
rect 16778 3236 16782 3292
rect 16718 3232 16782 3236
rect 16798 3292 16862 3296
rect 16798 3236 16802 3292
rect 16802 3236 16858 3292
rect 16858 3236 16862 3292
rect 16798 3232 16862 3236
rect 16878 3292 16942 3296
rect 16878 3236 16882 3292
rect 16882 3236 16938 3292
rect 16938 3236 16942 3292
rect 16878 3232 16942 3236
rect 16958 3292 17022 3296
rect 16958 3236 16962 3292
rect 16962 3236 17018 3292
rect 17018 3236 17022 3292
rect 16958 3232 17022 3236
rect 7258 2748 7322 2752
rect 7258 2692 7262 2748
rect 7262 2692 7318 2748
rect 7318 2692 7322 2748
rect 7258 2688 7322 2692
rect 7338 2748 7402 2752
rect 7338 2692 7342 2748
rect 7342 2692 7398 2748
rect 7398 2692 7402 2748
rect 7338 2688 7402 2692
rect 7418 2748 7482 2752
rect 7418 2692 7422 2748
rect 7422 2692 7478 2748
rect 7478 2692 7482 2748
rect 7418 2688 7482 2692
rect 7498 2748 7562 2752
rect 7498 2692 7502 2748
rect 7502 2692 7558 2748
rect 7558 2692 7562 2748
rect 7498 2688 7562 2692
rect 13565 2748 13629 2752
rect 13565 2692 13569 2748
rect 13569 2692 13625 2748
rect 13625 2692 13629 2748
rect 13565 2688 13629 2692
rect 13645 2748 13709 2752
rect 13645 2692 13649 2748
rect 13649 2692 13705 2748
rect 13705 2692 13709 2748
rect 13645 2688 13709 2692
rect 13725 2748 13789 2752
rect 13725 2692 13729 2748
rect 13729 2692 13785 2748
rect 13785 2692 13789 2748
rect 13725 2688 13789 2692
rect 13805 2748 13869 2752
rect 13805 2692 13809 2748
rect 13809 2692 13865 2748
rect 13865 2692 13869 2748
rect 13805 2688 13869 2692
rect 4105 2204 4169 2208
rect 4105 2148 4109 2204
rect 4109 2148 4165 2204
rect 4165 2148 4169 2204
rect 4105 2144 4169 2148
rect 4185 2204 4249 2208
rect 4185 2148 4189 2204
rect 4189 2148 4245 2204
rect 4245 2148 4249 2204
rect 4185 2144 4249 2148
rect 4265 2204 4329 2208
rect 4265 2148 4269 2204
rect 4269 2148 4325 2204
rect 4325 2148 4329 2204
rect 4265 2144 4329 2148
rect 4345 2204 4409 2208
rect 4345 2148 4349 2204
rect 4349 2148 4405 2204
rect 4405 2148 4409 2204
rect 4345 2144 4409 2148
rect 10411 2204 10475 2208
rect 10411 2148 10415 2204
rect 10415 2148 10471 2204
rect 10471 2148 10475 2204
rect 10411 2144 10475 2148
rect 10491 2204 10555 2208
rect 10491 2148 10495 2204
rect 10495 2148 10551 2204
rect 10551 2148 10555 2204
rect 10491 2144 10555 2148
rect 10571 2204 10635 2208
rect 10571 2148 10575 2204
rect 10575 2148 10631 2204
rect 10631 2148 10635 2204
rect 10571 2144 10635 2148
rect 10651 2204 10715 2208
rect 10651 2148 10655 2204
rect 10655 2148 10711 2204
rect 10711 2148 10715 2204
rect 10651 2144 10715 2148
rect 16718 2204 16782 2208
rect 16718 2148 16722 2204
rect 16722 2148 16778 2204
rect 16778 2148 16782 2204
rect 16718 2144 16782 2148
rect 16798 2204 16862 2208
rect 16798 2148 16802 2204
rect 16802 2148 16858 2204
rect 16858 2148 16862 2204
rect 16798 2144 16862 2148
rect 16878 2204 16942 2208
rect 16878 2148 16882 2204
rect 16882 2148 16938 2204
rect 16938 2148 16942 2204
rect 16878 2144 16942 2148
rect 16958 2204 17022 2208
rect 16958 2148 16962 2204
rect 16962 2148 17018 2204
rect 17018 2148 17022 2204
rect 16958 2144 17022 2148
<< metal4 >>
rect 4097 18528 4417 18544
rect 4097 18464 4105 18528
rect 4169 18464 4185 18528
rect 4249 18464 4265 18528
rect 4329 18464 4345 18528
rect 4409 18464 4417 18528
rect 4097 17440 4417 18464
rect 4097 17376 4105 17440
rect 4169 17376 4185 17440
rect 4249 17376 4265 17440
rect 4329 17376 4345 17440
rect 4409 17376 4417 17440
rect 4097 16352 4417 17376
rect 4097 16288 4105 16352
rect 4169 16288 4185 16352
rect 4249 16288 4265 16352
rect 4329 16288 4345 16352
rect 4409 16288 4417 16352
rect 4097 15264 4417 16288
rect 4097 15200 4105 15264
rect 4169 15200 4185 15264
rect 4249 15200 4265 15264
rect 4329 15200 4345 15264
rect 4409 15200 4417 15264
rect 4097 14176 4417 15200
rect 4097 14112 4105 14176
rect 4169 14112 4185 14176
rect 4249 14112 4265 14176
rect 4329 14112 4345 14176
rect 4409 14112 4417 14176
rect 4097 13088 4417 14112
rect 4097 13024 4105 13088
rect 4169 13024 4185 13088
rect 4249 13024 4265 13088
rect 4329 13024 4345 13088
rect 4409 13024 4417 13088
rect 4097 12000 4417 13024
rect 4097 11936 4105 12000
rect 4169 11936 4185 12000
rect 4249 11936 4265 12000
rect 4329 11936 4345 12000
rect 4409 11936 4417 12000
rect 4097 10912 4417 11936
rect 4097 10848 4105 10912
rect 4169 10848 4185 10912
rect 4249 10848 4265 10912
rect 4329 10848 4345 10912
rect 4409 10848 4417 10912
rect 4097 9824 4417 10848
rect 4097 9760 4105 9824
rect 4169 9760 4185 9824
rect 4249 9760 4265 9824
rect 4329 9760 4345 9824
rect 4409 9760 4417 9824
rect 4097 8736 4417 9760
rect 4097 8672 4105 8736
rect 4169 8672 4185 8736
rect 4249 8672 4265 8736
rect 4329 8672 4345 8736
rect 4409 8672 4417 8736
rect 4097 7648 4417 8672
rect 4097 7584 4105 7648
rect 4169 7584 4185 7648
rect 4249 7584 4265 7648
rect 4329 7584 4345 7648
rect 4409 7584 4417 7648
rect 4097 6560 4417 7584
rect 4097 6496 4105 6560
rect 4169 6496 4185 6560
rect 4249 6496 4265 6560
rect 4329 6496 4345 6560
rect 4409 6496 4417 6560
rect 4097 5472 4417 6496
rect 4097 5408 4105 5472
rect 4169 5408 4185 5472
rect 4249 5408 4265 5472
rect 4329 5408 4345 5472
rect 4409 5408 4417 5472
rect 4097 4384 4417 5408
rect 4097 4320 4105 4384
rect 4169 4320 4185 4384
rect 4249 4320 4265 4384
rect 4329 4320 4345 4384
rect 4409 4320 4417 4384
rect 4097 3296 4417 4320
rect 4097 3232 4105 3296
rect 4169 3232 4185 3296
rect 4249 3232 4265 3296
rect 4329 3232 4345 3296
rect 4409 3232 4417 3296
rect 4097 2208 4417 3232
rect 4097 2144 4105 2208
rect 4169 2144 4185 2208
rect 4249 2144 4265 2208
rect 4329 2144 4345 2208
rect 4409 2144 4417 2208
rect 4097 2128 4417 2144
rect 7250 17984 7570 18544
rect 7250 17920 7258 17984
rect 7322 17920 7338 17984
rect 7402 17920 7418 17984
rect 7482 17920 7498 17984
rect 7562 17920 7570 17984
rect 7250 16896 7570 17920
rect 7250 16832 7258 16896
rect 7322 16832 7338 16896
rect 7402 16832 7418 16896
rect 7482 16832 7498 16896
rect 7562 16832 7570 16896
rect 7250 15808 7570 16832
rect 7250 15744 7258 15808
rect 7322 15744 7338 15808
rect 7402 15744 7418 15808
rect 7482 15744 7498 15808
rect 7562 15744 7570 15808
rect 7250 14720 7570 15744
rect 7250 14656 7258 14720
rect 7322 14656 7338 14720
rect 7402 14656 7418 14720
rect 7482 14656 7498 14720
rect 7562 14656 7570 14720
rect 7250 13632 7570 14656
rect 7250 13568 7258 13632
rect 7322 13568 7338 13632
rect 7402 13568 7418 13632
rect 7482 13568 7498 13632
rect 7562 13568 7570 13632
rect 7250 12544 7570 13568
rect 7250 12480 7258 12544
rect 7322 12480 7338 12544
rect 7402 12480 7418 12544
rect 7482 12480 7498 12544
rect 7562 12480 7570 12544
rect 7250 11456 7570 12480
rect 7250 11392 7258 11456
rect 7322 11392 7338 11456
rect 7402 11392 7418 11456
rect 7482 11392 7498 11456
rect 7562 11392 7570 11456
rect 7250 10368 7570 11392
rect 7250 10304 7258 10368
rect 7322 10304 7338 10368
rect 7402 10304 7418 10368
rect 7482 10304 7498 10368
rect 7562 10304 7570 10368
rect 7250 9280 7570 10304
rect 7250 9216 7258 9280
rect 7322 9216 7338 9280
rect 7402 9216 7418 9280
rect 7482 9216 7498 9280
rect 7562 9216 7570 9280
rect 7250 8192 7570 9216
rect 7250 8128 7258 8192
rect 7322 8128 7338 8192
rect 7402 8128 7418 8192
rect 7482 8128 7498 8192
rect 7562 8128 7570 8192
rect 7250 7104 7570 8128
rect 7250 7040 7258 7104
rect 7322 7040 7338 7104
rect 7402 7040 7418 7104
rect 7482 7040 7498 7104
rect 7562 7040 7570 7104
rect 7250 6016 7570 7040
rect 7250 5952 7258 6016
rect 7322 5952 7338 6016
rect 7402 5952 7418 6016
rect 7482 5952 7498 6016
rect 7562 5952 7570 6016
rect 7250 4928 7570 5952
rect 7250 4864 7258 4928
rect 7322 4864 7338 4928
rect 7402 4864 7418 4928
rect 7482 4864 7498 4928
rect 7562 4864 7570 4928
rect 7250 3840 7570 4864
rect 7250 3776 7258 3840
rect 7322 3776 7338 3840
rect 7402 3776 7418 3840
rect 7482 3776 7498 3840
rect 7562 3776 7570 3840
rect 7250 2752 7570 3776
rect 7250 2688 7258 2752
rect 7322 2688 7338 2752
rect 7402 2688 7418 2752
rect 7482 2688 7498 2752
rect 7562 2688 7570 2752
rect 7250 2128 7570 2688
rect 10403 18528 10723 18544
rect 10403 18464 10411 18528
rect 10475 18464 10491 18528
rect 10555 18464 10571 18528
rect 10635 18464 10651 18528
rect 10715 18464 10723 18528
rect 10403 17440 10723 18464
rect 10403 17376 10411 17440
rect 10475 17376 10491 17440
rect 10555 17376 10571 17440
rect 10635 17376 10651 17440
rect 10715 17376 10723 17440
rect 10403 16352 10723 17376
rect 10403 16288 10411 16352
rect 10475 16288 10491 16352
rect 10555 16288 10571 16352
rect 10635 16288 10651 16352
rect 10715 16288 10723 16352
rect 10403 15264 10723 16288
rect 10403 15200 10411 15264
rect 10475 15200 10491 15264
rect 10555 15200 10571 15264
rect 10635 15200 10651 15264
rect 10715 15200 10723 15264
rect 10403 14176 10723 15200
rect 10403 14112 10411 14176
rect 10475 14112 10491 14176
rect 10555 14112 10571 14176
rect 10635 14112 10651 14176
rect 10715 14112 10723 14176
rect 10403 13088 10723 14112
rect 10403 13024 10411 13088
rect 10475 13024 10491 13088
rect 10555 13024 10571 13088
rect 10635 13024 10651 13088
rect 10715 13024 10723 13088
rect 10403 12000 10723 13024
rect 10403 11936 10411 12000
rect 10475 11936 10491 12000
rect 10555 11936 10571 12000
rect 10635 11936 10651 12000
rect 10715 11936 10723 12000
rect 10403 10912 10723 11936
rect 10403 10848 10411 10912
rect 10475 10848 10491 10912
rect 10555 10848 10571 10912
rect 10635 10848 10651 10912
rect 10715 10848 10723 10912
rect 10403 9824 10723 10848
rect 10403 9760 10411 9824
rect 10475 9760 10491 9824
rect 10555 9760 10571 9824
rect 10635 9760 10651 9824
rect 10715 9760 10723 9824
rect 10403 8736 10723 9760
rect 10403 8672 10411 8736
rect 10475 8672 10491 8736
rect 10555 8672 10571 8736
rect 10635 8672 10651 8736
rect 10715 8672 10723 8736
rect 10403 7648 10723 8672
rect 10403 7584 10411 7648
rect 10475 7584 10491 7648
rect 10555 7584 10571 7648
rect 10635 7584 10651 7648
rect 10715 7584 10723 7648
rect 10403 6560 10723 7584
rect 10403 6496 10411 6560
rect 10475 6496 10491 6560
rect 10555 6496 10571 6560
rect 10635 6496 10651 6560
rect 10715 6496 10723 6560
rect 10403 5472 10723 6496
rect 10403 5408 10411 5472
rect 10475 5408 10491 5472
rect 10555 5408 10571 5472
rect 10635 5408 10651 5472
rect 10715 5408 10723 5472
rect 10403 4384 10723 5408
rect 10403 4320 10411 4384
rect 10475 4320 10491 4384
rect 10555 4320 10571 4384
rect 10635 4320 10651 4384
rect 10715 4320 10723 4384
rect 10403 3296 10723 4320
rect 10403 3232 10411 3296
rect 10475 3232 10491 3296
rect 10555 3232 10571 3296
rect 10635 3232 10651 3296
rect 10715 3232 10723 3296
rect 10403 2208 10723 3232
rect 10403 2144 10411 2208
rect 10475 2144 10491 2208
rect 10555 2144 10571 2208
rect 10635 2144 10651 2208
rect 10715 2144 10723 2208
rect 10403 2128 10723 2144
rect 13557 17984 13877 18544
rect 13557 17920 13565 17984
rect 13629 17920 13645 17984
rect 13709 17920 13725 17984
rect 13789 17920 13805 17984
rect 13869 17920 13877 17984
rect 13557 16896 13877 17920
rect 13557 16832 13565 16896
rect 13629 16832 13645 16896
rect 13709 16832 13725 16896
rect 13789 16832 13805 16896
rect 13869 16832 13877 16896
rect 13557 15808 13877 16832
rect 13557 15744 13565 15808
rect 13629 15744 13645 15808
rect 13709 15744 13725 15808
rect 13789 15744 13805 15808
rect 13869 15744 13877 15808
rect 13557 14720 13877 15744
rect 13557 14656 13565 14720
rect 13629 14656 13645 14720
rect 13709 14656 13725 14720
rect 13789 14656 13805 14720
rect 13869 14656 13877 14720
rect 13557 13632 13877 14656
rect 13557 13568 13565 13632
rect 13629 13568 13645 13632
rect 13709 13568 13725 13632
rect 13789 13568 13805 13632
rect 13869 13568 13877 13632
rect 13557 12544 13877 13568
rect 13557 12480 13565 12544
rect 13629 12480 13645 12544
rect 13709 12480 13725 12544
rect 13789 12480 13805 12544
rect 13869 12480 13877 12544
rect 13557 11456 13877 12480
rect 13557 11392 13565 11456
rect 13629 11392 13645 11456
rect 13709 11392 13725 11456
rect 13789 11392 13805 11456
rect 13869 11392 13877 11456
rect 13557 10368 13877 11392
rect 13557 10304 13565 10368
rect 13629 10304 13645 10368
rect 13709 10304 13725 10368
rect 13789 10304 13805 10368
rect 13869 10304 13877 10368
rect 13557 9280 13877 10304
rect 13557 9216 13565 9280
rect 13629 9216 13645 9280
rect 13709 9216 13725 9280
rect 13789 9216 13805 9280
rect 13869 9216 13877 9280
rect 13557 8192 13877 9216
rect 13557 8128 13565 8192
rect 13629 8128 13645 8192
rect 13709 8128 13725 8192
rect 13789 8128 13805 8192
rect 13869 8128 13877 8192
rect 13557 7104 13877 8128
rect 13557 7040 13565 7104
rect 13629 7040 13645 7104
rect 13709 7040 13725 7104
rect 13789 7040 13805 7104
rect 13869 7040 13877 7104
rect 13557 6016 13877 7040
rect 13557 5952 13565 6016
rect 13629 5952 13645 6016
rect 13709 5952 13725 6016
rect 13789 5952 13805 6016
rect 13869 5952 13877 6016
rect 13557 4928 13877 5952
rect 13557 4864 13565 4928
rect 13629 4864 13645 4928
rect 13709 4864 13725 4928
rect 13789 4864 13805 4928
rect 13869 4864 13877 4928
rect 13557 3840 13877 4864
rect 13557 3776 13565 3840
rect 13629 3776 13645 3840
rect 13709 3776 13725 3840
rect 13789 3776 13805 3840
rect 13869 3776 13877 3840
rect 13557 2752 13877 3776
rect 13557 2688 13565 2752
rect 13629 2688 13645 2752
rect 13709 2688 13725 2752
rect 13789 2688 13805 2752
rect 13869 2688 13877 2752
rect 13557 2128 13877 2688
rect 16710 18528 17030 18544
rect 16710 18464 16718 18528
rect 16782 18464 16798 18528
rect 16862 18464 16878 18528
rect 16942 18464 16958 18528
rect 17022 18464 17030 18528
rect 16710 17440 17030 18464
rect 16710 17376 16718 17440
rect 16782 17376 16798 17440
rect 16862 17376 16878 17440
rect 16942 17376 16958 17440
rect 17022 17376 17030 17440
rect 16710 16352 17030 17376
rect 16710 16288 16718 16352
rect 16782 16288 16798 16352
rect 16862 16288 16878 16352
rect 16942 16288 16958 16352
rect 17022 16288 17030 16352
rect 16710 15264 17030 16288
rect 16710 15200 16718 15264
rect 16782 15200 16798 15264
rect 16862 15200 16878 15264
rect 16942 15200 16958 15264
rect 17022 15200 17030 15264
rect 16710 14176 17030 15200
rect 16710 14112 16718 14176
rect 16782 14112 16798 14176
rect 16862 14112 16878 14176
rect 16942 14112 16958 14176
rect 17022 14112 17030 14176
rect 16710 13088 17030 14112
rect 16710 13024 16718 13088
rect 16782 13024 16798 13088
rect 16862 13024 16878 13088
rect 16942 13024 16958 13088
rect 17022 13024 17030 13088
rect 16710 12000 17030 13024
rect 16710 11936 16718 12000
rect 16782 11936 16798 12000
rect 16862 11936 16878 12000
rect 16942 11936 16958 12000
rect 17022 11936 17030 12000
rect 16710 10912 17030 11936
rect 16710 10848 16718 10912
rect 16782 10848 16798 10912
rect 16862 10848 16878 10912
rect 16942 10848 16958 10912
rect 17022 10848 17030 10912
rect 16710 9824 17030 10848
rect 16710 9760 16718 9824
rect 16782 9760 16798 9824
rect 16862 9760 16878 9824
rect 16942 9760 16958 9824
rect 17022 9760 17030 9824
rect 16710 8736 17030 9760
rect 16710 8672 16718 8736
rect 16782 8672 16798 8736
rect 16862 8672 16878 8736
rect 16942 8672 16958 8736
rect 17022 8672 17030 8736
rect 16710 7648 17030 8672
rect 16710 7584 16718 7648
rect 16782 7584 16798 7648
rect 16862 7584 16878 7648
rect 16942 7584 16958 7648
rect 17022 7584 17030 7648
rect 16710 6560 17030 7584
rect 16710 6496 16718 6560
rect 16782 6496 16798 6560
rect 16862 6496 16878 6560
rect 16942 6496 16958 6560
rect 17022 6496 17030 6560
rect 16710 5472 17030 6496
rect 16710 5408 16718 5472
rect 16782 5408 16798 5472
rect 16862 5408 16878 5472
rect 16942 5408 16958 5472
rect 17022 5408 17030 5472
rect 16710 4384 17030 5408
rect 16710 4320 16718 4384
rect 16782 4320 16798 4384
rect 16862 4320 16878 4384
rect 16942 4320 16958 4384
rect 17022 4320 17030 4384
rect 16710 3296 17030 4320
rect 16710 3232 16718 3296
rect 16782 3232 16798 3296
rect 16862 3232 16878 3296
rect 16942 3232 16958 3296
rect 17022 3232 17030 3296
rect 16710 2208 17030 3232
rect 16710 2144 16718 2208
rect 16782 2144 16798 2208
rect 16862 2144 16878 2208
rect 16942 2144 16958 2208
rect 17022 2144 17030 2208
rect 16710 2128 17030 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_7
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_19
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_60 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_43
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_55
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_1_67
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_73 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 130 592
use scs8hd_buf_2  _36_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_79
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_83
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_94 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_90
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_94
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_107
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_121
timestamp 1586364061
transform 1 0 12236 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_135
timestamp 1586364061
transform 1 0 13524 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_4  FILLER_1_133
timestamp 1586364061
transform 1 0 13340 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_139
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_143
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_150
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_166
timestamp 1586364061
transform 1 0 16376 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_156
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 17756 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 17756 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_167
timestamp 1586364061
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_177
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_18
timestamp 1586364061
transform 1 0 2760 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_79
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_12  FILLER_2_119
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13708 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_2_140
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_152
timestamp 1586364061
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 17756 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_175
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_12
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_24
timestamp 1586364061
transform 1 0 3312 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_48
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_60
timestamp 1586364061
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 774 592
use scs8hd_conb_1  _31_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_120
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_126
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_130
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_148
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_152
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16284 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_163
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 17756 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_167
timestamp 1586364061
transform 1 0 16468 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_7
timestamp 1586364061
transform 1 0 1748 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_conb_1  _33_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_96
timestamp 1586364061
transform 1 0 9936 0 -1 4896
box -38 -48 774 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_126
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_138
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_150
timestamp 1586364061
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 17756 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6256 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_55
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_58
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_79
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_87
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 314 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_130
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_142
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_166
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 17756 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_6
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_10
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_14
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_46
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_49
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_59
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_conb_1  _20_
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_6_71
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_6  FILLER_7_77
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10304 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_99
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_8  FILLER_6_103
timestamp 1586364061
transform 1 0 10580 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_7_106
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_120
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13708 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_131
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_139
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_143
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_151
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_163
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 17756 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 17756 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_16
timestamp 1586364061
transform 1 0 2576 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_28
timestamp 1586364061
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_50
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_74
timestamp 1586364061
transform 1 0 7912 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_8_86
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12144 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13708 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 17756 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 14076 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_145
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_163
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 17756 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_168
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_172
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_8
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_20
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_28
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_122
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_6  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_1  FILLER_10_160
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 17756 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_170
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_11_18
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_29
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_45
timestamp 1586364061
transform 1 0 5244 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_127
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_131
timestamp 1586364061
transform 1 0 13156 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_163
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 17756 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_172
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 590 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_11
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 406 592
use scs8hd_conb_1  _23_
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_158
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 17756 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_170
timestamp 1586364061
transform 1 0 16744 0 -1 9248
box -38 -48 774 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_23
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_17
timestamp 1586364061
transform 1 0 2668 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_29
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_141
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 130 592
use scs8hd_conb_1  _30_
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_144
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_13_165
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 17756 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 17756 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_177
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_175
timestamp 1586364061
transform 1 0 17204 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_14
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_18
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_31
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_42
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_46
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_155
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 17756 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_168
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_176
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_14
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_26
timestamp 1586364061
transform 1 0 3496 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 17756 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_167
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_175
timestamp 1586364061
transform 1 0 17204 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_12
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_17_24
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_38
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_42
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_45
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 406 592
use scs8hd_decap_4  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_139
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_144
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_148
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_154
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 17756 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_167
timestamp 1586364061
transform 1 0 16468 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 314 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_13
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_17
timestamp 1586364061
transform 1 0 2668 0 -1 12512
box -38 -48 1142 592
use scs8hd_conb_1  _21_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_29
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_35
timestamp 1586364061
transform 1 0 4324 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_57
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_69
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_81
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 17756 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_175
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_6
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_10
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_18
timestamp 1586364061
transform 1 0 2760 0 -1 13600
box -38 -48 1142 592
use scs8hd_conb_1  _35_
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_30
timestamp 1586364061
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_35
timestamp 1586364061
transform 1 0 4324 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_47
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_47
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_59
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_83
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_139
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_143
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 774 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16008 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_157
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_161
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_164
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 17756 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 17756 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_169
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_177
timestamp 1586364061
transform 1 0 17388 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_6
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_10
timestamp 1586364061
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_21_14
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_25
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_36
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_47
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_55
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_78
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_90
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_102
timestamp 1586364061
transform 1 0 10488 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 17756 0 1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_177
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_13
timestamp 1586364061
transform 1 0 2300 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_18
timestamp 1586364061
transform 1 0 2760 0 -1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_30
timestamp 1586364061
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_52
timestamp 1586364061
transform 1 0 5888 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_63
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_75
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_91
timestamp 1586364061
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 17756 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_17
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_21
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 866 592
use scs8hd_decap_6  FILLER_23_35
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _32_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_52
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_56
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_60
timestamp 1586364061
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_65
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 590 592
use scs8hd_conb_1  _19_
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_106
timestamp 1586364061
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_161
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_166
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 17756 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_170
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _18_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_35
timestamp 1586364061
transform 1 0 4324 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_47
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_62
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_81
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_110
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_122
timestamp 1586364061
transform 1 0 12328 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_134
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_146
timestamp 1586364061
transform 1 0 14536 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_158
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 17756 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_176
timestamp 1586364061
transform 1 0 17296 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_16
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_20
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_28
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_41
timestamp 1586364061
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_45
timestamp 1586364061
transform 1 0 5244 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_82
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_99
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_103
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_131
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_25_137
timestamp 1586364061
transform 1 0 13708 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_149
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_154
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 17756 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_167
timestamp 1586364061
transform 1 0 16468 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 866 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_20
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_24
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 590 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 4508 0 -1 16864
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_36
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_41
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_49
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 130 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_57
timestamp 1586364061
transform 1 0 6348 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_69
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_75
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_115
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_122
timestamp 1586364061
transform 1 0 12328 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_121
timestamp 1586364061
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_127
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_132
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_138
timestamp 1586364061
transform 1 0 13800 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_27_139
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 16284 0 1 16864
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_162
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 17756 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 17756 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_175
timestamp 1586364061
transform 1 0 17204 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_169
timestamp 1586364061
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_173
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_177
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 130 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5704 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_42
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_59
timestamp 1586364061
transform 1 0 6532 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  FILLER_28_71
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_78
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_101
timestamp 1586364061
transform 1 0 10396 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  FILLER_28_109
timestamp 1586364061
transform 1 0 11132 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_121
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 774 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_135
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_147
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 130 592
use scs8hd_conb_1  _22_
timestamp 1586364061
transform 1 0 15364 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_158
timestamp 1586364061
transform 1 0 15640 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 17756 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_169
timestamp 1586364061
transform 1 0 16652 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_177
timestamp 1586364061
transform 1 0 17388 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_6
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_10
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_17
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_21
timestamp 1586364061
transform 1 0 3036 0 1 17952
box -38 -48 774 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 3956 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_29
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_46
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_50
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 1142 592
use scs8hd_conb_1  _34_
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_63
timestamp 1586364061
transform 1 0 6900 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_67
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_78
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_82
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 774 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_90
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_94
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_99
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 12512 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_122
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_125
timestamp 1586364061
transform 1 0 12604 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_137
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_141
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_145
timestamp 1586364061
transform 1 0 14444 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_153
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_156
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 17756 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_168
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_176
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 222 592
<< labels >>
rlabel metal2 s 3054 0 3110 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 478 20583 534 21063 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 416 480 536 6 address[2]
port 2 nsew default input
rlabel metal3 s 0 1368 480 1488 6 address[3]
port 3 nsew default input
rlabel metal2 s 4342 0 4398 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 5538 0 5594 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 1398 20583 1454 21063 6 bottom_left_grid_pin_13_
port 6 nsew default input
rlabel metal3 s 0 4632 480 4752 6 bottom_right_grid_pin_11_
port 7 nsew default input
rlabel metal3 s 0 5584 480 5704 6 bottom_right_grid_pin_13_
port 8 nsew default input
rlabel metal3 s 0 6672 480 6792 6 bottom_right_grid_pin_15_
port 9 nsew default input
rlabel metal2 s 2410 20583 2466 21063 6 bottom_right_grid_pin_1_
port 10 nsew default input
rlabel metal2 s 6826 0 6882 480 6 bottom_right_grid_pin_3_
port 11 nsew default input
rlabel metal3 s 0 2456 480 2576 6 bottom_right_grid_pin_5_
port 12 nsew default input
rlabel metal3 s 18439 1232 18919 1352 6 bottom_right_grid_pin_7_
port 13 nsew default input
rlabel metal3 s 0 3544 480 3664 6 bottom_right_grid_pin_9_
port 14 nsew default input
rlabel metal3 s 18439 3816 18919 3936 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[1]
port 16 nsew default input
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[2]
port 17 nsew default input
rlabel metal3 s 18439 6400 18919 6520 6 chanx_left_in[3]
port 18 nsew default input
rlabel metal2 s 3422 20583 3478 21063 6 chanx_left_in[4]
port 19 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_left_in[5]
port 20 nsew default input
rlabel metal2 s 4434 20583 4490 21063 6 chanx_left_in[6]
port 21 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chanx_left_in[7]
port 22 nsew default input
rlabel metal3 s 0 10888 480 11008 6 chanx_left_in[8]
port 23 nsew default input
rlabel metal2 s 5446 20583 5502 21063 6 chanx_left_out[0]
port 24 nsew default tristate
rlabel metal2 s 6458 20583 6514 21063 6 chanx_left_out[1]
port 25 nsew default tristate
rlabel metal2 s 7378 20583 7434 21063 6 chanx_left_out[2]
port 26 nsew default tristate
rlabel metal2 s 8390 20583 8446 21063 6 chanx_left_out[3]
port 27 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_left_out[4]
port 28 nsew default tristate
rlabel metal2 s 9402 20583 9458 21063 6 chanx_left_out[5]
port 29 nsew default tristate
rlabel metal2 s 10414 20583 10470 21063 6 chanx_left_out[6]
port 30 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 chanx_left_out[7]
port 31 nsew default tristate
rlabel metal2 s 9402 0 9458 480 6 chanx_left_out[8]
port 32 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chany_bottom_in[0]
port 33 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[1]
port 34 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[2]
port 35 nsew default input
rlabel metal3 s 0 15104 480 15224 6 chany_bottom_in[3]
port 36 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_in[4]
port 37 nsew default input
rlabel metal2 s 11426 20583 11482 21063 6 chany_bottom_in[5]
port 38 nsew default input
rlabel metal3 s 18439 9120 18919 9240 6 chany_bottom_in[6]
port 39 nsew default input
rlabel metal2 s 14462 0 14518 480 6 chany_bottom_in[7]
port 40 nsew default input
rlabel metal2 s 12438 20583 12494 21063 6 chany_bottom_in[8]
port 41 nsew default input
rlabel metal3 s 0 16192 480 16312 6 chany_bottom_out[0]
port 42 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chany_bottom_out[1]
port 43 nsew default tristate
rlabel metal2 s 13358 20583 13414 21063 6 chany_bottom_out[2]
port 44 nsew default tristate
rlabel metal3 s 18439 11704 18919 11824 6 chany_bottom_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chany_bottom_out[4]
port 46 nsew default tristate
rlabel metal2 s 14370 20583 14426 21063 6 chany_bottom_out[5]
port 47 nsew default tristate
rlabel metal2 s 15382 20583 15438 21063 6 chany_bottom_out[6]
port 48 nsew default tristate
rlabel metal2 s 16394 20583 16450 21063 6 chany_bottom_out[7]
port 49 nsew default tristate
rlabel metal2 s 17406 20583 17462 21063 6 chany_bottom_out[8]
port 50 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 data_in
port 51 nsew default input
rlabel metal2 s 570 0 626 480 6 enable
port 52 nsew default input
rlabel metal3 s 18439 14288 18919 14408 6 left_bottom_grid_pin_12_
port 53 nsew default input
rlabel metal2 s 16946 0 17002 480 6 left_top_grid_pin_11_
port 54 nsew default input
rlabel metal2 s 18418 20583 18474 21063 6 left_top_grid_pin_13_
port 55 nsew default input
rlabel metal2 s 18234 0 18290 480 6 left_top_grid_pin_15_
port 56 nsew default input
rlabel metal3 s 0 19320 480 19440 6 left_top_grid_pin_1_
port 57 nsew default input
rlabel metal3 s 18439 17008 18919 17128 6 left_top_grid_pin_3_
port 58 nsew default input
rlabel metal2 s 15658 0 15714 480 6 left_top_grid_pin_5_
port 59 nsew default input
rlabel metal3 s 0 20408 480 20528 6 left_top_grid_pin_7_
port 60 nsew default input
rlabel metal3 s 18439 19592 18919 19712 6 left_top_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 4097 2128 4417 18544 6 vpwr
port 62 nsew default input
rlabel metal4 s 7250 2128 7570 18544 6 vgnd
port 63 nsew default input
<< end >>
