* NGSPICE file created from sb_1__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 D Q CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt sb_1__0_ ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11]
+ chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16]
+ chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2]
+ chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11]
+ chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16]
+ chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2]
+ chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7]
+ chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10] chanx_right_in[11]
+ chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15] chanx_right_in[16]
+ chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10] chanx_right_out[11]
+ chanx_right_out[12] chanx_right_out[13] chanx_right_out[14] chanx_right_out[15]
+ chanx_right_out[16] chanx_right_out[17] chanx_right_out[18] chanx_right_out[19]
+ chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5]
+ chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9] chany_top_in[0]
+ chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14]
+ chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19]
+ chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5]
+ chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0]
+ chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14]
+ chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19]
+ chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5]
+ chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9] left_bottom_grid_pin_11_
+ left_bottom_grid_pin_13_ left_bottom_grid_pin_15_ left_bottom_grid_pin_17_ left_bottom_grid_pin_1_
+ left_bottom_grid_pin_3_ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_
+ prog_clk right_bottom_grid_pin_11_ right_bottom_grid_pin_13_ right_bottom_grid_pin_15_
+ right_bottom_grid_pin_17_ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_
+ right_bottom_grid_pin_7_ right_bottom_grid_pin_9_ top_left_grid_pin_42_ top_left_grid_pin_43_
+ top_left_grid_pin_44_ top_left_grid_pin_45_ top_left_grid_pin_46_ top_left_grid_pin_47_
+ top_left_grid_pin_48_ top_left_grid_pin_49_ VPWR VGND
XFILLER_22_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_0.mux_l4_in_0_/S mux_right_track_2.mux_l1_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_9.mux_l4_in_0_/S mux_left_track_17.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_12_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_062_ chanx_right_in[12] chanx_left_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_8.mux_l1_in_0_/S mux_right_track_8.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_10.mux_l3_in_0_ mux_top_track_10.mux_l2_in_1_/X mux_top_track_10.mux_l2_in_0_/X
+ mux_top_track_10.mux_l3_in_0_/S mux_top_track_10.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_prog_clk clkbuf_2_2_0_prog_clk/X clkbuf_3_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
X_114_ _114_/A chany_top_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_045_ _045_/HI _045_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_10.mux_l2_in_1_ _030_/HI chanx_left_in[9] mux_top_track_10.mux_l2_in_0_/S
+ mux_top_track_10.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_028_ _028_/HI _028_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_061_ chanx_right_in[13] chanx_left_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_10.mux_l2_in_0_/S mux_top_track_10.mux_l3_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_4.mux_l4_in_0_/S mux_right_track_8.mux_l1_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l4_in_0_/X _071_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_113_ _113_/A chany_top_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_044_ _044_/HI _044_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_10.mux_l2_in_0_ chanx_right_in[19] mux_top_track_10.mux_l1_in_0_/X
+ mux_top_track_10.mux_l2_in_0_/S mux_top_track_10.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_3_ _028_/HI chanx_left_in[16] mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l3_in_0_/X _063_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_0.mux_l2_in_3_ _029_/HI chanx_left_in[2] mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l4_in_0_ mux_right_track_8.mux_l3_in_1_/X mux_right_track_8.mux_l3_in_0_/X
+ mux_right_track_8.mux_l4_in_0_/S mux_right_track_8.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_060_ chanx_right_in[14] chanx_left_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_10.mux_l1_in_0_/S mux_top_track_10.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ mux_top_track_0.mux_l4_in_0_/S mux_top_track_0.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_112_ _112_/A chany_top_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_043_ _043_/HI _043_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_8.mux_l3_in_1_ mux_right_track_8.mux_l2_in_3_/X mux_right_track_8.mux_l2_in_2_/X
+ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_1_/S mux_top_track_0.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_8.mux_l2_in_2_ chanx_left_in[6] right_bottom_grid_pin_17_ mux_right_track_8.mux_l2_in_0_/S
+ mux_right_track_8.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_0.mux_l2_in_2_ chanx_left_in[0] chanx_right_in[2] mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_22.mux_l2_in_0_ mux_top_track_22.mux_l1_in_1_/X mux_top_track_22.mux_l1_in_0_/X
+ mux_top_track_22.mux_l2_in_0_/S mux_top_track_22.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_10.mux_l1_in_0_ chanx_right_in[9] top_left_grid_pin_43_ mux_top_track_10.mux_l1_in_0_/S
+ mux_top_track_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_22.mux_l1_in_1_ _037_/HI chanx_left_in[17] mux_top_track_22.mux_l1_in_0_/S
+ mux_top_track_22.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_8.mux_l3_in_0_/S mux_top_track_10.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_111_ _111_/A chany_top_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_042_ _042_/HI _042_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_1_/S mux_top_track_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_16.mux_l1_in_0_/S mux_top_track_16.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_1_ right_bottom_grid_pin_9_ right_bottom_grid_pin_1_
+ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_0.mux_l2_in_1_ chanx_right_in[1] top_left_grid_pin_48_ mux_top_track_0.mux_l2_in_0_/S
+ mux_top_track_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_22.sky130_fd_sc_hd__buf_4_0_ mux_top_track_22.mux_l2_in_0_/X _104_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l2_in_0_/X _107_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_track_22.mux_l1_in_0_ chanx_right_in[17] top_left_grid_pin_49_ mux_top_track_22.mux_l1_in_0_/S
+ mux_top_track_22.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_110_ _110_/A chany_top_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_041_ _041_/HI _041_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_14.mux_l2_in_0_/S mux_top_track_16.mux_l1_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l4_in_0_/X _115_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_8.mux_l2_in_0_ chany_top_in[16] mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ top_left_grid_pin_46_ mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_0_/S mux_top_track_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_38.sky130_fd_sc_hd__buf_4_0_ mux_top_track_38.mux_l2_in_0_/X _096_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_040_ _040_/HI _040_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_28_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_8.mux_l1_in_0_ chany_top_in[9] chany_top_in[2] mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_prog_clk clkbuf_2_1_0_prog_clk/A clkbuf_3_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_0.mux_l1_in_0_ top_left_grid_pin_44_ top_left_grid_pin_42_ mux_top_track_0.mux_l1_in_0_/S
+ mux_top_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l4_in_0_/X _091_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_099_ chanx_left_in[11] chany_top_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l3_in_0_/X _079_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_6_ chanx_left_in[14] chanx_left_in[5] mux_right_track_4.mux_l1_in_6_/S
+ mux_right_track_4.mux_l1_in_6_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_2_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_ mux_left_track_1.mux_l3_in_1_/S mux_left_track_1.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_3_ _046_/HI left_bottom_grid_pin_15_ mux_left_track_3.mux_l2_in_1_/S
+ mux_left_track_3.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_098_ chanx_left_in[7] chany_top_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l4_in_0_ mux_left_track_3.mux_l3_in_1_/X mux_left_track_3.mux_l3_in_0_/X
+ mux_left_track_3.mux_l4_in_0_/S mux_left_track_3.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_4.mux_l1_in_5_ right_bottom_grid_pin_17_ right_bottom_grid_pin_15_
+ mux_right_track_4.mux_l1_in_6_/S mux_right_track_4.mux_l1_in_5_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_1_ mux_left_track_3.mux_l2_in_3_/X mux_left_track_3.mux_l2_in_2_/X
+ mux_left_track_3.mux_l3_in_0_/S mux_left_track_3.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l4_in_0_/X _073_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_1.mux_l2_in_3_/S mux_left_track_1.mux_l3_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l2_in_2_ left_bottom_grid_pin_11_ left_bottom_grid_pin_7_ mux_left_track_3.mux_l2_in_1_/S
+ mux_left_track_3.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l2_in_3_ _055_/HI mux_right_track_4.mux_l1_in_6_/X mux_right_track_4.mux_l2_in_2_/S
+ mux_right_track_4.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_097_ chanx_left_in[3] chany_top_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l3_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_4_ right_bottom_grid_pin_13_ right_bottom_grid_pin_11_
+ mux_right_track_4.mux_l1_in_6_/S mux_right_track_4.mux_l1_in_4_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S mux_left_track_3.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l4_in_0_ mux_right_track_4.mux_l3_in_1_/X mux_right_track_4.mux_l3_in_0_/X
+ mux_right_track_4.mux_l4_in_0_/S mux_right_track_4.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_1.mux_l1_in_0_/S mux_left_track_1.mux_l2_in_3_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l2_in_1_ left_bottom_grid_pin_3_ chanx_right_in[13] mux_left_track_3.mux_l2_in_1_/S
+ mux_left_track_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l3_in_1_ mux_right_track_4.mux_l2_in_3_/X mux_right_track_4.mux_l2_in_2_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l4_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_096_ _096_/A chany_top_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_0_/S mux_top_track_16.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_2_ mux_right_track_4.mux_l1_in_5_/X mux_right_track_4.mux_l1_in_4_/X
+ mux_right_track_4.mux_l2_in_2_/S mux_right_track_4.mux_l2_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_4.mux_l1_in_3_/S mux_top_track_4.mux_l2_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_079_ _079_/A chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_16.mux_l1_in_3_ _051_/HI chanx_left_in[17] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_20.mux_l1_in_1_/S mux_top_track_20.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_16.mux_l1_in_1_ _033_/HI chanx_left_in[13] mux_top_track_16.mux_l1_in_0_/S
+ mux_top_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_3_ right_bottom_grid_pin_9_ right_bottom_grid_pin_7_
+ mux_right_track_4.mux_l1_in_6_/S mux_right_track_4.mux_l1_in_3_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_16.mux_l3_in_0_ mux_right_track_16.mux_l2_in_1_/X mux_right_track_16.mux_l2_in_0_/X
+ mux_right_track_16.mux_l3_in_0_/S mux_right_track_16.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_32.mux_l3_in_0_/S mux_left_track_1.mux_l1_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ chanx_right_in[4] mux_left_track_3.mux_l1_in_0_/X mux_left_track_3.mux_l2_in_1_/S
+ mux_left_track_3.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_3_1_0_prog_clk clkbuf_3_1_0_prog_clk/A clkbuf_3_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_4.mux_l2_in_2_/S mux_right_track_4.mux_l3_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_16.mux_l2_in_1_ mux_right_track_16.mux_l1_in_3_/X mux_right_track_16.mux_l1_in_2_/X
+ mux_right_track_16.mux_l2_in_1_/S mux_right_track_16.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_095_ _095_/A chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_2_/S mux_right_track_4.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_2.mux_l3_in_0_/S mux_top_track_4.mux_l1_in_3_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_078_ chanx_left_in[16] chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_track_12.sky130_fd_sc_hd__buf_4_0_ mux_top_track_12.mux_l2_in_0_/X _109_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_right_track_16.mux_l1_in_2_ chanx_left_in[8] right_bottom_grid_pin_11_ mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.mux_l1_in_2_ right_bottom_grid_pin_5_ right_bottom_grid_pin_3_
+ mux_right_track_4.mux_l1_in_6_/S mux_right_track_4.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_0_ chanx_right_in[13] top_left_grid_pin_46_ mux_top_track_16.mux_l1_in_0_/S
+ mux_top_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_18.mux_l2_in_0_/S mux_top_track_20.mux_l1_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_6.mux_l1_in_3_ _041_/HI chanx_left_in[6] mux_top_track_6.mux_l1_in_3_/S
+ mux_top_track_6.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_4.mux_l1_in_6_/S mux_right_track_4.mux_l2_in_2_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[6] mux_left_track_3.mux_l1_in_0_/S
+ mux_left_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_1_/S mux_right_track_16.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_094_ _094_/A chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_track_6.mux_l3_in_0_ mux_top_track_6.mux_l2_in_1_/X mux_top_track_6.mux_l2_in_0_/X
+ mux_top_track_6.mux_l3_in_0_/S mux_top_track_6.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_2_/S mux_right_track_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_077_ chanx_left_in[17] chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_16.mux_l1_in_1_ right_bottom_grid_pin_3_ chany_top_in[17] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_6.mux_l2_in_1_ mux_top_track_6.mux_l1_in_3_/X mux_top_track_6.mux_l1_in_2_/X
+ mux_top_track_6.mux_l2_in_1_/S mux_top_track_6.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_1_ right_bottom_grid_pin_1_ chany_top_in[15] mux_right_track_4.mux_l1_in_6_/S
+ mux_right_track_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_6.mux_l1_in_2_ chanx_right_in[11] chanx_right_in[6] mux_top_track_6.mux_l1_in_3_/S
+ mux_top_track_6.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_2.mux_l4_in_0_/S mux_right_track_4.mux_l1_in_6_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_093_ _093_/A chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
X_076_ chanx_left_in[18] chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_0_ chany_top_in[10] chany_top_in[3] mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_6.mux_l2_in_0_ mux_top_track_6.mux_l1_in_1_/X mux_top_track_6.mux_l1_in_0_/X
+ mux_top_track_6.mux_l2_in_1_/S mux_top_track_6.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_4.mux_l1_in_0_ chany_top_in[8] chany_top_in[1] mux_right_track_4.mux_l1_in_6_/S
+ mux_right_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l4_in_0_/X _093_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_21_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ _059_/A chanx_left_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_6.sky130_fd_sc_hd__buf_4_0_ mux_top_track_6.mux_l3_in_0_/X _112_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_track_6.mux_l1_in_1_ top_left_grid_pin_49_ top_left_grid_pin_47_ mux_top_track_6.mux_l1_in_3_/S
+ mux_top_track_6.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_0_0_prog_clk clkbuf_3_1_0_prog_clk/A clkbuf_3_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_092_ chanx_left_in[2] chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_075_ _075_/A chanx_left_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l3_in_0_/X _087_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_058_ chanx_right_in[16] chanx_left_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_30_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_6.mux_l1_in_0_ top_left_grid_pin_45_ top_left_grid_pin_43_ mux_top_track_6.mux_l1_in_3_/S
+ mux_top_track_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l4_in_0_/X _075_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_24_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_091_ _091_/A chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_074_ _074_/A chanx_left_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_12.mux_l1_in_1_/S mux_top_track_12.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_18_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_057_ chanx_right_in[17] chanx_left_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_109_ _109_/A chany_top_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_26_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l2_in_3_ _049_/HI left_bottom_grid_pin_17_ mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_3_ _050_/HI chanx_left_in[12] mux_right_track_0.mux_l2_in_3_/S
+ mux_right_track_0.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_9.mux_l4_in_0_ mux_left_track_9.mux_l3_in_1_/X mux_left_track_9.mux_l3_in_0_/X
+ mux_left_track_9.mux_l4_in_0_/S mux_left_track_9.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
X_090_ chanx_left_in[4] chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l4_in_0_ mux_right_track_0.mux_l3_in_1_/X mux_right_track_0.mux_l3_in_0_/X
+ mux_right_track_0.mux_l4_in_0_/S mux_right_track_0.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_10.mux_l3_in_0_/S mux_top_track_12.mux_l1_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_073_ _073_/A chanx_left_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_056_ chanx_right_in[18] chanx_left_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_9.mux_l3_in_1_ mux_left_track_9.mux_l2_in_3_/X mux_left_track_9.mux_l2_in_2_/X
+ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l3_in_1_ mux_right_track_0.mux_l2_in_3_/X mux_right_track_0.mux_l2_in_2_/X
+ mux_right_track_0.mux_l3_in_1_/S mux_right_track_0.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_108_ _108_/A chany_top_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l1_in_3_ _044_/HI left_bottom_grid_pin_11_ mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_039_ _039_/HI _039_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_18.mux_l1_in_1_/S mux_top_track_18.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_27_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_9.mux_l2_in_2_ left_bottom_grid_pin_9_ left_bottom_grid_pin_1_ mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l2_in_2_ chanx_left_in[2] right_bottom_grid_pin_17_ mux_right_track_0.mux_l2_in_3_/S
+ mux_right_track_0.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_12.mux_l2_in_0_ mux_top_track_12.mux_l1_in_1_/X mux_top_track_12.mux_l1_in_0_/X
+ mux_top_track_12.mux_l2_in_0_/S mux_top_track_12.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l3_in_0_/X _059_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_17.mux_l3_in_0_ mux_left_track_17.mux_l2_in_1_/X mux_left_track_17.mux_l2_in_0_/X
+ mux_left_track_17.mux_l3_in_0_/S mux_left_track_17.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_12.mux_l1_in_1_ _031_/HI chanx_left_in[10] mux_top_track_12.mux_l1_in_1_/S
+ mux_top_track_12.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_072_ chanx_right_in[2] chanx_left_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l2_in_1_ mux_left_track_17.mux_l1_in_3_/X mux_left_track_17.mux_l1_in_2_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_055_ _055_/HI _055_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_1_/S mux_right_track_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_107_ _107_/A chany_top_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l1_in_2_ left_bottom_grid_pin_3_ chanx_right_in[17] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_038_ _038_/HI _038_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_16.mux_l2_in_0_/S mux_top_track_18.mux_l1_in_1_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_9.mux_l2_in_1_ chanx_right_in[16] chanx_right_in[6] mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_0.mux_l2_in_1_ right_bottom_grid_pin_13_ right_bottom_grid_pin_9_
+ mux_right_track_0.mux_l2_in_3_/S mux_right_track_0.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_12.mux_l1_in_0_ chanx_right_in[10] top_left_grid_pin_44_ mux_top_track_12.mux_l1_in_1_/S
+ mux_top_track_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_0_/S mux_top_track_24.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_071_ _071_/A chanx_left_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_2.mux_l1_in_3_ _035_/HI chanx_left_in[4] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l1_in_3_ _053_/HI chanx_left_in[18] mux_right_track_24.mux_l1_in_2_/S
+ mux_right_track_24.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l1_in_1_ _038_/HI chanx_left_in[18] mux_top_track_24.mux_l1_in_1_/S
+ mux_top_track_24.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_054_ _054_/HI _054_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_106_ _106_/A chany_top_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_17.mux_l1_in_1_ chanx_right_in[8] chany_top_in[17] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_037_ _037_/HI _037_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_9.mux_l2_in_0_ chany_top_in[18] mux_left_track_9.mux_l1_in_0_/X mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_3_/S mux_right_track_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S mux_top_track_2.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_5_ right_bottom_grid_pin_1_
+ mux_right_track_0.mux_l1_in_0_/S mux_right_track_0.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_1_ mux_right_track_24.mux_l1_in_3_/X mux_right_track_24.mux_l1_in_2_/X
+ mux_right_track_24.mux_l2_in_0_/S mux_right_track_24.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_1_ mux_top_track_2.mux_l1_in_3_/X mux_top_track_2.mux_l1_in_2_/X
+ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_070_ chanx_right_in[4] chanx_left_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_top_track_0.mux_l3_in_1_/S mux_top_track_0.mux_l4_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l2_in_0_/X _103_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_24.mux_l1_in_2_ chanx_left_in[9] right_bottom_grid_pin_13_ mux_right_track_24.mux_l1_in_2_/S
+ mux_right_track_24.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l1_in_2_ chanx_right_in[4] chanx_right_in[3] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_053_ _053_/HI _053_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_top_track_24.mux_l1_in_0_ chanx_right_in[18] top_left_grid_pin_42_ mux_top_track_24.mux_l1_in_1_/S
+ mux_top_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_32.mux_l3_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_18.sky130_fd_sc_hd__buf_4_0_ mux_top_track_18.mux_l2_in_0_/X _106_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_14_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_105_ _105_/A chany_top_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_036_ _036_/HI _036_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_0_ chany_top_in[10] chany_top_in[3] mux_left_track_17.mux_l1_in_0_/S
+ mux_left_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l4_in_0_/X _095_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_left_track_9.mux_l1_in_0_ chany_top_in[11] chany_top_in[4] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_0.mux_l1_in_0_ chany_top_in[13] chany_top_in[6] mux_right_track_0.mux_l1_in_0_/S
+ mux_right_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_24.mux_l2_in_0_ mux_right_track_24.mux_l1_in_1_/X mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S mux_right_track_24.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X _114_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_ mux_left_track_3.mux_l3_in_0_/S mux_left_track_3.mux_l4_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_0.mux_l2_in_0_/S mux_top_track_0.mux_l3_in_1_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_18_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_24.mux_l1_in_1_ right_bottom_grid_pin_5_ chany_top_in[18] mux_right_track_24.mux_l1_in_2_/S
+ mux_right_track_24.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l1_in_1_ top_left_grid_pin_49_ top_left_grid_pin_47_ mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_052_ _052_/HI _052_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l2_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_104_ _104_/A chany_top_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_6_ left_bottom_grid_pin_17_ left_bottom_grid_pin_15_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_6_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_035_ _035_/HI _035_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_track_0.mux_l3_in_1_/S mux_right_track_0.mux_l4_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_3.mux_l2_in_1_/S mux_left_track_3.mux_l3_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_0.mux_l1_in_0_/S mux_top_track_0.mux_l2_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.mux_l1_in_0_ chany_top_in[11] chany_top_in[4] mux_right_track_24.mux_l1_in_2_/S
+ mux_right_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l1_in_0_ top_left_grid_pin_45_ top_left_grid_pin_43_ mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_051_ _051_/HI _051_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_24.mux_l3_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l4_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_20_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_034_ _034_/HI _034_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_103_ _103_/A chany_top_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_6.mux_l2_in_1_/S mux_top_track_6.mux_l3_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l1_in_5_ left_bottom_grid_pin_13_ left_bottom_grid_pin_11_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_5_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_0.mux_l2_in_3_/S mux_right_track_0.mux_l3_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_3.mux_l1_in_0_/S mux_left_track_3.mux_l2_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ ccff_head mux_top_track_0.mux_l1_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_050_ _050_/HI _050_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_left_track_5.mux_l2_in_3_ _048_/HI mux_left_track_5.mux_l1_in_6_/X mux_left_track_5.mux_l2_in_0_/S
+ mux_left_track_5.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_9.mux_l2_in_0_/S mux_left_track_9.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_033_ _033_/HI _033_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_28_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_102_ top_left_grid_pin_43_ chany_top_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_6.mux_l1_in_3_/S mux_top_track_6.mux_l2_in_1_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l1_in_4_ left_bottom_grid_pin_9_ left_bottom_grid_pin_7_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_4_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_5.mux_l4_in_0_ mux_left_track_5.mux_l3_in_1_/X mux_left_track_5.mux_l3_in_0_/X
+ mux_left_track_5.mux_l4_in_0_/S mux_left_track_5.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_22.mux_l1_in_0_/S mux_top_track_22.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_0.mux_l1_in_0_/S mux_right_track_0.mux_l2_in_3_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l3_in_1_ mux_left_track_5.mux_l2_in_3_/X mux_left_track_5.mux_l2_in_2_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_1.mux_l4_in_0_/S mux_left_track_3.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_2_ mux_left_track_5.mux_l1_in_5_/X mux_left_track_5.mux_l1_in_4_/X
+ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l2_in_2_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_101_ chanx_left_in[19] chany_top_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_032_ _032_/HI _032_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_3_ left_bottom_grid_pin_5_ left_bottom_grid_pin_3_ mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_4.mux_l3_in_0_/S mux_top_track_6.mux_l1_in_3_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_20.mux_l2_in_0_/S mux_top_track_22.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l3_in_0_/X _067_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_38.mux_l2_in_0_/S mux_right_track_0.mux_l1_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l3_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_100_ chanx_left_in[15] chany_top_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_031_ _031_/HI _031_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_5.mux_l4_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_25.mux_l1_in_3_ _045_/HI left_bottom_grid_pin_13_ mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.mux_l1_in_2_ left_bottom_grid_pin_1_ chanx_right_in[14] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_18.mux_l2_in_0_ mux_top_track_18.mux_l1_in_1_/X mux_top_track_18.mux_l1_in_0_/X
+ mux_top_track_18.mux_l2_in_0_/S mux_top_track_18.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_33.mux_l2_in_0_/S ccff_tail
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_20.mux_l2_in_0_ mux_top_track_20.mux_l1_in_1_/X mux_top_track_20.mux_l1_in_0_/X
+ mux_top_track_20.mux_l2_in_0_/S mux_top_track_20.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_18.mux_l1_in_1_ _034_/HI chanx_left_in[14] mux_top_track_18.mux_l1_in_1_/S
+ mux_top_track_18.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_20.mux_l1_in_1_ _036_/HI chanx_left_in[16] mux_top_track_20.mux_l1_in_1_/S
+ mux_top_track_20.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l3_in_0_ mux_left_track_25.mux_l2_in_1_/X mux_left_track_25.mux_l2_in_0_/X
+ mux_left_track_25.mux_l3_in_0_/S mux_left_track_25.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_24.mux_l1_in_2_/S
+ mux_right_track_24.mux_l2_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l2_in_1_ mux_left_track_25.mux_l1_in_3_/X mux_left_track_25.mux_l1_in_2_/X
+ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_030_ _030_/HI _030_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_5.mux_l1_in_1_ chanx_right_in[5] chany_top_in[19] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_2_ left_bottom_grid_pin_5_ chanx_right_in[18] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_20.sky130_fd_sc_hd__buf_4_0_ mux_top_track_20.mux_l2_in_0_/X _105_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_31_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_33.mux_l1_in_1_/S mux_left_track_33.mux_l2_in_0_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_18.mux_l1_in_0_ chanx_right_in[14] top_left_grid_pin_47_ mux_top_track_18.mux_l1_in_1_/S
+ mux_top_track_18.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_14.sky130_fd_sc_hd__buf_4_0_ mux_top_track_14.mux_l2_in_0_/X _108_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_top_track_20.mux_l1_in_0_ chanx_right_in[16] top_left_grid_pin_48_ mux_top_track_20.mux_l1_in_1_/S
+ mux_top_track_20.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_16.mux_l3_in_0_/S
+ mux_right_track_24.mux_l1_in_2_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_0_ chany_top_in[12] chany_top_in[5] mux_left_track_5.mux_l1_in_0_/S
+ mux_left_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l1_in_1_ chanx_right_in[9] chany_top_in[16] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_089_ chanx_left_in[5] chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S mux_top_track_8.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_25.mux_l3_in_0_/S mux_left_track_33.mux_l1_in_1_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_right_track_32.mux_l3_in_0_ mux_right_track_32.mux_l2_in_1_/X mux_right_track_32.mux_l2_in_0_/X
+ mux_right_track_32.mux_l3_in_0_/S mux_right_track_32.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_8.mux_l2_in_1_ _042_/HI chanx_left_in[8] mux_top_track_8.mux_l2_in_1_/S
+ mux_top_track_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_7_0_prog_clk clkbuf_3_6_0_prog_clk/A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_32.mux_l2_in_1_ _054_/HI mux_right_track_32.mux_l1_in_2_/X mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_32.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_32.mux_l1_in_2_ chanx_left_in[10] right_bottom_grid_pin_15_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_088_ chanx_left_in[6] chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l1_in_0_ chany_top_in[9] chany_top_in[2] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_14.mux_l1_in_0_/S mux_top_track_14.mux_l2_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_8.mux_l2_in_0_ chanx_right_in[15] mux_top_track_8.mux_l1_in_0_/X mux_top_track_8.mux_l2_in_1_/S
+ mux_top_track_8.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l2_in_0_ mux_right_track_32.mux_l1_in_1_/X mux_right_track_32.mux_l1_in_0_/X
+ mux_right_track_32.mux_l2_in_0_/S mux_right_track_32.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_26_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l3_in_0_/X _111_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l1_in_1_ right_bottom_grid_pin_7_ chany_top_in[19] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_087_ _087_/A chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_12.mux_l2_in_0_/S mux_top_track_14.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X _083_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_1.mux_l2_in_3_ _043_/HI left_bottom_grid_pin_17_ mux_left_track_1.mux_l2_in_3_/S
+ mux_left_track_1.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_16.mux_l2_in_1_/S
+ mux_right_track_16.mux_l3_in_0_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_0_ chanx_right_in[8] top_left_grid_pin_42_ mux_top_track_8.mux_l1_in_0_/S
+ mux_top_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_32.mux_l1_in_0_ chany_top_in[12] chany_top_in[5] mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l4_in_0_ mux_left_track_1.mux_l3_in_1_/X mux_left_track_1.mux_l3_in_0_/X
+ mux_left_track_1.mux_l4_in_0_/S mux_left_track_1.mux_l4_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ chanx_left_in[8] chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_25.mux_l2_in_0_/S mux_left_track_25.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l4_in_0_/X _074_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmux_left_track_1.mux_l3_in_1_ mux_left_track_1.mux_l2_in_3_/X mux_left_track_1.mux_l2_in_2_/X
+ mux_left_track_1.mux_l3_in_1_/S mux_left_track_1.mux_l3_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_069_ chanx_right_in[5] chanx_left_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_1.mux_l2_in_2_ left_bottom_grid_pin_13_ left_bottom_grid_pin_9_ mux_left_track_1.mux_l2_in_3_/S
+ mux_left_track_1.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_16.mux_l1_in_3_/S
+ mux_right_track_16.mux_l2_in_1_/S clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_prog_clk clkbuf_3_6_0_prog_clk/A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_2.mux_l2_in_3_ _052_/HI chanx_left_in[13] mux_right_track_2.mux_l2_in_2_/S
+ mux_right_track_2.mux_l2_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_085_ chanx_left_in[9] chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_25.mux_l1_in_0_/S mux_left_track_25.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_1_/S mux_left_track_1.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_068_ chanx_right_in[6] chanx_left_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_2.mux_l4_in_0_ mux_right_track_2.mux_l3_in_1_/X mux_right_track_2.mux_l3_in_0_/X
+ mux_right_track_2.mux_l4_in_0_/S mux_right_track_2.mux_l4_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_1.mux_l2_in_1_ left_bottom_grid_pin_5_ mux_left_track_1.mux_l1_in_2_/X
+ mux_left_track_1.mux_l2_in_3_/S mux_left_track_1.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l3_in_1_ mux_right_track_2.mux_l2_in_3_/X mux_right_track_2.mux_l2_in_2_/X
+ mux_right_track_2.mux_l3_in_1_/S mux_right_track_2.mux_l3_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_ mux_right_track_8.mux_l4_in_0_/S mux_right_track_16.mux_l1_in_3_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_left_track_1.mux_l1_in_2_ left_bottom_grid_pin_1_ chanx_right_in[12] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_2_ chanx_left_in[4] right_bottom_grid_pin_15_ mux_right_track_2.mux_l2_in_2_/S
+ mux_right_track_2.mux_l2_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_14.mux_l2_in_0_ mux_top_track_14.mux_l1_in_1_/X mux_top_track_14.mux_l1_in_0_/X
+ mux_top_track_14.mux_l2_in_0_/S mux_top_track_14.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_084_ chanx_left_in[10] chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_17.mux_l3_in_0_/S mux_left_track_25.mux_l1_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_14.mux_l1_in_1_ _032_/HI chanx_left_in[12] mux_top_track_14.mux_l1_in_0_/S
+ mux_top_track_14.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_38.mux_l1_in_0_/S mux_top_track_38.mux_l2_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_067_ _067_/A chanx_left_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_3_/S mux_left_track_1.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_1_/S mux_right_track_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_0 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_1.mux_l1_in_1_ chanx_right_in[2] chany_top_in[14] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_1_ right_bottom_grid_pin_11_ right_bottom_grid_pin_7_
+ mux_right_track_2.mux_l2_in_2_/S mux_right_track_2.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_10.sky130_fd_sc_hd__buf_4_0_ mux_top_track_10.mux_l3_in_0_/X _110_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_083_ _083_/A chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l4_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_14.mux_l1_in_0_ chanx_right_in[12] top_left_grid_pin_45_ mux_top_track_14.mux_l1_in_0_/S
+ mux_top_track_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_2.mux_l2_in_0_/S mux_top_track_2.mux_l3_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_24.mux_l2_in_0_/S mux_top_track_38.mux_l1_in_0_/S
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
X_066_ chanx_right_in[8] chanx_left_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_3_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_3_6_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_049_ _049_/HI _049_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_4.mux_l1_in_3_ _040_/HI chanx_left_in[5] mux_top_track_4.mux_l1_in_3_/S
+ mux_top_track_4.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l3_in_0_ mux_left_track_33.mux_l2_in_1_/X mux_left_track_33.mux_l2_in_0_/X
+ ccff_tail mux_left_track_33.mux_l3_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l1_in_0_ chany_top_in[7] chany_top_in[0] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_2_/S mux_right_track_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l2_in_1_ _047_/HI mux_left_track_33.mux_l1_in_2_/X mux_left_track_33.mux_l2_in_0_/S
+ mux_left_track_33.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_track_2.mux_l3_in_1_/S mux_right_track_2.mux_l4_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_082_ chanx_left_in[12] chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_5.mux_l2_in_0_/S mux_left_track_5.mux_l3_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_5_0_prog_clk clkbuf_2_2_0_prog_clk/X clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_10_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_2.mux_l1_in_1_ right_bottom_grid_pin_3_ chany_top_in[14] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_2.mux_l1_in_1_/S mux_top_track_2.mux_l2_in_0_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_1_ mux_top_track_4.mux_l1_in_3_/X mux_top_track_4.mux_l1_in_2_/X
+ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l2_in_1_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l1_in_2_ left_bottom_grid_pin_15_ left_bottom_grid_pin_7_ mux_left_track_33.mux_l1_in_1_/S
+ mux_left_track_33.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_065_ chanx_right_in[9] chanx_left_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_4.mux_l1_in_2_ chanx_right_in[7] chanx_right_in[5] mux_top_track_4.mux_l1_in_3_/S
+ mux_top_track_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ mux_top_track_8.mux_l2_in_1_/S mux_top_track_8.mux_l3_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_048_ _048_/HI _048_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_38.mux_l2_in_0_ _039_/HI mux_top_track_38.mux_l1_in_0_/X mux_top_track_38.mux_l2_in_0_/S
+ mux_top_track_38.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_2 top_left_grid_pin_49_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l1_in_1_/X mux_left_track_33.mux_l1_in_0_/X
+ mux_left_track_33.mux_l2_in_0_/S mux_left_track_33.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_2.mux_l2_in_2_/S mux_right_track_2.mux_l3_in_1_/S
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l3_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_081_ chanx_left_in[13] chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l4_in_0_/X _094_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_5.mux_l1_in_0_/S mux_left_track_5.mux_l2_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l1_in_0_ chany_top_in[7] chany_top_in[0] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l1_in_1_ chanx_right_in[10] chany_top_in[15] mux_left_track_33.mux_l1_in_1_/S
+ mux_left_track_33.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_0.mux_l4_in_0_/S mux_top_track_2.mux_l1_in_1_/S
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_064_ chanx_right_in[10] chanx_left_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X _113_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l4_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l1_in_1_ top_left_grid_pin_48_ top_left_grid_pin_46_ mux_top_track_4.mux_l1_in_3_/S
+ mux_top_track_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_047_ _047_/HI _047_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_8.mux_l1_in_0_/S mux_top_track_8.mux_l2_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_29_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ mux_top_track_24.mux_l1_in_1_/S mux_top_track_24.mux_l2_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_2_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_16_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_ mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l2_in_2_/S
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_38.mux_l1_in_0_ chanx_left_in[1] chanx_right_in[0] mux_top_track_38.mux_l1_in_0_/S
+ mux_top_track_38.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ mux_left_track_17.mux_l1_in_0_/S mux_left_track_17.mux_l2_in_0_/S
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_080_ chanx_left_in[14] chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_27_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ mux_left_track_3.mux_l4_in_0_/S mux_left_track_5.mux_l1_in_0_/S
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_33.mux_l1_in_0_ chany_top_in[8] chany_top_in[1] mux_left_track_33.mux_l1_in_1_/S
+ mux_left_track_33.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_063_ _063_/A chanx_left_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_ mux_right_track_8.mux_l2_in_0_/S mux_right_track_8.mux_l3_in_0_/S
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l1_in_0_ top_left_grid_pin_44_ top_left_grid_pin_42_ mux_top_track_4.mux_l1_in_3_/S
+ mux_top_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_115_ _115_/A chany_top_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_046_ _046_/HI _046_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_6.mux_l3_in_0_/S mux_top_track_8.mux_l1_in_0_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_prog_clk clkbuf_2_3_0_prog_clk/A clkbuf_2_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_029_ _029_/HI _029_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ mux_top_track_22.mux_l2_in_0_/S mux_top_track_24.mux_l1_in_1_/S
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxtp_1
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

