VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_right_right
  CLASS BLOCK ;
  FOREIGN grid_io_right_right ;
  ORIGIN 0.000 0.000 ;
  SIZE 45.000 BY 76.800 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END IO_ISOL_N
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 2.400 ;
    END
  END ccff_tail
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 42.600 42.200 45.000 42.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 2.400 76.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
  PIN left_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END left_width_0_height_0__pin_0_
  PIN left_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END left_width_0_height_0__pin_1_lower
  PIN left_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 2.400 42.800 ;
    END
  END left_width_0_height_0__pin_1_upper
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 2.400 ;
    END
  END prog_clk
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.380 10.640 11.980 73.680 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 16.040 10.640 17.640 73.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 39.100 73.525 ;
      LAYER met1 ;
        RECT 5.520 10.640 39.490 73.680 ;
      LAYER met2 ;
        RECT 5.620 2.680 39.460 76.685 ;
        RECT 6.170 2.400 16.370 2.680 ;
        RECT 17.210 2.400 27.870 2.680 ;
        RECT 28.710 2.400 38.910 2.680 ;
      LAYER met3 ;
        RECT 2.800 75.800 42.600 76.665 ;
        RECT 2.400 60.200 42.600 75.800 ;
        RECT 2.800 58.800 42.600 60.200 ;
        RECT 2.400 43.200 42.600 58.800 ;
        RECT 2.800 41.800 42.200 43.200 ;
        RECT 2.400 26.200 42.600 41.800 ;
        RECT 2.800 24.800 42.600 26.200 ;
        RECT 2.400 9.200 42.600 24.800 ;
        RECT 2.800 8.335 42.600 9.200 ;
      LAYER met4 ;
        RECT 21.700 10.640 34.620 73.680 ;
  END
END grid_io_right_right
END LIBRARY

