magic
tech sky130A
magscale 1 2
timestamp 1606426228
<< locali >>
rect 10149 10523 10183 10761
<< viali >>
rect 4261 15657 4295 15691
rect 4077 15521 4111 15555
rect 4629 15521 4663 15555
rect 5365 15521 5399 15555
rect 4813 15385 4847 15419
rect 5549 15385 5583 15419
rect 7297 15113 7331 15147
rect 9413 15113 9447 15147
rect 7113 14909 7147 14943
rect 9229 14909 9263 14943
rect 15209 14025 15243 14059
rect 5641 13957 5675 13991
rect 4261 13821 4295 13855
rect 4517 13821 4551 13855
rect 15025 13821 15059 13855
rect 4813 13481 4847 13515
rect 2697 13345 2731 13379
rect 3065 13345 3099 13379
rect 4997 13345 5031 13379
rect 3157 13141 3191 13175
rect 7573 12869 7607 12903
rect 8125 12801 8159 12835
rect 8033 12733 8067 12767
rect 7941 12665 7975 12699
rect 7297 12393 7331 12427
rect 8217 12325 8251 12359
rect 6009 12257 6043 12291
rect 8309 12189 8343 12223
rect 8401 12189 8435 12223
rect 7849 12121 7883 12155
rect 9137 11849 9171 11883
rect 7481 11713 7515 11747
rect 7757 11645 7791 11679
rect 7205 11577 7239 11611
rect 8002 11577 8036 11611
rect 6837 11509 6871 11543
rect 7297 11509 7331 11543
rect 6745 11305 6779 11339
rect 10149 11305 10183 11339
rect 4169 11237 4203 11271
rect 4261 11237 4295 11271
rect 6653 11237 6687 11271
rect 7297 11169 7331 11203
rect 7564 11169 7598 11203
rect 10057 11169 10091 11203
rect 5181 11101 5215 11135
rect 6929 11101 6963 11135
rect 10241 11101 10275 11135
rect 6285 11033 6319 11067
rect 8677 10965 8711 10999
rect 9689 10965 9723 10999
rect 2927 10761 2961 10795
rect 7297 10761 7331 10795
rect 10149 10761 10183 10795
rect 8953 10693 8987 10727
rect 2421 10625 2455 10659
rect 7573 10625 7607 10659
rect 9781 10625 9815 10659
rect 2840 10557 2874 10591
rect 7481 10557 7515 10591
rect 9597 10557 9631 10591
rect 10793 10625 10827 10659
rect 10609 10557 10643 10591
rect 1501 10489 1535 10523
rect 1593 10489 1627 10523
rect 7840 10489 7874 10523
rect 10149 10489 10183 10523
rect 9229 10421 9263 10455
rect 9689 10421 9723 10455
rect 10241 10421 10275 10455
rect 10701 10421 10735 10455
rect 6561 10217 6595 10251
rect 9781 10217 9815 10251
rect 7472 10149 7506 10183
rect 6653 10081 6687 10115
rect 7205 10081 7239 10115
rect 6837 10013 6871 10047
rect 6193 9877 6227 9911
rect 8585 9877 8619 9911
rect 7205 9605 7239 9639
rect 7757 9537 7791 9571
rect 8677 9537 8711 9571
rect 8769 9537 8803 9571
rect 7665 9469 7699 9503
rect 7573 9401 7607 9435
rect 8217 9333 8251 9367
rect 8585 9333 8619 9367
rect 12357 8993 12391 9027
rect 12633 8925 12667 8959
rect 3249 7293 3283 7327
rect 3525 7225 3559 7259
rect 8125 5865 8159 5899
rect 9137 5865 9171 5899
rect 4353 5729 4387 5763
rect 5181 5729 5215 5763
rect 6837 5729 6871 5763
rect 7389 5729 7423 5763
rect 7941 5729 7975 5763
rect 8953 5729 8987 5763
rect 9689 5729 9723 5763
rect 10241 5729 10275 5763
rect 11529 5729 11563 5763
rect 9873 5593 9907 5627
rect 11713 5593 11747 5627
rect 4537 5525 4571 5559
rect 5365 5525 5399 5559
rect 7021 5525 7055 5559
rect 7573 5525 7607 5559
rect 10425 5525 10459 5559
rect 8493 5321 8527 5355
rect 10333 5321 10367 5355
rect 11437 5321 11471 5355
rect 11989 5321 12023 5355
rect 9781 5253 9815 5287
rect 3709 5117 3743 5151
rect 4813 5117 4847 5151
rect 5641 5117 5675 5151
rect 6193 5117 6227 5151
rect 6837 5117 6871 5151
rect 7389 5117 7423 5151
rect 8309 5117 8343 5151
rect 9045 5117 9079 5151
rect 9597 5117 9631 5151
rect 10149 5117 10183 5151
rect 10701 5117 10735 5151
rect 11253 5117 11287 5151
rect 11805 5117 11839 5151
rect 12449 5117 12483 5151
rect 13001 5117 13035 5151
rect 3893 4981 3927 5015
rect 4997 4981 5031 5015
rect 5825 4981 5859 5015
rect 6377 4981 6411 5015
rect 7021 4981 7055 5015
rect 7573 4981 7607 5015
rect 9229 4981 9263 5015
rect 10885 4981 10919 5015
rect 12633 4981 12667 5015
rect 13185 4981 13219 5015
rect 5089 4777 5123 4811
rect 5917 4777 5951 4811
rect 9229 4777 9263 4811
rect 9873 4777 9907 4811
rect 4905 4641 4939 4675
rect 5733 4641 5767 4675
rect 7021 4641 7055 4675
rect 7849 4641 7883 4675
rect 8401 4641 8435 4675
rect 9045 4641 9079 4675
rect 9689 4641 9723 4675
rect 10701 4641 10735 4675
rect 11897 4641 11931 4675
rect 7205 4437 7239 4471
rect 8033 4437 8067 4471
rect 8585 4437 8619 4471
rect 10885 4437 10919 4471
rect 12081 4437 12115 4471
rect 7757 4029 7791 4063
rect 9873 4029 9907 4063
rect 7941 3893 7975 3927
rect 10057 3893 10091 3927
<< metal1 >>
rect 3050 17892 3056 17944
rect 3108 17932 3114 17944
rect 4890 17932 4896 17944
rect 3108 17904 4896 17932
rect 3108 17892 3114 17904
rect 4890 17892 4896 17904
rect 4948 17892 4954 17944
rect 1104 17434 15824 17456
rect 1104 17382 3447 17434
rect 3499 17382 3511 17434
rect 3563 17382 3575 17434
rect 3627 17382 3639 17434
rect 3691 17382 8378 17434
rect 8430 17382 8442 17434
rect 8494 17382 8506 17434
rect 8558 17382 8570 17434
rect 8622 17382 13308 17434
rect 13360 17382 13372 17434
rect 13424 17382 13436 17434
rect 13488 17382 13500 17434
rect 13552 17382 15824 17434
rect 1104 17360 15824 17382
rect 1104 16890 15824 16912
rect 1104 16838 5912 16890
rect 5964 16838 5976 16890
rect 6028 16838 6040 16890
rect 6092 16838 6104 16890
rect 6156 16838 10843 16890
rect 10895 16838 10907 16890
rect 10959 16838 10971 16890
rect 11023 16838 11035 16890
rect 11087 16838 15824 16890
rect 1104 16816 15824 16838
rect 6270 16532 6276 16584
rect 6328 16572 6334 16584
rect 10410 16572 10416 16584
rect 6328 16544 10416 16572
rect 6328 16532 6334 16544
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 5534 16464 5540 16516
rect 5592 16504 5598 16516
rect 9950 16504 9956 16516
rect 5592 16476 9956 16504
rect 5592 16464 5598 16476
rect 9950 16464 9956 16476
rect 10008 16464 10014 16516
rect 6362 16396 6368 16448
rect 6420 16436 6426 16448
rect 10318 16436 10324 16448
rect 6420 16408 10324 16436
rect 6420 16396 6426 16408
rect 10318 16396 10324 16408
rect 10376 16396 10382 16448
rect 1104 16346 15824 16368
rect 1104 16294 3447 16346
rect 3499 16294 3511 16346
rect 3563 16294 3575 16346
rect 3627 16294 3639 16346
rect 3691 16294 8378 16346
rect 8430 16294 8442 16346
rect 8494 16294 8506 16346
rect 8558 16294 8570 16346
rect 8622 16294 13308 16346
rect 13360 16294 13372 16346
rect 13424 16294 13436 16346
rect 13488 16294 13500 16346
rect 13552 16294 15824 16346
rect 1104 16272 15824 16294
rect 7650 16192 7656 16244
rect 7708 16232 7714 16244
rect 10502 16232 10508 16244
rect 7708 16204 10508 16232
rect 7708 16192 7714 16204
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 6822 16124 6828 16176
rect 6880 16164 6886 16176
rect 9766 16164 9772 16176
rect 6880 16136 9772 16164
rect 6880 16124 6886 16136
rect 9766 16124 9772 16136
rect 9824 16124 9830 16176
rect 7282 16056 7288 16108
rect 7340 16096 7346 16108
rect 8846 16096 8852 16108
rect 7340 16068 8852 16096
rect 7340 16056 7346 16068
rect 8846 16056 8852 16068
rect 8904 16056 8910 16108
rect 10502 16056 10508 16108
rect 10560 16096 10566 16108
rect 11330 16096 11336 16108
rect 10560 16068 11336 16096
rect 10560 16056 10566 16068
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 8662 15988 8668 16040
rect 8720 16028 8726 16040
rect 9582 16028 9588 16040
rect 8720 16000 9588 16028
rect 8720 15988 8726 16000
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 10686 15988 10692 16040
rect 10744 16028 10750 16040
rect 11790 16028 11796 16040
rect 10744 16000 11796 16028
rect 10744 15988 10750 16000
rect 11790 15988 11796 16000
rect 11848 15988 11854 16040
rect 13078 15988 13084 16040
rect 13136 16028 13142 16040
rect 16298 16028 16304 16040
rect 13136 16000 16304 16028
rect 13136 15988 13142 16000
rect 16298 15988 16304 16000
rect 16356 15988 16362 16040
rect 8202 15920 8208 15972
rect 8260 15960 8266 15972
rect 9674 15960 9680 15972
rect 8260 15932 9680 15960
rect 8260 15920 8266 15932
rect 9674 15920 9680 15932
rect 9732 15920 9738 15972
rect 13814 15960 13820 15972
rect 9784 15932 13820 15960
rect 1854 15852 1860 15904
rect 1912 15892 1918 15904
rect 2682 15892 2688 15904
rect 1912 15864 2688 15892
rect 1912 15852 1918 15864
rect 2682 15852 2688 15864
rect 2740 15852 2746 15904
rect 4338 15852 4344 15904
rect 4396 15892 4402 15904
rect 5350 15892 5356 15904
rect 4396 15864 5356 15892
rect 4396 15852 4402 15864
rect 5350 15852 5356 15864
rect 5408 15852 5414 15904
rect 9306 15852 9312 15904
rect 9364 15892 9370 15904
rect 9784 15892 9812 15932
rect 13814 15920 13820 15932
rect 13872 15920 13878 15972
rect 9364 15864 9812 15892
rect 9364 15852 9370 15864
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 13170 15892 13176 15904
rect 9916 15864 13176 15892
rect 9916 15852 9922 15864
rect 13170 15852 13176 15864
rect 13228 15852 13234 15904
rect 1104 15802 15824 15824
rect 1104 15750 5912 15802
rect 5964 15750 5976 15802
rect 6028 15750 6040 15802
rect 6092 15750 6104 15802
rect 6156 15750 10843 15802
rect 10895 15750 10907 15802
rect 10959 15750 10971 15802
rect 11023 15750 11035 15802
rect 11087 15750 15824 15802
rect 1104 15728 15824 15750
rect 566 15648 572 15700
rect 624 15688 630 15700
rect 4249 15691 4307 15697
rect 4249 15688 4261 15691
rect 624 15660 4261 15688
rect 624 15648 630 15660
rect 4249 15657 4261 15660
rect 4295 15657 4307 15691
rect 7098 15688 7104 15700
rect 4249 15651 4307 15657
rect 4540 15660 7104 15688
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4540 15552 4568 15660
rect 7098 15648 7104 15660
rect 7156 15648 7162 15700
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 12986 15688 12992 15700
rect 9548 15660 12992 15688
rect 9548 15648 9554 15660
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 6270 15620 6276 15632
rect 4632 15592 6276 15620
rect 4632 15561 4660 15592
rect 6270 15580 6276 15592
rect 6328 15580 6334 15632
rect 9214 15580 9220 15632
rect 9272 15620 9278 15632
rect 9858 15620 9864 15632
rect 9272 15592 9864 15620
rect 9272 15580 9278 15592
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 4111 15524 4568 15552
rect 4617 15555 4675 15561
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 4617 15521 4629 15555
rect 4663 15521 4675 15555
rect 4617 15515 4675 15521
rect 5353 15555 5411 15561
rect 5353 15521 5365 15555
rect 5399 15552 5411 15555
rect 7834 15552 7840 15564
rect 5399 15524 7840 15552
rect 5399 15521 5411 15524
rect 5353 15515 5411 15521
rect 7834 15512 7840 15524
rect 7892 15512 7898 15564
rect 8018 15512 8024 15564
rect 8076 15552 8082 15564
rect 10594 15552 10600 15564
rect 8076 15524 10600 15552
rect 8076 15512 8082 15524
rect 10594 15512 10600 15524
rect 10652 15512 10658 15564
rect 15102 15552 15108 15564
rect 13740 15524 15108 15552
rect 2222 15444 2228 15496
rect 2280 15484 2286 15496
rect 2280 15456 5580 15484
rect 2280 15444 2286 15456
rect 1394 15376 1400 15428
rect 1452 15416 1458 15428
rect 5552 15425 5580 15456
rect 7742 15444 7748 15496
rect 7800 15484 7806 15496
rect 11422 15484 11428 15496
rect 7800 15456 11428 15484
rect 7800 15444 7806 15456
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 11974 15444 11980 15496
rect 12032 15484 12038 15496
rect 13740 15484 13768 15524
rect 15102 15512 15108 15524
rect 15160 15512 15166 15564
rect 12032 15456 13768 15484
rect 12032 15444 12038 15456
rect 14458 15444 14464 15496
rect 14516 15484 14522 15496
rect 15930 15484 15936 15496
rect 14516 15456 15936 15484
rect 14516 15444 14522 15456
rect 15930 15444 15936 15456
rect 15988 15444 15994 15496
rect 4801 15419 4859 15425
rect 4801 15416 4813 15419
rect 1452 15388 4813 15416
rect 1452 15376 1458 15388
rect 4801 15385 4813 15388
rect 4847 15385 4859 15419
rect 4801 15379 4859 15385
rect 5537 15419 5595 15425
rect 5537 15385 5549 15419
rect 5583 15385 5595 15419
rect 5537 15379 5595 15385
rect 8110 15376 8116 15428
rect 8168 15416 8174 15428
rect 12158 15416 12164 15428
rect 8168 15388 12164 15416
rect 8168 15376 8174 15388
rect 12158 15376 12164 15388
rect 12216 15376 12222 15428
rect 12986 15376 12992 15428
rect 13044 15416 13050 15428
rect 16758 15416 16764 15428
rect 13044 15388 16764 15416
rect 13044 15376 13050 15388
rect 16758 15376 16764 15388
rect 16816 15376 16822 15428
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 6822 15348 6828 15360
rect 4764 15320 6828 15348
rect 4764 15308 4770 15320
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 7190 15308 7196 15360
rect 7248 15348 7254 15360
rect 9398 15348 9404 15360
rect 7248 15320 9404 15348
rect 7248 15308 7254 15320
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 1104 15258 15824 15280
rect 1104 15206 3447 15258
rect 3499 15206 3511 15258
rect 3563 15206 3575 15258
rect 3627 15206 3639 15258
rect 3691 15206 8378 15258
rect 8430 15206 8442 15258
rect 8494 15206 8506 15258
rect 8558 15206 8570 15258
rect 8622 15206 13308 15258
rect 13360 15206 13372 15258
rect 13424 15206 13436 15258
rect 13488 15206 13500 15258
rect 13552 15206 15824 15258
rect 1104 15184 15824 15206
rect 6822 15104 6828 15156
rect 6880 15144 6886 15156
rect 7285 15147 7343 15153
rect 7285 15144 7297 15147
rect 6880 15116 7297 15144
rect 6880 15104 6886 15116
rect 7285 15113 7297 15116
rect 7331 15113 7343 15147
rect 9398 15144 9404 15156
rect 9359 15116 9404 15144
rect 7285 15107 7343 15113
rect 9398 15104 9404 15116
rect 9456 15104 9462 15156
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14909 7159 14943
rect 7101 14903 7159 14909
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14940 9275 14943
rect 10594 14940 10600 14952
rect 9263 14912 10600 14940
rect 9263 14909 9275 14912
rect 9217 14903 9275 14909
rect 7116 14872 7144 14903
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 9398 14872 9404 14884
rect 7116 14844 9404 14872
rect 9398 14832 9404 14844
rect 9456 14832 9462 14884
rect 1104 14714 15824 14736
rect 1104 14662 5912 14714
rect 5964 14662 5976 14714
rect 6028 14662 6040 14714
rect 6092 14662 6104 14714
rect 6156 14662 10843 14714
rect 10895 14662 10907 14714
rect 10959 14662 10971 14714
rect 11023 14662 11035 14714
rect 11087 14662 15824 14714
rect 1104 14640 15824 14662
rect 1104 14170 15824 14192
rect 1104 14118 3447 14170
rect 3499 14118 3511 14170
rect 3563 14118 3575 14170
rect 3627 14118 3639 14170
rect 3691 14118 8378 14170
rect 8430 14118 8442 14170
rect 8494 14118 8506 14170
rect 8558 14118 8570 14170
rect 8622 14118 13308 14170
rect 13360 14118 13372 14170
rect 13424 14118 13436 14170
rect 13488 14118 13500 14170
rect 13552 14118 15824 14170
rect 1104 14096 15824 14118
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 15197 14059 15255 14065
rect 15197 14056 15209 14059
rect 13780 14028 15209 14056
rect 13780 14016 13786 14028
rect 15197 14025 15209 14028
rect 15243 14025 15255 14059
rect 15197 14019 15255 14025
rect 5629 13991 5687 13997
rect 5629 13957 5641 13991
rect 5675 13988 5687 13991
rect 8110 13988 8116 14000
rect 5675 13960 8116 13988
rect 5675 13957 5687 13960
rect 5629 13951 5687 13957
rect 8110 13948 8116 13960
rect 8168 13948 8174 14000
rect 3970 13880 3976 13932
rect 4028 13920 4034 13932
rect 4028 13892 4384 13920
rect 4028 13880 4034 13892
rect 4246 13852 4252 13864
rect 4207 13824 4252 13852
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 4356 13852 4384 13892
rect 4505 13855 4563 13861
rect 4505 13852 4517 13855
rect 4356 13824 4517 13852
rect 4505 13821 4517 13824
rect 4551 13821 4563 13855
rect 4505 13815 4563 13821
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 15013 13855 15071 13861
rect 15013 13852 15025 13855
rect 13688 13824 15025 13852
rect 13688 13812 13694 13824
rect 15013 13821 15025 13824
rect 15059 13821 15071 13855
rect 15013 13815 15071 13821
rect 1104 13626 15824 13648
rect 1104 13574 5912 13626
rect 5964 13574 5976 13626
rect 6028 13574 6040 13626
rect 6092 13574 6104 13626
rect 6156 13574 10843 13626
rect 10895 13574 10907 13626
rect 10959 13574 10971 13626
rect 11023 13574 11035 13626
rect 11087 13574 15824 13626
rect 1104 13552 15824 13574
rect 4246 13472 4252 13524
rect 4304 13512 4310 13524
rect 4801 13515 4859 13521
rect 4801 13512 4813 13515
rect 4304 13484 4813 13512
rect 4304 13472 4310 13484
rect 4801 13481 4813 13484
rect 4847 13481 4859 13515
rect 4801 13475 4859 13481
rect 198 13336 204 13388
rect 256 13376 262 13388
rect 2685 13379 2743 13385
rect 2685 13376 2697 13379
rect 256 13348 2697 13376
rect 256 13336 262 13348
rect 2685 13345 2697 13348
rect 2731 13345 2743 13379
rect 2685 13339 2743 13345
rect 3053 13379 3111 13385
rect 3053 13345 3065 13379
rect 3099 13345 3111 13379
rect 4982 13376 4988 13388
rect 4943 13348 4988 13376
rect 3053 13339 3111 13345
rect 3068 13308 3096 13339
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 9122 13308 9128 13320
rect 3068 13280 9128 13308
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 2866 13132 2872 13184
rect 2924 13172 2930 13184
rect 3145 13175 3203 13181
rect 3145 13172 3157 13175
rect 2924 13144 3157 13172
rect 2924 13132 2930 13144
rect 3145 13141 3157 13144
rect 3191 13141 3203 13175
rect 3145 13135 3203 13141
rect 1104 13082 15824 13104
rect 1104 13030 3447 13082
rect 3499 13030 3511 13082
rect 3563 13030 3575 13082
rect 3627 13030 3639 13082
rect 3691 13030 8378 13082
rect 8430 13030 8442 13082
rect 8494 13030 8506 13082
rect 8558 13030 8570 13082
rect 8622 13030 13308 13082
rect 13360 13030 13372 13082
rect 13424 13030 13436 13082
rect 13488 13030 13500 13082
rect 13552 13030 15824 13082
rect 1104 13008 15824 13030
rect 7561 12903 7619 12909
rect 7561 12869 7573 12903
rect 7607 12900 7619 12903
rect 8662 12900 8668 12912
rect 7607 12872 8668 12900
rect 7607 12869 7619 12872
rect 7561 12863 7619 12869
rect 8662 12860 8668 12872
rect 8720 12860 8726 12912
rect 8110 12832 8116 12844
rect 8071 12804 8116 12832
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 8021 12767 8079 12773
rect 8021 12764 8033 12767
rect 7892 12736 8033 12764
rect 7892 12724 7898 12736
rect 8021 12733 8033 12736
rect 8067 12733 8079 12767
rect 8021 12727 8079 12733
rect 7650 12656 7656 12708
rect 7708 12696 7714 12708
rect 7929 12699 7987 12705
rect 7929 12696 7941 12699
rect 7708 12668 7941 12696
rect 7708 12656 7714 12668
rect 7929 12665 7941 12668
rect 7975 12665 7987 12699
rect 7929 12659 7987 12665
rect 9122 12588 9128 12640
rect 9180 12628 9186 12640
rect 13446 12628 13452 12640
rect 9180 12600 13452 12628
rect 9180 12588 9186 12600
rect 13446 12588 13452 12600
rect 13504 12588 13510 12640
rect 1104 12538 15824 12560
rect 1104 12486 5912 12538
rect 5964 12486 5976 12538
rect 6028 12486 6040 12538
rect 6092 12486 6104 12538
rect 6156 12486 10843 12538
rect 10895 12486 10907 12538
rect 10959 12486 10971 12538
rect 11023 12486 11035 12538
rect 11087 12486 15824 12538
rect 1104 12464 15824 12486
rect 4982 12384 4988 12436
rect 5040 12424 5046 12436
rect 7285 12427 7343 12433
rect 7285 12424 7297 12427
rect 5040 12396 7297 12424
rect 5040 12384 5046 12396
rect 7285 12393 7297 12396
rect 7331 12424 7343 12427
rect 7374 12424 7380 12436
rect 7331 12396 7380 12424
rect 7331 12393 7343 12396
rect 7285 12387 7343 12393
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 9030 12424 9036 12436
rect 8904 12396 9036 12424
rect 8904 12384 8910 12396
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 4338 12316 4344 12368
rect 4396 12356 4402 12368
rect 8202 12356 8208 12368
rect 4396 12328 8208 12356
rect 4396 12316 4402 12328
rect 8202 12316 8208 12328
rect 8260 12316 8266 12368
rect 5997 12291 6055 12297
rect 5997 12257 6009 12291
rect 6043 12288 6055 12291
rect 11146 12288 11152 12300
rect 6043 12260 11152 12288
rect 6043 12257 6055 12260
rect 5997 12251 6055 12257
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 6270 12180 6276 12232
rect 6328 12220 6334 12232
rect 6638 12220 6644 12232
rect 6328 12192 6644 12220
rect 6328 12180 6334 12192
rect 6638 12180 6644 12192
rect 6696 12220 6702 12232
rect 8297 12223 8355 12229
rect 8297 12220 8309 12223
rect 6696 12192 8309 12220
rect 6696 12180 6702 12192
rect 8297 12189 8309 12192
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 7837 12155 7895 12161
rect 7837 12152 7849 12155
rect 6972 12124 7849 12152
rect 6972 12112 6978 12124
rect 7837 12121 7849 12124
rect 7883 12121 7895 12155
rect 7837 12115 7895 12121
rect 8110 12112 8116 12164
rect 8168 12152 8174 12164
rect 8404 12152 8432 12183
rect 8168 12124 8432 12152
rect 8168 12112 8174 12124
rect 1104 11994 15824 12016
rect 1104 11942 3447 11994
rect 3499 11942 3511 11994
rect 3563 11942 3575 11994
rect 3627 11942 3639 11994
rect 3691 11942 8378 11994
rect 8430 11942 8442 11994
rect 8494 11942 8506 11994
rect 8558 11942 8570 11994
rect 8622 11942 13308 11994
rect 13360 11942 13372 11994
rect 13424 11942 13436 11994
rect 13488 11942 13500 11994
rect 13552 11942 15824 11994
rect 1104 11920 15824 11942
rect 8110 11880 8116 11892
rect 7484 11852 8116 11880
rect 7484 11753 7512 11852
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 9122 11880 9128 11892
rect 9083 11852 9128 11880
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11744 7527 11747
rect 7558 11744 7564 11756
rect 7515 11716 7564 11744
rect 7515 11713 7527 11716
rect 7469 11707 7527 11713
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 7282 11636 7288 11688
rect 7340 11676 7346 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 7340 11648 7757 11676
rect 7340 11636 7346 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 7745 11639 7803 11645
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 7190 11608 7196 11620
rect 4120 11580 7196 11608
rect 4120 11568 4126 11580
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 7926 11568 7932 11620
rect 7984 11617 7990 11620
rect 7984 11611 8048 11617
rect 7984 11577 8002 11611
rect 8036 11577 8048 11611
rect 7984 11571 8048 11577
rect 7984 11568 7990 11571
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6788 11512 6837 11540
rect 6788 11500 6794 11512
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7285 11543 7343 11549
rect 7285 11540 7297 11543
rect 7156 11512 7297 11540
rect 7156 11500 7162 11512
rect 7285 11509 7297 11512
rect 7331 11540 7343 11543
rect 8202 11540 8208 11552
rect 7331 11512 8208 11540
rect 7331 11509 7343 11512
rect 7285 11503 7343 11509
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 1104 11450 15824 11472
rect 1104 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 6104 11450
rect 6156 11398 10843 11450
rect 10895 11398 10907 11450
rect 10959 11398 10971 11450
rect 11023 11398 11035 11450
rect 11087 11398 15824 11450
rect 1104 11376 15824 11398
rect 6730 11336 6736 11348
rect 6691 11308 6736 11336
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 10134 11336 10140 11348
rect 10047 11308 10140 11336
rect 10134 11296 10140 11308
rect 10192 11336 10198 11348
rect 15470 11336 15476 11348
rect 10192 11308 15476 11336
rect 10192 11296 10198 11308
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 3142 11228 3148 11280
rect 3200 11268 3206 11280
rect 4157 11271 4215 11277
rect 4157 11268 4169 11271
rect 3200 11240 4169 11268
rect 3200 11228 3206 11240
rect 4157 11237 4169 11240
rect 4203 11237 4215 11271
rect 4157 11231 4215 11237
rect 4246 11228 4252 11280
rect 4304 11268 4310 11280
rect 6641 11271 6699 11277
rect 4304 11240 4349 11268
rect 4304 11228 4310 11240
rect 6641 11237 6653 11271
rect 6687 11268 6699 11271
rect 6914 11268 6920 11280
rect 6687 11240 6920 11268
rect 6687 11237 6699 11240
rect 6641 11231 6699 11237
rect 6914 11228 6920 11240
rect 6972 11228 6978 11280
rect 13630 11268 13636 11280
rect 7116 11240 13636 11268
rect 7116 11200 7144 11240
rect 13630 11228 13636 11240
rect 13688 11228 13694 11280
rect 7282 11200 7288 11212
rect 5184 11172 7144 11200
rect 7243 11172 7288 11200
rect 5184 11141 5212 11172
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 7558 11209 7564 11212
rect 7552 11200 7564 11209
rect 7519 11172 7564 11200
rect 7552 11163 7564 11172
rect 7558 11160 7564 11163
rect 7616 11160 7622 11212
rect 10042 11200 10048 11212
rect 10003 11172 10048 11200
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11101 5227 11135
rect 5169 11095 5227 11101
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 10229 11135 10287 11141
rect 6963 11104 7328 11132
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 6273 11067 6331 11073
rect 6273 11033 6285 11067
rect 6319 11064 6331 11067
rect 7190 11064 7196 11076
rect 6319 11036 7196 11064
rect 6319 11033 6331 11036
rect 6273 11027 6331 11033
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 7300 10996 7328 11104
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 10244 11064 10272 11095
rect 8772 11036 10272 11064
rect 8772 11008 8800 11036
rect 8665 10999 8723 11005
rect 8665 10996 8677 10999
rect 7300 10968 8677 10996
rect 8665 10965 8677 10968
rect 8711 10996 8723 10999
rect 8754 10996 8760 11008
rect 8711 10968 8760 10996
rect 8711 10965 8723 10968
rect 8665 10959 8723 10965
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 9674 10996 9680 11008
rect 9635 10968 9680 10996
rect 9674 10956 9680 10968
rect 9732 10956 9738 11008
rect 1104 10906 15824 10928
rect 1104 10854 3447 10906
rect 3499 10854 3511 10906
rect 3563 10854 3575 10906
rect 3627 10854 3639 10906
rect 3691 10854 8378 10906
rect 8430 10854 8442 10906
rect 8494 10854 8506 10906
rect 8558 10854 8570 10906
rect 8622 10854 13308 10906
rect 13360 10854 13372 10906
rect 13424 10854 13436 10906
rect 13488 10854 13500 10906
rect 13552 10854 15824 10906
rect 1104 10832 15824 10854
rect 2915 10795 2973 10801
rect 2915 10761 2927 10795
rect 2961 10792 2973 10795
rect 4246 10792 4252 10804
rect 2961 10764 4252 10792
rect 2961 10761 2973 10764
rect 2915 10755 2973 10761
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 7282 10792 7288 10804
rect 7243 10764 7288 10792
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 8846 10752 8852 10804
rect 8904 10792 8910 10804
rect 9490 10792 9496 10804
rect 8904 10764 9496 10792
rect 8904 10752 8910 10764
rect 9490 10752 9496 10764
rect 9548 10792 9554 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 9548 10764 10149 10792
rect 9548 10752 9554 10764
rect 10137 10761 10149 10764
rect 10183 10761 10195 10795
rect 10137 10755 10195 10761
rect 10226 10752 10232 10804
rect 10284 10792 10290 10804
rect 10686 10792 10692 10804
rect 10284 10764 10692 10792
rect 10284 10752 10290 10764
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 2774 10724 2780 10736
rect 2424 10696 2780 10724
rect 2424 10665 2452 10696
rect 2774 10684 2780 10696
rect 2832 10684 2838 10736
rect 2409 10659 2467 10665
rect 2409 10625 2421 10659
rect 2455 10625 2467 10659
rect 7300 10656 7328 10752
rect 8941 10727 8999 10733
rect 8941 10693 8953 10727
rect 8987 10693 8999 10727
rect 8941 10687 8999 10693
rect 7561 10659 7619 10665
rect 7561 10656 7573 10659
rect 2409 10619 2467 10625
rect 2608 10628 2912 10656
rect 7300 10628 7573 10656
rect 1489 10523 1547 10529
rect 1489 10489 1501 10523
rect 1535 10489 1547 10523
rect 1489 10483 1547 10489
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 2608 10520 2636 10628
rect 2884 10600 2912 10628
rect 7561 10625 7573 10628
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 8956 10656 8984 10687
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 8956 10628 9781 10656
rect 2866 10597 2872 10600
rect 2828 10591 2872 10597
rect 2828 10557 2840 10591
rect 2828 10551 2872 10557
rect 2866 10548 2872 10551
rect 2924 10548 2930 10600
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 7432 10560 7481 10588
rect 7432 10548 7438 10560
rect 7469 10557 7481 10560
rect 7515 10557 7527 10591
rect 7469 10551 7527 10557
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 8956 10588 8984 10628
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 10781 10659 10839 10665
rect 10781 10656 10793 10659
rect 9769 10619 9827 10625
rect 9876 10628 10793 10656
rect 7708 10560 8984 10588
rect 9585 10591 9643 10597
rect 7708 10548 7714 10560
rect 9585 10557 9597 10591
rect 9631 10588 9643 10591
rect 9674 10588 9680 10600
rect 9631 10560 9680 10588
rect 9631 10557 9643 10560
rect 9585 10551 9643 10557
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 1627 10492 2636 10520
rect 7828 10523 7886 10529
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 7828 10489 7840 10523
rect 7874 10520 7886 10523
rect 8754 10520 8760 10532
rect 7874 10492 8760 10520
rect 7874 10489 7886 10492
rect 7828 10483 7886 10489
rect 1504 10452 1532 10483
rect 8754 10480 8760 10492
rect 8812 10520 8818 10532
rect 9876 10520 9904 10628
rect 10781 10625 10793 10628
rect 10827 10625 10839 10659
rect 10781 10619 10839 10625
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10588 10655 10591
rect 10686 10588 10692 10600
rect 10643 10560 10692 10588
rect 10643 10557 10655 10560
rect 10597 10551 10655 10557
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 8812 10492 9904 10520
rect 10137 10523 10195 10529
rect 8812 10480 8818 10492
rect 10137 10489 10149 10523
rect 10183 10520 10195 10523
rect 10183 10492 10732 10520
rect 10183 10489 10195 10492
rect 10137 10483 10195 10489
rect 2958 10452 2964 10464
rect 1504 10424 2964 10452
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 9214 10452 9220 10464
rect 9175 10424 9220 10452
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 10704 10461 10732 10492
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10452 9735 10455
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 9723 10424 10241 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 10229 10415 10287 10421
rect 10689 10455 10747 10461
rect 10689 10421 10701 10455
rect 10735 10421 10747 10455
rect 10689 10415 10747 10421
rect 1104 10362 15824 10384
rect 1104 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 6104 10362
rect 6156 10310 10843 10362
rect 10895 10310 10907 10362
rect 10959 10310 10971 10362
rect 11023 10310 11035 10362
rect 11087 10310 15824 10362
rect 1104 10288 15824 10310
rect 6549 10251 6607 10257
rect 6549 10217 6561 10251
rect 6595 10248 6607 10251
rect 9214 10248 9220 10260
rect 6595 10220 9220 10248
rect 6595 10217 6607 10220
rect 6549 10211 6607 10217
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 9769 10251 9827 10257
rect 9769 10217 9781 10251
rect 9815 10248 9827 10251
rect 10042 10248 10048 10260
rect 9815 10220 10048 10248
rect 9815 10217 9827 10220
rect 9769 10211 9827 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 7460 10183 7518 10189
rect 7460 10149 7472 10183
rect 7506 10180 7518 10183
rect 7650 10180 7656 10192
rect 7506 10152 7656 10180
rect 7506 10149 7518 10152
rect 7460 10143 7518 10149
rect 7650 10140 7656 10152
rect 7708 10140 7714 10192
rect 6641 10115 6699 10121
rect 6641 10081 6653 10115
rect 6687 10112 6699 10115
rect 7098 10112 7104 10124
rect 6687 10084 7104 10112
rect 6687 10081 6699 10084
rect 6641 10075 6699 10081
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10112 7251 10115
rect 7282 10112 7288 10124
rect 7239 10084 7288 10112
rect 7239 10081 7251 10084
rect 7193 10075 7251 10081
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10013 6883 10047
rect 6825 10007 6883 10013
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 6181 9911 6239 9917
rect 6181 9908 6193 9911
rect 5592 9880 6193 9908
rect 5592 9868 5598 9880
rect 6181 9877 6193 9880
rect 6227 9877 6239 9911
rect 6840 9908 6868 10007
rect 7926 9908 7932 9920
rect 6840 9880 7932 9908
rect 6181 9871 6239 9877
rect 7926 9868 7932 9880
rect 7984 9908 7990 9920
rect 8573 9911 8631 9917
rect 8573 9908 8585 9911
rect 7984 9880 8585 9908
rect 7984 9868 7990 9880
rect 8573 9877 8585 9880
rect 8619 9877 8631 9911
rect 8573 9871 8631 9877
rect 1104 9818 15824 9840
rect 1104 9766 3447 9818
rect 3499 9766 3511 9818
rect 3563 9766 3575 9818
rect 3627 9766 3639 9818
rect 3691 9766 8378 9818
rect 8430 9766 8442 9818
rect 8494 9766 8506 9818
rect 8558 9766 8570 9818
rect 8622 9766 13308 9818
rect 13360 9766 13372 9818
rect 13424 9766 13436 9818
rect 13488 9766 13500 9818
rect 13552 9766 15824 9818
rect 1104 9744 15824 9766
rect 3326 9664 3332 9716
rect 3384 9704 3390 9716
rect 3786 9704 3792 9716
rect 3384 9676 3792 9704
rect 3384 9664 3390 9676
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 6730 9664 6736 9716
rect 6788 9704 6794 9716
rect 8018 9704 8024 9716
rect 6788 9676 8024 9704
rect 6788 9664 6794 9676
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 12066 9704 12072 9716
rect 11296 9676 12072 9704
rect 11296 9664 11302 9676
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 7098 9596 7104 9648
rect 7156 9636 7162 9648
rect 7193 9639 7251 9645
rect 7193 9636 7205 9639
rect 7156 9608 7205 9636
rect 7156 9596 7162 9608
rect 7193 9605 7205 9608
rect 7239 9605 7251 9639
rect 7193 9599 7251 9605
rect 7742 9568 7748 9580
rect 7703 9540 7748 9568
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 8662 9568 8668 9580
rect 8623 9540 8668 9568
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 8754 9528 8760 9580
rect 8812 9568 8818 9580
rect 8812 9540 8857 9568
rect 8812 9528 8818 9540
rect 4890 9460 4896 9512
rect 4948 9500 4954 9512
rect 6730 9500 6736 9512
rect 4948 9472 6736 9500
rect 4948 9460 4954 9472
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 7190 9460 7196 9512
rect 7248 9500 7254 9512
rect 7653 9503 7711 9509
rect 7653 9500 7665 9503
rect 7248 9472 7665 9500
rect 7248 9460 7254 9472
rect 7653 9469 7665 9472
rect 7699 9469 7711 9503
rect 7653 9463 7711 9469
rect 7561 9435 7619 9441
rect 7561 9401 7573 9435
rect 7607 9432 7619 9435
rect 7607 9404 8248 9432
rect 7607 9401 7619 9404
rect 7561 9395 7619 9401
rect 8220 9373 8248 9404
rect 8205 9367 8263 9373
rect 8205 9333 8217 9367
rect 8251 9333 8263 9367
rect 8205 9327 8263 9333
rect 8573 9367 8631 9373
rect 8573 9333 8585 9367
rect 8619 9364 8631 9367
rect 8754 9364 8760 9376
rect 8619 9336 8760 9364
rect 8619 9333 8631 9336
rect 8573 9327 8631 9333
rect 8754 9324 8760 9336
rect 8812 9364 8818 9376
rect 9398 9364 9404 9376
rect 8812 9336 9404 9364
rect 8812 9324 8818 9336
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 1104 9274 15824 9296
rect 1104 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 6104 9274
rect 6156 9222 10843 9274
rect 10895 9222 10907 9274
rect 10959 9222 10971 9274
rect 11023 9222 11035 9274
rect 11087 9222 15824 9274
rect 1104 9200 15824 9222
rect 12345 9027 12403 9033
rect 12345 8993 12357 9027
rect 12391 9024 12403 9027
rect 12434 9024 12440 9036
rect 12391 8996 12440 9024
rect 12391 8993 12403 8996
rect 12345 8987 12403 8993
rect 12434 8984 12440 8996
rect 12492 8984 12498 9036
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 12621 8959 12679 8965
rect 12621 8956 12633 8959
rect 11204 8928 12633 8956
rect 11204 8916 11210 8928
rect 12621 8925 12633 8928
rect 12667 8925 12679 8959
rect 12621 8919 12679 8925
rect 1104 8730 15824 8752
rect 1104 8678 3447 8730
rect 3499 8678 3511 8730
rect 3563 8678 3575 8730
rect 3627 8678 3639 8730
rect 3691 8678 8378 8730
rect 8430 8678 8442 8730
rect 8494 8678 8506 8730
rect 8558 8678 8570 8730
rect 8622 8678 13308 8730
rect 13360 8678 13372 8730
rect 13424 8678 13436 8730
rect 13488 8678 13500 8730
rect 13552 8678 15824 8730
rect 1104 8656 15824 8678
rect 1104 8186 15824 8208
rect 1104 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 6104 8186
rect 6156 8134 10843 8186
rect 10895 8134 10907 8186
rect 10959 8134 10971 8186
rect 11023 8134 11035 8186
rect 11087 8134 15824 8186
rect 1104 8112 15824 8134
rect 1104 7642 15824 7664
rect 1104 7590 3447 7642
rect 3499 7590 3511 7642
rect 3563 7590 3575 7642
rect 3627 7590 3639 7642
rect 3691 7590 8378 7642
rect 8430 7590 8442 7642
rect 8494 7590 8506 7642
rect 8558 7590 8570 7642
rect 8622 7590 13308 7642
rect 13360 7590 13372 7642
rect 13424 7590 13436 7642
rect 13488 7590 13500 7642
rect 13552 7590 15824 7642
rect 1104 7568 15824 7590
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 9030 7392 9036 7404
rect 5316 7364 9036 7392
rect 5316 7352 5322 7364
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 3237 7327 3295 7333
rect 3237 7293 3249 7327
rect 3283 7324 3295 7327
rect 5534 7324 5540 7336
rect 3283 7296 5540 7324
rect 3283 7293 3295 7296
rect 3237 7287 3295 7293
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 3050 7216 3056 7268
rect 3108 7256 3114 7268
rect 3513 7259 3571 7265
rect 3513 7256 3525 7259
rect 3108 7228 3525 7256
rect 3108 7216 3114 7228
rect 3513 7225 3525 7228
rect 3559 7225 3571 7259
rect 3513 7219 3571 7225
rect 3878 7148 3884 7200
rect 3936 7188 3942 7200
rect 7834 7188 7840 7200
rect 3936 7160 7840 7188
rect 3936 7148 3942 7160
rect 7834 7148 7840 7160
rect 7892 7148 7898 7200
rect 13906 7148 13912 7200
rect 13964 7188 13970 7200
rect 14642 7188 14648 7200
rect 13964 7160 14648 7188
rect 13964 7148 13970 7160
rect 14642 7148 14648 7160
rect 14700 7148 14706 7200
rect 1104 7098 15824 7120
rect 1104 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 6104 7098
rect 6156 7046 10843 7098
rect 10895 7046 10907 7098
rect 10959 7046 10971 7098
rect 11023 7046 11035 7098
rect 11087 7046 15824 7098
rect 1104 7024 15824 7046
rect 1104 6554 15824 6576
rect 1104 6502 3447 6554
rect 3499 6502 3511 6554
rect 3563 6502 3575 6554
rect 3627 6502 3639 6554
rect 3691 6502 8378 6554
rect 8430 6502 8442 6554
rect 8494 6502 8506 6554
rect 8558 6502 8570 6554
rect 8622 6502 13308 6554
rect 13360 6502 13372 6554
rect 13424 6502 13436 6554
rect 13488 6502 13500 6554
rect 13552 6502 15824 6554
rect 1104 6480 15824 6502
rect 7190 6128 7196 6180
rect 7248 6168 7254 6180
rect 10226 6168 10232 6180
rect 7248 6140 10232 6168
rect 7248 6128 7254 6140
rect 10226 6128 10232 6140
rect 10284 6128 10290 6180
rect 7374 6060 7380 6112
rect 7432 6100 7438 6112
rect 11606 6100 11612 6112
rect 7432 6072 11612 6100
rect 7432 6060 7438 6072
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 1104 6010 15824 6032
rect 1104 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 6104 6010
rect 6156 5958 10843 6010
rect 10895 5958 10907 6010
rect 10959 5958 10971 6010
rect 11023 5958 11035 6010
rect 11087 5958 15824 6010
rect 1104 5936 15824 5958
rect 4430 5856 4436 5908
rect 4488 5896 4494 5908
rect 8113 5899 8171 5905
rect 8113 5896 8125 5899
rect 4488 5868 8125 5896
rect 4488 5856 4494 5868
rect 8113 5865 8125 5868
rect 8159 5865 8171 5899
rect 8113 5859 8171 5865
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 7558 5828 7564 5840
rect 5184 5800 7564 5828
rect 4338 5760 4344 5772
rect 4299 5732 4344 5760
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 5184 5769 5212 5800
rect 7558 5788 7564 5800
rect 7616 5788 7622 5840
rect 9140 5828 9168 5859
rect 13906 5828 13912 5840
rect 7668 5800 9168 5828
rect 10244 5800 13912 5828
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5729 5227 5763
rect 5169 5723 5227 5729
rect 6825 5763 6883 5769
rect 6825 5729 6837 5763
rect 6871 5760 6883 5763
rect 7190 5760 7196 5772
rect 6871 5732 7196 5760
rect 6871 5729 6883 5732
rect 6825 5723 6883 5729
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 7374 5760 7380 5772
rect 7335 5732 7380 5760
rect 7374 5720 7380 5732
rect 7432 5720 7438 5772
rect 4798 5652 4804 5704
rect 4856 5692 4862 5704
rect 7668 5692 7696 5800
rect 7929 5763 7987 5769
rect 7929 5729 7941 5763
rect 7975 5760 7987 5763
rect 8846 5760 8852 5772
rect 7975 5732 8852 5760
rect 7975 5729 7987 5732
rect 7929 5723 7987 5729
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5760 8999 5763
rect 9122 5760 9128 5772
rect 8987 5732 9128 5760
rect 8987 5729 8999 5732
rect 8941 5723 8999 5729
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5760 9735 5763
rect 10134 5760 10140 5772
rect 9723 5732 10140 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 10134 5720 10140 5732
rect 10192 5720 10198 5772
rect 10244 5769 10272 5800
rect 13906 5788 13912 5800
rect 13964 5788 13970 5840
rect 10229 5763 10287 5769
rect 10229 5729 10241 5763
rect 10275 5729 10287 5763
rect 10229 5723 10287 5729
rect 11517 5763 11575 5769
rect 11517 5729 11529 5763
rect 11563 5760 11575 5763
rect 14458 5760 14464 5772
rect 11563 5732 14464 5760
rect 11563 5729 11575 5732
rect 11517 5723 11575 5729
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 4856 5664 7696 5692
rect 7760 5664 11744 5692
rect 4856 5652 4862 5664
rect 3786 5584 3792 5636
rect 3844 5624 3850 5636
rect 3844 5596 7144 5624
rect 3844 5584 3850 5596
rect 4522 5556 4528 5568
rect 4483 5528 4528 5556
rect 4522 5516 4528 5528
rect 4580 5516 4586 5568
rect 5350 5556 5356 5568
rect 5311 5528 5356 5556
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 7006 5556 7012 5568
rect 6967 5528 7012 5556
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 7116 5556 7144 5596
rect 7466 5584 7472 5636
rect 7524 5624 7530 5636
rect 7760 5624 7788 5664
rect 7524 5596 7788 5624
rect 7524 5584 7530 5596
rect 8018 5584 8024 5636
rect 8076 5624 8082 5636
rect 11716 5633 11744 5664
rect 9861 5627 9919 5633
rect 9861 5624 9873 5627
rect 8076 5596 9873 5624
rect 8076 5584 8082 5596
rect 9861 5593 9873 5596
rect 9907 5593 9919 5627
rect 9861 5587 9919 5593
rect 11701 5627 11759 5633
rect 11701 5593 11713 5627
rect 11747 5593 11759 5627
rect 11701 5587 11759 5593
rect 7561 5559 7619 5565
rect 7561 5556 7573 5559
rect 7116 5528 7573 5556
rect 7561 5525 7573 5528
rect 7607 5525 7619 5559
rect 7561 5519 7619 5525
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 10413 5559 10471 5565
rect 10413 5556 10425 5559
rect 9732 5528 10425 5556
rect 9732 5516 9738 5528
rect 10413 5525 10425 5528
rect 10459 5525 10471 5559
rect 10413 5519 10471 5525
rect 1104 5466 15824 5488
rect 1104 5414 3447 5466
rect 3499 5414 3511 5466
rect 3563 5414 3575 5466
rect 3627 5414 3639 5466
rect 3691 5414 8378 5466
rect 8430 5414 8442 5466
rect 8494 5414 8506 5466
rect 8558 5414 8570 5466
rect 8622 5414 13308 5466
rect 13360 5414 13372 5466
rect 13424 5414 13436 5466
rect 13488 5414 13500 5466
rect 13552 5414 15824 5466
rect 1104 5392 15824 5414
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 8481 5355 8539 5361
rect 8481 5352 8493 5355
rect 5500 5324 8493 5352
rect 5500 5312 5506 5324
rect 8481 5321 8493 5324
rect 8527 5321 8539 5355
rect 10134 5352 10140 5364
rect 8481 5315 8539 5321
rect 9692 5324 10140 5352
rect 9692 5284 9720 5324
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10318 5352 10324 5364
rect 10279 5324 10324 5352
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 11422 5352 11428 5364
rect 11383 5324 11428 5352
rect 11422 5312 11428 5324
rect 11480 5312 11486 5364
rect 11977 5355 12035 5361
rect 11977 5321 11989 5355
rect 12023 5352 12035 5355
rect 12158 5352 12164 5364
rect 12023 5324 12164 5352
rect 12023 5321 12035 5324
rect 11977 5315 12035 5321
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 8220 5256 9720 5284
rect 9769 5287 9827 5293
rect 3697 5151 3755 5157
rect 3697 5117 3709 5151
rect 3743 5148 3755 5151
rect 4062 5148 4068 5160
rect 3743 5120 4068 5148
rect 3743 5117 3755 5120
rect 3697 5111 3755 5117
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4801 5151 4859 5157
rect 4801 5117 4813 5151
rect 4847 5148 4859 5151
rect 5258 5148 5264 5160
rect 4847 5120 5264 5148
rect 4847 5117 4859 5120
rect 4801 5111 4859 5117
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 5718 5148 5724 5160
rect 5675 5120 5724 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 6181 5151 6239 5157
rect 6181 5117 6193 5151
rect 6227 5148 6239 5151
rect 6825 5151 6883 5157
rect 6227 5120 6684 5148
rect 6227 5117 6239 5120
rect 6181 5111 6239 5117
rect 2590 5040 2596 5092
rect 2648 5080 2654 5092
rect 6656 5080 6684 5120
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 6914 5148 6920 5160
rect 6871 5120 6920 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 8220 5148 8248 5256
rect 9769 5253 9781 5287
rect 9815 5284 9827 5287
rect 10410 5284 10416 5296
rect 9815 5256 10416 5284
rect 9815 5253 9827 5256
rect 9769 5247 9827 5253
rect 10410 5244 10416 5256
rect 10468 5244 10474 5296
rect 15930 5284 15936 5296
rect 11256 5256 15936 5284
rect 10318 5216 10324 5228
rect 8312 5188 10324 5216
rect 8312 5157 8340 5188
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 7423 5120 8248 5148
rect 8297 5151 8355 5157
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 8297 5117 8309 5151
rect 8343 5117 8355 5151
rect 8297 5111 8355 5117
rect 9033 5151 9091 5157
rect 9033 5117 9045 5151
rect 9079 5117 9091 5151
rect 9033 5111 9091 5117
rect 8110 5080 8116 5092
rect 2648 5052 6408 5080
rect 6656 5052 8116 5080
rect 2648 5040 2654 5052
rect 3878 5012 3884 5024
rect 3839 4984 3884 5012
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 4982 5012 4988 5024
rect 4943 4984 4988 5012
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 5810 5012 5816 5024
rect 5771 4984 5816 5012
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 6380 5021 6408 5052
rect 8110 5040 8116 5052
rect 8168 5040 8174 5092
rect 9048 5080 9076 5111
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 9585 5151 9643 5157
rect 9585 5148 9597 5151
rect 9456 5120 9597 5148
rect 9456 5108 9462 5120
rect 9585 5117 9597 5120
rect 9631 5117 9643 5151
rect 9585 5111 9643 5117
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 10100 5120 10149 5148
rect 10100 5108 10106 5120
rect 10137 5117 10149 5120
rect 10183 5117 10195 5151
rect 10137 5111 10195 5117
rect 10226 5108 10232 5160
rect 10284 5148 10290 5160
rect 10502 5148 10508 5160
rect 10284 5120 10508 5148
rect 10284 5108 10290 5120
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 11256 5157 11284 5256
rect 15930 5244 15936 5256
rect 15988 5244 15994 5296
rect 16298 5216 16304 5228
rect 11808 5188 16304 5216
rect 11808 5157 11836 5188
rect 16298 5176 16304 5188
rect 16356 5176 16362 5228
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5117 10747 5151
rect 10689 5111 10747 5117
rect 11241 5151 11299 5157
rect 11241 5117 11253 5151
rect 11287 5117 11299 5151
rect 11241 5111 11299 5117
rect 11793 5151 11851 5157
rect 11793 5117 11805 5151
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5117 12495 5151
rect 12986 5148 12992 5160
rect 12947 5120 12992 5148
rect 12437 5111 12495 5117
rect 10594 5080 10600 5092
rect 9048 5052 10600 5080
rect 10594 5040 10600 5052
rect 10652 5040 10658 5092
rect 10704 5080 10732 5111
rect 12452 5080 12480 5111
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 16758 5080 16764 5092
rect 10704 5052 11560 5080
rect 12452 5052 16764 5080
rect 6365 5015 6423 5021
rect 6365 4981 6377 5015
rect 6411 4981 6423 5015
rect 7006 5012 7012 5024
rect 6967 4984 7012 5012
rect 6365 4975 6423 4981
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 7558 5012 7564 5024
rect 7519 4984 7564 5012
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 9217 5015 9275 5021
rect 9217 5012 9229 5015
rect 7708 4984 9229 5012
rect 7708 4972 7714 4984
rect 9217 4981 9229 4984
rect 9263 4981 9275 5015
rect 9217 4975 9275 4981
rect 9766 4972 9772 5024
rect 9824 5012 9830 5024
rect 10873 5015 10931 5021
rect 10873 5012 10885 5015
rect 9824 4984 10885 5012
rect 9824 4972 9830 4984
rect 10873 4981 10885 4984
rect 10919 4981 10931 5015
rect 11532 5012 11560 5052
rect 16758 5040 16764 5052
rect 16816 5040 16822 5092
rect 12526 5012 12532 5024
rect 11532 4984 12532 5012
rect 10873 4975 10931 4981
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 12618 4972 12624 5024
rect 12676 5012 12682 5024
rect 13170 5012 13176 5024
rect 12676 4984 12721 5012
rect 13131 4984 13176 5012
rect 12676 4972 12682 4984
rect 13170 4972 13176 4984
rect 13228 4972 13234 5024
rect 1104 4922 15824 4944
rect 1104 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 6104 4922
rect 6156 4870 10843 4922
rect 10895 4870 10907 4922
rect 10959 4870 10971 4922
rect 11023 4870 11035 4922
rect 11087 4870 15824 4922
rect 1104 4848 15824 4870
rect 934 4768 940 4820
rect 992 4808 998 4820
rect 5077 4811 5135 4817
rect 5077 4808 5089 4811
rect 992 4780 5089 4808
rect 992 4768 998 4780
rect 5077 4777 5089 4780
rect 5123 4777 5135 4811
rect 5905 4811 5963 4817
rect 5905 4808 5917 4811
rect 5077 4771 5135 4777
rect 5184 4780 5917 4808
rect 2774 4700 2780 4752
rect 2832 4740 2838 4752
rect 5184 4740 5212 4780
rect 5905 4777 5917 4780
rect 5951 4777 5963 4811
rect 5905 4771 5963 4777
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 9217 4811 9275 4817
rect 9217 4808 9229 4811
rect 6880 4780 9229 4808
rect 6880 4768 6886 4780
rect 9217 4777 9229 4780
rect 9263 4777 9275 4811
rect 9217 4771 9275 4777
rect 9398 4768 9404 4820
rect 9456 4808 9462 4820
rect 9858 4808 9864 4820
rect 9456 4780 9720 4808
rect 9819 4780 9864 4808
rect 9456 4768 9462 4780
rect 2832 4712 5212 4740
rect 2832 4700 2838 4712
rect 5442 4700 5448 4752
rect 5500 4740 5506 4752
rect 7650 4740 7656 4752
rect 5500 4712 7656 4740
rect 5500 4700 5506 4712
rect 7650 4700 7656 4712
rect 7708 4700 7714 4752
rect 9582 4740 9588 4752
rect 7852 4712 9588 4740
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4672 4951 4675
rect 5626 4672 5632 4684
rect 4939 4644 5632 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 5721 4675 5779 4681
rect 5721 4641 5733 4675
rect 5767 4672 5779 4675
rect 6914 4672 6920 4684
rect 5767 4644 6920 4672
rect 5767 4641 5779 4644
rect 5721 4635 5779 4641
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7852 4681 7880 4712
rect 9582 4700 9588 4712
rect 9640 4700 9646 4752
rect 9692 4740 9720 4780
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 14182 4808 14188 4820
rect 10612 4780 14188 4808
rect 10612 4740 10640 4780
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 11974 4740 11980 4752
rect 9692 4712 10640 4740
rect 10704 4712 11980 4740
rect 7009 4675 7067 4681
rect 7009 4641 7021 4675
rect 7055 4641 7067 4675
rect 7009 4635 7067 4641
rect 7837 4675 7895 4681
rect 7837 4641 7849 4675
rect 7883 4641 7895 4675
rect 7837 4635 7895 4641
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4641 8447 4675
rect 8389 4635 8447 4641
rect 9033 4675 9091 4681
rect 9033 4641 9045 4675
rect 9079 4672 9091 4675
rect 9306 4672 9312 4684
rect 9079 4644 9312 4672
rect 9079 4641 9091 4644
rect 9033 4635 9091 4641
rect 7024 4604 7052 4635
rect 8294 4604 8300 4616
rect 7024 4576 8300 4604
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 6362 4496 6368 4548
rect 6420 4536 6426 4548
rect 8404 4536 8432 4635
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 10704 4681 10732 4712
rect 11974 4700 11980 4712
rect 12032 4700 12038 4752
rect 12158 4700 12164 4752
rect 12216 4740 12222 4752
rect 12618 4740 12624 4752
rect 12216 4712 12624 4740
rect 12216 4700 12222 4712
rect 12618 4700 12624 4712
rect 12676 4700 12682 4752
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4641 10747 4675
rect 10689 4635 10747 4641
rect 11885 4675 11943 4681
rect 11885 4641 11897 4675
rect 11931 4672 11943 4675
rect 13078 4672 13084 4684
rect 11931 4644 13084 4672
rect 11931 4641 11943 4644
rect 11885 4635 11943 4641
rect 9692 4604 9720 4635
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13722 4604 13728 4616
rect 9692 4576 13728 4604
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 12434 4536 12440 4548
rect 6420 4508 8156 4536
rect 8404 4508 12440 4536
rect 6420 4496 6426 4508
rect 6730 4428 6736 4480
rect 6788 4468 6794 4480
rect 7193 4471 7251 4477
rect 7193 4468 7205 4471
rect 6788 4440 7205 4468
rect 6788 4428 6794 4440
rect 7193 4437 7205 4440
rect 7239 4437 7251 4471
rect 7193 4431 7251 4437
rect 7834 4428 7840 4480
rect 7892 4468 7898 4480
rect 8021 4471 8079 4477
rect 8021 4468 8033 4471
rect 7892 4440 8033 4468
rect 7892 4428 7898 4440
rect 8021 4437 8033 4440
rect 8067 4437 8079 4471
rect 8128 4468 8156 4508
rect 12434 4496 12440 4508
rect 12492 4496 12498 4548
rect 8573 4471 8631 4477
rect 8573 4468 8585 4471
rect 8128 4440 8585 4468
rect 8021 4431 8079 4437
rect 8573 4437 8585 4440
rect 8619 4437 8631 4471
rect 10870 4468 10876 4480
rect 10831 4440 10876 4468
rect 8573 4431 8631 4437
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 12066 4468 12072 4480
rect 12027 4440 12072 4468
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 1104 4378 15824 4400
rect 1104 4326 3447 4378
rect 3499 4326 3511 4378
rect 3563 4326 3575 4378
rect 3627 4326 3639 4378
rect 3691 4326 8378 4378
rect 8430 4326 8442 4378
rect 8494 4326 8506 4378
rect 8558 4326 8570 4378
rect 8622 4326 13308 4378
rect 13360 4326 13372 4378
rect 13424 4326 13436 4378
rect 13488 4326 13500 4378
rect 13552 4326 15824 4378
rect 1104 4304 15824 4326
rect 5718 4224 5724 4276
rect 5776 4264 5782 4276
rect 9950 4264 9956 4276
rect 5776 4236 9956 4264
rect 5776 4224 5782 4236
rect 9950 4224 9956 4236
rect 10008 4224 10014 4276
rect 10226 4224 10232 4276
rect 10284 4264 10290 4276
rect 10284 4236 13768 4264
rect 10284 4224 10290 4236
rect 9490 4156 9496 4208
rect 9548 4196 9554 4208
rect 12158 4196 12164 4208
rect 9548 4168 12164 4196
rect 9548 4156 9554 4168
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 6546 4088 6552 4140
rect 6604 4128 6610 4140
rect 10870 4128 10876 4140
rect 6604 4100 10876 4128
rect 6604 4088 6610 4100
rect 10870 4088 10876 4100
rect 10928 4088 10934 4140
rect 13740 4128 13768 4236
rect 14642 4128 14648 4140
rect 13740 4100 14648 4128
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 3142 4020 3148 4072
rect 3200 4060 3206 4072
rect 7098 4060 7104 4072
rect 3200 4032 7104 4060
rect 3200 4020 3206 4032
rect 7098 4020 7104 4032
rect 7156 4020 7162 4072
rect 7745 4063 7803 4069
rect 7745 4029 7757 4063
rect 7791 4060 7803 4063
rect 9766 4060 9772 4072
rect 7791 4032 9772 4060
rect 7791 4029 7803 4032
rect 7745 4023 7803 4029
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4060 9919 4063
rect 13998 4060 14004 4072
rect 9907 4032 14004 4060
rect 9907 4029 9919 4032
rect 9861 4023 9919 4029
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 5718 3952 5724 4004
rect 5776 3992 5782 4004
rect 5776 3964 10088 3992
rect 5776 3952 5782 3964
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 10060 3933 10088 3964
rect 7929 3927 7987 3933
rect 7929 3924 7941 3927
rect 3844 3896 7941 3924
rect 3844 3884 3850 3896
rect 7929 3893 7941 3896
rect 7975 3893 7987 3927
rect 7929 3887 7987 3893
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3893 10103 3927
rect 10045 3887 10103 3893
rect 1104 3834 15824 3856
rect 1104 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 6104 3834
rect 6156 3782 10843 3834
rect 10895 3782 10907 3834
rect 10959 3782 10971 3834
rect 11023 3782 11035 3834
rect 11087 3782 15824 3834
rect 1104 3760 15824 3782
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 9122 3720 9128 3732
rect 5684 3692 9128 3720
rect 5684 3680 5690 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 11974 3720 11980 3732
rect 9640 3692 11980 3720
rect 9640 3680 9646 3692
rect 11974 3680 11980 3692
rect 12032 3680 12038 3732
rect 7834 3612 7840 3664
rect 7892 3652 7898 3664
rect 12066 3652 12072 3664
rect 7892 3624 12072 3652
rect 7892 3612 7898 3624
rect 12066 3612 12072 3624
rect 12124 3612 12130 3664
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 9950 3584 9956 3596
rect 6972 3556 9956 3584
rect 6972 3544 6978 3556
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 1394 3476 1400 3528
rect 1452 3516 1458 3528
rect 5810 3516 5816 3528
rect 1452 3488 5816 3516
rect 1452 3476 1458 3488
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 11238 3516 11244 3528
rect 8720 3488 11244 3516
rect 8720 3476 8726 3488
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 6822 3448 6828 3460
rect 5316 3420 6828 3448
rect 5316 3408 5322 3420
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 7926 3408 7932 3460
rect 7984 3448 7990 3460
rect 10410 3448 10416 3460
rect 7984 3420 10416 3448
rect 7984 3408 7990 3420
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 2682 3340 2688 3392
rect 2740 3380 2746 3392
rect 7558 3380 7564 3392
rect 2740 3352 7564 3380
rect 2740 3340 2746 3352
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 8202 3340 8208 3392
rect 8260 3380 8266 3392
rect 8662 3380 8668 3392
rect 8260 3352 8668 3380
rect 8260 3340 8266 3352
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 8754 3340 8760 3392
rect 8812 3380 8818 3392
rect 10502 3380 10508 3392
rect 8812 3352 10508 3380
rect 8812 3340 8818 3352
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 10594 3340 10600 3392
rect 10652 3380 10658 3392
rect 13078 3380 13084 3392
rect 10652 3352 13084 3380
rect 10652 3340 10658 3352
rect 13078 3340 13084 3352
rect 13136 3340 13142 3392
rect 1104 3290 15824 3312
rect 1104 3238 3447 3290
rect 3499 3238 3511 3290
rect 3563 3238 3575 3290
rect 3627 3238 3639 3290
rect 3691 3238 8378 3290
rect 8430 3238 8442 3290
rect 8494 3238 8506 3290
rect 8558 3238 8570 3290
rect 8622 3238 13308 3290
rect 13360 3238 13372 3290
rect 13424 3238 13436 3290
rect 13488 3238 13500 3290
rect 13552 3238 15824 3290
rect 1104 3216 15824 3238
rect 2314 3136 2320 3188
rect 2372 3176 2378 3188
rect 7006 3176 7012 3188
rect 2372 3148 7012 3176
rect 2372 3136 2378 3148
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 10686 3136 10692 3188
rect 10744 3176 10750 3188
rect 15470 3176 15476 3188
rect 10744 3148 15476 3176
rect 10744 3136 10750 3148
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 8202 3068 8208 3120
rect 8260 3108 8266 3120
rect 13170 3108 13176 3120
rect 8260 3080 13176 3108
rect 8260 3068 8266 3080
rect 13170 3068 13176 3080
rect 13228 3068 13234 3120
rect 1854 3000 1860 3052
rect 1912 3040 1918 3052
rect 5350 3040 5356 3052
rect 1912 3012 5356 3040
rect 1912 3000 1918 3012
rect 5350 3000 5356 3012
rect 5408 3000 5414 3052
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 9674 3040 9680 3052
rect 6328 3012 9680 3040
rect 6328 3000 6334 3012
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 12434 3040 12440 3052
rect 10376 3012 12440 3040
rect 10376 3000 10382 3012
rect 12434 3000 12440 3012
rect 12492 3000 12498 3052
rect 566 2932 572 2984
rect 624 2972 630 2984
rect 4982 2972 4988 2984
rect 624 2944 4988 2972
rect 624 2932 630 2944
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 8110 2932 8116 2984
rect 8168 2972 8174 2984
rect 10686 2972 10692 2984
rect 8168 2944 10692 2972
rect 8168 2932 8174 2944
rect 10686 2932 10692 2944
rect 10744 2932 10750 2984
rect 1026 2864 1032 2916
rect 1084 2904 1090 2916
rect 4522 2904 4528 2916
rect 1084 2876 4528 2904
rect 1084 2864 1090 2876
rect 4522 2864 4528 2876
rect 4580 2864 4586 2916
rect 6638 2864 6644 2916
rect 6696 2904 6702 2916
rect 9490 2904 9496 2916
rect 6696 2876 9496 2904
rect 6696 2864 6702 2876
rect 9490 2864 9496 2876
rect 9548 2864 9554 2916
rect 10502 2864 10508 2916
rect 10560 2904 10566 2916
rect 12894 2904 12900 2916
rect 10560 2876 12900 2904
rect 10560 2864 10566 2876
rect 12894 2864 12900 2876
rect 12952 2864 12958 2916
rect 198 2796 204 2848
rect 256 2836 262 2848
rect 3878 2836 3884 2848
rect 256 2808 3884 2836
rect 256 2796 262 2808
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 12526 2796 12532 2848
rect 12584 2836 12590 2848
rect 15010 2836 15016 2848
rect 12584 2808 15016 2836
rect 12584 2796 12590 2808
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 1104 2746 15824 2768
rect 1104 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 6104 2746
rect 6156 2694 10843 2746
rect 10895 2694 10907 2746
rect 10959 2694 10971 2746
rect 11023 2694 11035 2746
rect 11087 2694 15824 2746
rect 1104 2672 15824 2694
rect 1104 2202 15824 2224
rect 1104 2150 3447 2202
rect 3499 2150 3511 2202
rect 3563 2150 3575 2202
rect 3627 2150 3639 2202
rect 3691 2150 8378 2202
rect 8430 2150 8442 2202
rect 8494 2150 8506 2202
rect 8558 2150 8570 2202
rect 8622 2150 13308 2202
rect 13360 2150 13372 2202
rect 13424 2150 13436 2202
rect 13488 2150 13500 2202
rect 13552 2150 15824 2202
rect 1104 2128 15824 2150
rect 7006 2048 7012 2100
rect 7064 2088 7070 2100
rect 8018 2088 8024 2100
rect 7064 2060 8024 2088
rect 7064 2048 7070 2060
rect 8018 2048 8024 2060
rect 8076 2048 8082 2100
rect 3970 552 3976 604
rect 4028 592 4034 604
rect 6362 592 6368 604
rect 4028 564 6368 592
rect 4028 552 4034 564
rect 6362 552 6368 564
rect 6420 552 6426 604
<< via1 >>
rect 3056 17892 3108 17944
rect 4896 17892 4948 17944
rect 3447 17382 3499 17434
rect 3511 17382 3563 17434
rect 3575 17382 3627 17434
rect 3639 17382 3691 17434
rect 8378 17382 8430 17434
rect 8442 17382 8494 17434
rect 8506 17382 8558 17434
rect 8570 17382 8622 17434
rect 13308 17382 13360 17434
rect 13372 17382 13424 17434
rect 13436 17382 13488 17434
rect 13500 17382 13552 17434
rect 5912 16838 5964 16890
rect 5976 16838 6028 16890
rect 6040 16838 6092 16890
rect 6104 16838 6156 16890
rect 10843 16838 10895 16890
rect 10907 16838 10959 16890
rect 10971 16838 11023 16890
rect 11035 16838 11087 16890
rect 6276 16532 6328 16584
rect 10416 16532 10468 16584
rect 5540 16464 5592 16516
rect 9956 16464 10008 16516
rect 6368 16396 6420 16448
rect 10324 16396 10376 16448
rect 3447 16294 3499 16346
rect 3511 16294 3563 16346
rect 3575 16294 3627 16346
rect 3639 16294 3691 16346
rect 8378 16294 8430 16346
rect 8442 16294 8494 16346
rect 8506 16294 8558 16346
rect 8570 16294 8622 16346
rect 13308 16294 13360 16346
rect 13372 16294 13424 16346
rect 13436 16294 13488 16346
rect 13500 16294 13552 16346
rect 7656 16192 7708 16244
rect 10508 16192 10560 16244
rect 6828 16124 6880 16176
rect 9772 16124 9824 16176
rect 7288 16056 7340 16108
rect 8852 16056 8904 16108
rect 10508 16056 10560 16108
rect 11336 16056 11388 16108
rect 8668 15988 8720 16040
rect 9588 15988 9640 16040
rect 10692 15988 10744 16040
rect 11796 15988 11848 16040
rect 13084 15988 13136 16040
rect 16304 15988 16356 16040
rect 8208 15920 8260 15972
rect 9680 15920 9732 15972
rect 1860 15852 1912 15904
rect 2688 15852 2740 15904
rect 4344 15852 4396 15904
rect 5356 15852 5408 15904
rect 9312 15852 9364 15904
rect 13820 15920 13872 15972
rect 9864 15852 9916 15904
rect 13176 15852 13228 15904
rect 5912 15750 5964 15802
rect 5976 15750 6028 15802
rect 6040 15750 6092 15802
rect 6104 15750 6156 15802
rect 10843 15750 10895 15802
rect 10907 15750 10959 15802
rect 10971 15750 11023 15802
rect 11035 15750 11087 15802
rect 572 15648 624 15700
rect 7104 15648 7156 15700
rect 9496 15648 9548 15700
rect 12992 15648 13044 15700
rect 6276 15580 6328 15632
rect 9220 15580 9272 15632
rect 9864 15580 9916 15632
rect 7840 15512 7892 15564
rect 8024 15512 8076 15564
rect 10600 15512 10652 15564
rect 2228 15444 2280 15496
rect 1400 15376 1452 15428
rect 7748 15444 7800 15496
rect 11428 15444 11480 15496
rect 11980 15444 12032 15496
rect 15108 15512 15160 15564
rect 14464 15444 14516 15496
rect 15936 15444 15988 15496
rect 8116 15376 8168 15428
rect 12164 15376 12216 15428
rect 12992 15376 13044 15428
rect 16764 15376 16816 15428
rect 4712 15308 4764 15360
rect 6828 15308 6880 15360
rect 7196 15308 7248 15360
rect 9404 15308 9456 15360
rect 3447 15206 3499 15258
rect 3511 15206 3563 15258
rect 3575 15206 3627 15258
rect 3639 15206 3691 15258
rect 8378 15206 8430 15258
rect 8442 15206 8494 15258
rect 8506 15206 8558 15258
rect 8570 15206 8622 15258
rect 13308 15206 13360 15258
rect 13372 15206 13424 15258
rect 13436 15206 13488 15258
rect 13500 15206 13552 15258
rect 6828 15104 6880 15156
rect 9404 15147 9456 15156
rect 9404 15113 9413 15147
rect 9413 15113 9447 15147
rect 9447 15113 9456 15147
rect 9404 15104 9456 15113
rect 10600 14900 10652 14952
rect 9404 14832 9456 14884
rect 5912 14662 5964 14714
rect 5976 14662 6028 14714
rect 6040 14662 6092 14714
rect 6104 14662 6156 14714
rect 10843 14662 10895 14714
rect 10907 14662 10959 14714
rect 10971 14662 11023 14714
rect 11035 14662 11087 14714
rect 3447 14118 3499 14170
rect 3511 14118 3563 14170
rect 3575 14118 3627 14170
rect 3639 14118 3691 14170
rect 8378 14118 8430 14170
rect 8442 14118 8494 14170
rect 8506 14118 8558 14170
rect 8570 14118 8622 14170
rect 13308 14118 13360 14170
rect 13372 14118 13424 14170
rect 13436 14118 13488 14170
rect 13500 14118 13552 14170
rect 13728 14016 13780 14068
rect 8116 13948 8168 14000
rect 3976 13880 4028 13932
rect 4252 13855 4304 13864
rect 4252 13821 4261 13855
rect 4261 13821 4295 13855
rect 4295 13821 4304 13855
rect 4252 13812 4304 13821
rect 13636 13812 13688 13864
rect 5912 13574 5964 13626
rect 5976 13574 6028 13626
rect 6040 13574 6092 13626
rect 6104 13574 6156 13626
rect 10843 13574 10895 13626
rect 10907 13574 10959 13626
rect 10971 13574 11023 13626
rect 11035 13574 11087 13626
rect 4252 13472 4304 13524
rect 204 13336 256 13388
rect 4988 13379 5040 13388
rect 4988 13345 4997 13379
rect 4997 13345 5031 13379
rect 5031 13345 5040 13379
rect 4988 13336 5040 13345
rect 9128 13268 9180 13320
rect 2872 13132 2924 13184
rect 3447 13030 3499 13082
rect 3511 13030 3563 13082
rect 3575 13030 3627 13082
rect 3639 13030 3691 13082
rect 8378 13030 8430 13082
rect 8442 13030 8494 13082
rect 8506 13030 8558 13082
rect 8570 13030 8622 13082
rect 13308 13030 13360 13082
rect 13372 13030 13424 13082
rect 13436 13030 13488 13082
rect 13500 13030 13552 13082
rect 8668 12860 8720 12912
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 7840 12724 7892 12776
rect 7656 12656 7708 12708
rect 9128 12588 9180 12640
rect 13452 12588 13504 12640
rect 5912 12486 5964 12538
rect 5976 12486 6028 12538
rect 6040 12486 6092 12538
rect 6104 12486 6156 12538
rect 10843 12486 10895 12538
rect 10907 12486 10959 12538
rect 10971 12486 11023 12538
rect 11035 12486 11087 12538
rect 4988 12384 5040 12436
rect 7380 12384 7432 12436
rect 8852 12384 8904 12436
rect 9036 12384 9088 12436
rect 4344 12316 4396 12368
rect 8208 12359 8260 12368
rect 8208 12325 8217 12359
rect 8217 12325 8251 12359
rect 8251 12325 8260 12359
rect 8208 12316 8260 12325
rect 11152 12248 11204 12300
rect 6276 12180 6328 12232
rect 6644 12180 6696 12232
rect 6920 12112 6972 12164
rect 8116 12112 8168 12164
rect 3447 11942 3499 11994
rect 3511 11942 3563 11994
rect 3575 11942 3627 11994
rect 3639 11942 3691 11994
rect 8378 11942 8430 11994
rect 8442 11942 8494 11994
rect 8506 11942 8558 11994
rect 8570 11942 8622 11994
rect 13308 11942 13360 11994
rect 13372 11942 13424 11994
rect 13436 11942 13488 11994
rect 13500 11942 13552 11994
rect 8116 11840 8168 11892
rect 9128 11883 9180 11892
rect 9128 11849 9137 11883
rect 9137 11849 9171 11883
rect 9171 11849 9180 11883
rect 9128 11840 9180 11849
rect 7564 11704 7616 11756
rect 7288 11636 7340 11688
rect 4068 11568 4120 11620
rect 7196 11611 7248 11620
rect 7196 11577 7205 11611
rect 7205 11577 7239 11611
rect 7239 11577 7248 11611
rect 7196 11568 7248 11577
rect 7932 11568 7984 11620
rect 6736 11500 6788 11552
rect 7104 11500 7156 11552
rect 8208 11500 8260 11552
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 6104 11398 6156 11450
rect 10843 11398 10895 11450
rect 10907 11398 10959 11450
rect 10971 11398 11023 11450
rect 11035 11398 11087 11450
rect 6736 11339 6788 11348
rect 6736 11305 6745 11339
rect 6745 11305 6779 11339
rect 6779 11305 6788 11339
rect 6736 11296 6788 11305
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 15476 11296 15528 11348
rect 3148 11228 3200 11280
rect 4252 11271 4304 11280
rect 4252 11237 4261 11271
rect 4261 11237 4295 11271
rect 4295 11237 4304 11271
rect 4252 11228 4304 11237
rect 6920 11228 6972 11280
rect 13636 11228 13688 11280
rect 7288 11203 7340 11212
rect 7288 11169 7297 11203
rect 7297 11169 7331 11203
rect 7331 11169 7340 11203
rect 7288 11160 7340 11169
rect 7564 11203 7616 11212
rect 7564 11169 7598 11203
rect 7598 11169 7616 11203
rect 7564 11160 7616 11169
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 7196 11024 7248 11076
rect 8760 10956 8812 11008
rect 9680 10999 9732 11008
rect 9680 10965 9689 10999
rect 9689 10965 9723 10999
rect 9723 10965 9732 10999
rect 9680 10956 9732 10965
rect 3447 10854 3499 10906
rect 3511 10854 3563 10906
rect 3575 10854 3627 10906
rect 3639 10854 3691 10906
rect 8378 10854 8430 10906
rect 8442 10854 8494 10906
rect 8506 10854 8558 10906
rect 8570 10854 8622 10906
rect 13308 10854 13360 10906
rect 13372 10854 13424 10906
rect 13436 10854 13488 10906
rect 13500 10854 13552 10906
rect 4252 10752 4304 10804
rect 7288 10795 7340 10804
rect 7288 10761 7297 10795
rect 7297 10761 7331 10795
rect 7331 10761 7340 10795
rect 7288 10752 7340 10761
rect 8852 10752 8904 10804
rect 9496 10752 9548 10804
rect 10232 10752 10284 10804
rect 10692 10752 10744 10804
rect 2780 10684 2832 10736
rect 2872 10591 2924 10600
rect 2872 10557 2874 10591
rect 2874 10557 2924 10591
rect 2872 10548 2924 10557
rect 7380 10548 7432 10600
rect 7656 10548 7708 10600
rect 9680 10548 9732 10600
rect 8760 10480 8812 10532
rect 10692 10548 10744 10600
rect 2964 10412 3016 10464
rect 9220 10455 9272 10464
rect 9220 10421 9229 10455
rect 9229 10421 9263 10455
rect 9263 10421 9272 10455
rect 9220 10412 9272 10421
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 6104 10310 6156 10362
rect 10843 10310 10895 10362
rect 10907 10310 10959 10362
rect 10971 10310 11023 10362
rect 11035 10310 11087 10362
rect 9220 10208 9272 10260
rect 10048 10208 10100 10260
rect 7656 10140 7708 10192
rect 7104 10072 7156 10124
rect 7288 10072 7340 10124
rect 5540 9868 5592 9920
rect 7932 9868 7984 9920
rect 3447 9766 3499 9818
rect 3511 9766 3563 9818
rect 3575 9766 3627 9818
rect 3639 9766 3691 9818
rect 8378 9766 8430 9818
rect 8442 9766 8494 9818
rect 8506 9766 8558 9818
rect 8570 9766 8622 9818
rect 13308 9766 13360 9818
rect 13372 9766 13424 9818
rect 13436 9766 13488 9818
rect 13500 9766 13552 9818
rect 3332 9664 3384 9716
rect 3792 9664 3844 9716
rect 6736 9664 6788 9716
rect 8024 9664 8076 9716
rect 11244 9664 11296 9716
rect 12072 9664 12124 9716
rect 7104 9596 7156 9648
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 8760 9571 8812 9580
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 4896 9460 4948 9512
rect 6736 9460 6788 9512
rect 7196 9460 7248 9512
rect 8760 9324 8812 9376
rect 9404 9324 9456 9376
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 6104 9222 6156 9274
rect 10843 9222 10895 9274
rect 10907 9222 10959 9274
rect 10971 9222 11023 9274
rect 11035 9222 11087 9274
rect 12440 8984 12492 9036
rect 11152 8916 11204 8968
rect 3447 8678 3499 8730
rect 3511 8678 3563 8730
rect 3575 8678 3627 8730
rect 3639 8678 3691 8730
rect 8378 8678 8430 8730
rect 8442 8678 8494 8730
rect 8506 8678 8558 8730
rect 8570 8678 8622 8730
rect 13308 8678 13360 8730
rect 13372 8678 13424 8730
rect 13436 8678 13488 8730
rect 13500 8678 13552 8730
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 6104 8134 6156 8186
rect 10843 8134 10895 8186
rect 10907 8134 10959 8186
rect 10971 8134 11023 8186
rect 11035 8134 11087 8186
rect 3447 7590 3499 7642
rect 3511 7590 3563 7642
rect 3575 7590 3627 7642
rect 3639 7590 3691 7642
rect 8378 7590 8430 7642
rect 8442 7590 8494 7642
rect 8506 7590 8558 7642
rect 8570 7590 8622 7642
rect 13308 7590 13360 7642
rect 13372 7590 13424 7642
rect 13436 7590 13488 7642
rect 13500 7590 13552 7642
rect 5264 7352 5316 7404
rect 9036 7352 9088 7404
rect 5540 7284 5592 7336
rect 3056 7216 3108 7268
rect 3884 7148 3936 7200
rect 7840 7148 7892 7200
rect 13912 7148 13964 7200
rect 14648 7148 14700 7200
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 6104 7046 6156 7098
rect 10843 7046 10895 7098
rect 10907 7046 10959 7098
rect 10971 7046 11023 7098
rect 11035 7046 11087 7098
rect 3447 6502 3499 6554
rect 3511 6502 3563 6554
rect 3575 6502 3627 6554
rect 3639 6502 3691 6554
rect 8378 6502 8430 6554
rect 8442 6502 8494 6554
rect 8506 6502 8558 6554
rect 8570 6502 8622 6554
rect 13308 6502 13360 6554
rect 13372 6502 13424 6554
rect 13436 6502 13488 6554
rect 13500 6502 13552 6554
rect 7196 6128 7248 6180
rect 10232 6128 10284 6180
rect 7380 6060 7432 6112
rect 11612 6060 11664 6112
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 6104 5958 6156 6010
rect 10843 5958 10895 6010
rect 10907 5958 10959 6010
rect 10971 5958 11023 6010
rect 11035 5958 11087 6010
rect 4436 5856 4488 5908
rect 4344 5763 4396 5772
rect 4344 5729 4353 5763
rect 4353 5729 4387 5763
rect 4387 5729 4396 5763
rect 4344 5720 4396 5729
rect 7564 5788 7616 5840
rect 7196 5720 7248 5772
rect 7380 5763 7432 5772
rect 7380 5729 7389 5763
rect 7389 5729 7423 5763
rect 7423 5729 7432 5763
rect 7380 5720 7432 5729
rect 4804 5652 4856 5704
rect 8852 5720 8904 5772
rect 9128 5720 9180 5772
rect 10140 5720 10192 5772
rect 13912 5788 13964 5840
rect 14464 5720 14516 5772
rect 3792 5584 3844 5636
rect 4528 5559 4580 5568
rect 4528 5525 4537 5559
rect 4537 5525 4571 5559
rect 4571 5525 4580 5559
rect 4528 5516 4580 5525
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 7472 5584 7524 5636
rect 8024 5584 8076 5636
rect 9680 5516 9732 5568
rect 3447 5414 3499 5466
rect 3511 5414 3563 5466
rect 3575 5414 3627 5466
rect 3639 5414 3691 5466
rect 8378 5414 8430 5466
rect 8442 5414 8494 5466
rect 8506 5414 8558 5466
rect 8570 5414 8622 5466
rect 13308 5414 13360 5466
rect 13372 5414 13424 5466
rect 13436 5414 13488 5466
rect 13500 5414 13552 5466
rect 5448 5312 5500 5364
rect 10140 5312 10192 5364
rect 10324 5355 10376 5364
rect 10324 5321 10333 5355
rect 10333 5321 10367 5355
rect 10367 5321 10376 5355
rect 10324 5312 10376 5321
rect 11428 5355 11480 5364
rect 11428 5321 11437 5355
rect 11437 5321 11471 5355
rect 11471 5321 11480 5355
rect 11428 5312 11480 5321
rect 12164 5312 12216 5364
rect 4068 5108 4120 5160
rect 5264 5108 5316 5160
rect 5724 5108 5776 5160
rect 2596 5040 2648 5092
rect 6920 5108 6972 5160
rect 10416 5244 10468 5296
rect 10324 5176 10376 5228
rect 3884 5015 3936 5024
rect 3884 4981 3893 5015
rect 3893 4981 3927 5015
rect 3927 4981 3936 5015
rect 3884 4972 3936 4981
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 4988 4972 5040 4981
rect 5816 5015 5868 5024
rect 5816 4981 5825 5015
rect 5825 4981 5859 5015
rect 5859 4981 5868 5015
rect 5816 4972 5868 4981
rect 8116 5040 8168 5092
rect 9404 5108 9456 5160
rect 10048 5108 10100 5160
rect 10232 5108 10284 5160
rect 10508 5108 10560 5160
rect 15936 5244 15988 5296
rect 16304 5176 16356 5228
rect 12992 5151 13044 5160
rect 10600 5040 10652 5092
rect 12992 5117 13001 5151
rect 13001 5117 13035 5151
rect 13035 5117 13044 5151
rect 12992 5108 13044 5117
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 7564 5015 7616 5024
rect 7564 4981 7573 5015
rect 7573 4981 7607 5015
rect 7607 4981 7616 5015
rect 7564 4972 7616 4981
rect 7656 4972 7708 5024
rect 9772 4972 9824 5024
rect 16764 5040 16816 5092
rect 12532 4972 12584 5024
rect 12624 5015 12676 5024
rect 12624 4981 12633 5015
rect 12633 4981 12667 5015
rect 12667 4981 12676 5015
rect 13176 5015 13228 5024
rect 12624 4972 12676 4981
rect 13176 4981 13185 5015
rect 13185 4981 13219 5015
rect 13219 4981 13228 5015
rect 13176 4972 13228 4981
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 6104 4870 6156 4922
rect 10843 4870 10895 4922
rect 10907 4870 10959 4922
rect 10971 4870 11023 4922
rect 11035 4870 11087 4922
rect 940 4768 992 4820
rect 2780 4700 2832 4752
rect 6828 4768 6880 4820
rect 9404 4768 9456 4820
rect 9864 4811 9916 4820
rect 5448 4700 5500 4752
rect 7656 4700 7708 4752
rect 5632 4632 5684 4684
rect 6920 4632 6972 4684
rect 9588 4700 9640 4752
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 14188 4768 14240 4820
rect 8300 4564 8352 4616
rect 6368 4496 6420 4548
rect 9312 4632 9364 4684
rect 11980 4700 12032 4752
rect 12164 4700 12216 4752
rect 12624 4700 12676 4752
rect 13084 4632 13136 4684
rect 13728 4564 13780 4616
rect 6736 4428 6788 4480
rect 7840 4428 7892 4480
rect 12440 4496 12492 4548
rect 10876 4471 10928 4480
rect 10876 4437 10885 4471
rect 10885 4437 10919 4471
rect 10919 4437 10928 4471
rect 10876 4428 10928 4437
rect 12072 4471 12124 4480
rect 12072 4437 12081 4471
rect 12081 4437 12115 4471
rect 12115 4437 12124 4471
rect 12072 4428 12124 4437
rect 3447 4326 3499 4378
rect 3511 4326 3563 4378
rect 3575 4326 3627 4378
rect 3639 4326 3691 4378
rect 8378 4326 8430 4378
rect 8442 4326 8494 4378
rect 8506 4326 8558 4378
rect 8570 4326 8622 4378
rect 13308 4326 13360 4378
rect 13372 4326 13424 4378
rect 13436 4326 13488 4378
rect 13500 4326 13552 4378
rect 5724 4224 5776 4276
rect 9956 4224 10008 4276
rect 10232 4224 10284 4276
rect 9496 4156 9548 4208
rect 12164 4156 12216 4208
rect 6552 4088 6604 4140
rect 10876 4088 10928 4140
rect 14648 4088 14700 4140
rect 3148 4020 3200 4072
rect 7104 4020 7156 4072
rect 9772 4020 9824 4072
rect 14004 4020 14056 4072
rect 5724 3952 5776 4004
rect 3792 3884 3844 3936
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 6104 3782 6156 3834
rect 10843 3782 10895 3834
rect 10907 3782 10959 3834
rect 10971 3782 11023 3834
rect 11035 3782 11087 3834
rect 5632 3680 5684 3732
rect 9128 3680 9180 3732
rect 9588 3680 9640 3732
rect 11980 3680 12032 3732
rect 7840 3612 7892 3664
rect 12072 3612 12124 3664
rect 6920 3544 6972 3596
rect 9956 3544 10008 3596
rect 1400 3476 1452 3528
rect 5816 3476 5868 3528
rect 8668 3476 8720 3528
rect 11244 3476 11296 3528
rect 5264 3408 5316 3460
rect 6828 3408 6880 3460
rect 7932 3408 7984 3460
rect 10416 3408 10468 3460
rect 2688 3340 2740 3392
rect 7564 3340 7616 3392
rect 8208 3340 8260 3392
rect 8668 3340 8720 3392
rect 8760 3340 8812 3392
rect 10508 3340 10560 3392
rect 10600 3340 10652 3392
rect 13084 3340 13136 3392
rect 3447 3238 3499 3290
rect 3511 3238 3563 3290
rect 3575 3238 3627 3290
rect 3639 3238 3691 3290
rect 8378 3238 8430 3290
rect 8442 3238 8494 3290
rect 8506 3238 8558 3290
rect 8570 3238 8622 3290
rect 13308 3238 13360 3290
rect 13372 3238 13424 3290
rect 13436 3238 13488 3290
rect 13500 3238 13552 3290
rect 2320 3136 2372 3188
rect 7012 3136 7064 3188
rect 10692 3136 10744 3188
rect 15476 3136 15528 3188
rect 8208 3068 8260 3120
rect 13176 3068 13228 3120
rect 1860 3000 1912 3052
rect 5356 3000 5408 3052
rect 6276 3000 6328 3052
rect 9680 3000 9732 3052
rect 10324 3000 10376 3052
rect 12440 3000 12492 3052
rect 572 2932 624 2984
rect 4988 2932 5040 2984
rect 8116 2932 8168 2984
rect 10692 2932 10744 2984
rect 1032 2864 1084 2916
rect 4528 2864 4580 2916
rect 6644 2864 6696 2916
rect 9496 2864 9548 2916
rect 10508 2864 10560 2916
rect 12900 2864 12952 2916
rect 204 2796 256 2848
rect 3884 2796 3936 2848
rect 12532 2796 12584 2848
rect 15016 2796 15068 2848
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 6104 2694 6156 2746
rect 10843 2694 10895 2746
rect 10907 2694 10959 2746
rect 10971 2694 11023 2746
rect 11035 2694 11087 2746
rect 3447 2150 3499 2202
rect 3511 2150 3563 2202
rect 3575 2150 3627 2202
rect 3639 2150 3691 2202
rect 8378 2150 8430 2202
rect 8442 2150 8494 2202
rect 8506 2150 8558 2202
rect 8570 2150 8622 2202
rect 13308 2150 13360 2202
rect 13372 2150 13424 2202
rect 13436 2150 13488 2202
rect 13500 2150 13552 2202
rect 7012 2048 7064 2100
rect 8024 2048 8076 2100
rect 3976 552 4028 604
rect 6368 552 6420 604
<< metal2 >>
rect 202 19520 258 20000
rect 570 19520 626 20000
rect 1030 19520 1086 20000
rect 1398 19520 1454 20000
rect 1858 19520 1914 20000
rect 2226 19520 2282 20000
rect 2686 19520 2742 20000
rect 3054 19520 3110 20000
rect 3514 19520 3570 20000
rect 3882 19520 3938 20000
rect 4342 19520 4398 20000
rect 4710 19520 4766 20000
rect 5170 19520 5226 20000
rect 5538 19520 5594 20000
rect 5998 19520 6054 20000
rect 6366 19520 6422 20000
rect 6826 19520 6882 20000
rect 7194 19520 7250 20000
rect 7654 19520 7710 20000
rect 8022 19520 8078 20000
rect 8482 19520 8538 20000
rect 8850 19520 8906 20000
rect 9310 19520 9366 20000
rect 9678 19520 9734 20000
rect 10138 19520 10194 20000
rect 10506 19520 10562 20000
rect 10966 19520 11022 20000
rect 11334 19520 11390 20000
rect 11794 19520 11850 20000
rect 12162 19520 12218 20000
rect 12622 19520 12678 20000
rect 12990 19520 13046 20000
rect 13450 19520 13506 20000
rect 13818 19520 13874 20000
rect 14278 19530 14334 20000
rect 14016 19520 14334 19530
rect 14646 19520 14702 20000
rect 15106 19520 15162 20000
rect 15474 19520 15530 20000
rect 15934 19520 15990 20000
rect 16302 19520 16358 20000
rect 16762 19520 16818 20000
rect 216 13394 244 19520
rect 584 15706 612 19520
rect 572 15700 624 15706
rect 572 15642 624 15648
rect 204 13388 256 13394
rect 204 13330 256 13336
rect 1044 12458 1072 19520
rect 1412 15434 1440 19520
rect 1872 15910 1900 19520
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 2240 15502 2268 19520
rect 2700 15994 2728 19520
rect 3068 17950 3096 19520
rect 3056 17944 3108 17950
rect 3056 17886 3108 17892
rect 3528 17626 3556 19520
rect 2608 15966 2728 15994
rect 3344 17598 3556 17626
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 1400 15428 1452 15434
rect 1400 15370 1452 15376
rect 952 12430 1072 12458
rect 952 4826 980 12430
rect 2608 5098 2636 15966
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 940 4820 992 4826
rect 940 4762 992 4768
rect 2700 4740 2728 15846
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 10742 2820 14991
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 2884 10606 2912 13126
rect 3146 11656 3202 11665
rect 3146 11591 3202 11600
rect 3160 11286 3188 11591
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 2872 10600 2924 10606
rect 2792 10560 2872 10588
rect 2792 8401 2820 10560
rect 2872 10542 2924 10548
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2778 8392 2834 8401
rect 2778 8327 2834 8336
rect 2780 4752 2832 4758
rect 2700 4712 2780 4740
rect 2780 4694 2832 4700
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 572 2984 624 2990
rect 572 2926 624 2932
rect 204 2848 256 2854
rect 204 2790 256 2796
rect 216 480 244 2790
rect 584 480 612 2926
rect 1032 2916 1084 2922
rect 1032 2858 1084 2864
rect 1044 480 1072 2858
rect 1412 480 1440 3470
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1872 480 1900 2994
rect 2332 480 2360 3130
rect 2700 480 2728 3334
rect 2976 1737 3004 10406
rect 3344 9722 3372 17598
rect 3421 17436 3717 17456
rect 3477 17434 3501 17436
rect 3557 17434 3581 17436
rect 3637 17434 3661 17436
rect 3499 17382 3501 17434
rect 3563 17382 3575 17434
rect 3637 17382 3639 17434
rect 3477 17380 3501 17382
rect 3557 17380 3581 17382
rect 3637 17380 3661 17382
rect 3421 17360 3717 17380
rect 3421 16348 3717 16368
rect 3477 16346 3501 16348
rect 3557 16346 3581 16348
rect 3637 16346 3661 16348
rect 3499 16294 3501 16346
rect 3563 16294 3575 16346
rect 3637 16294 3639 16346
rect 3477 16292 3501 16294
rect 3557 16292 3581 16294
rect 3637 16292 3661 16294
rect 3421 16272 3717 16292
rect 3421 15260 3717 15280
rect 3477 15258 3501 15260
rect 3557 15258 3581 15260
rect 3637 15258 3661 15260
rect 3499 15206 3501 15258
rect 3563 15206 3575 15258
rect 3637 15206 3639 15258
rect 3477 15204 3501 15206
rect 3557 15204 3581 15206
rect 3637 15204 3661 15206
rect 3421 15184 3717 15204
rect 3421 14172 3717 14192
rect 3477 14170 3501 14172
rect 3557 14170 3581 14172
rect 3637 14170 3661 14172
rect 3499 14118 3501 14170
rect 3563 14118 3575 14170
rect 3637 14118 3639 14170
rect 3477 14116 3501 14118
rect 3557 14116 3581 14118
rect 3637 14116 3661 14118
rect 3421 14096 3717 14116
rect 3421 13084 3717 13104
rect 3477 13082 3501 13084
rect 3557 13082 3581 13084
rect 3637 13082 3661 13084
rect 3499 13030 3501 13082
rect 3563 13030 3575 13082
rect 3637 13030 3639 13082
rect 3477 13028 3501 13030
rect 3557 13028 3581 13030
rect 3637 13028 3661 13030
rect 3421 13008 3717 13028
rect 3421 11996 3717 12016
rect 3477 11994 3501 11996
rect 3557 11994 3581 11996
rect 3637 11994 3661 11996
rect 3499 11942 3501 11994
rect 3563 11942 3575 11994
rect 3637 11942 3639 11994
rect 3477 11940 3501 11942
rect 3557 11940 3581 11942
rect 3637 11940 3661 11942
rect 3421 11920 3717 11940
rect 3421 10908 3717 10928
rect 3477 10906 3501 10908
rect 3557 10906 3581 10908
rect 3637 10906 3661 10908
rect 3499 10854 3501 10906
rect 3563 10854 3575 10906
rect 3637 10854 3639 10906
rect 3477 10852 3501 10854
rect 3557 10852 3581 10854
rect 3637 10852 3661 10854
rect 3421 10832 3717 10852
rect 3421 9820 3717 9840
rect 3477 9818 3501 9820
rect 3557 9818 3581 9820
rect 3637 9818 3661 9820
rect 3499 9766 3501 9818
rect 3563 9766 3575 9818
rect 3637 9766 3639 9818
rect 3477 9764 3501 9766
rect 3557 9764 3581 9766
rect 3637 9764 3661 9766
rect 3421 9744 3717 9764
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3421 8732 3717 8752
rect 3477 8730 3501 8732
rect 3557 8730 3581 8732
rect 3637 8730 3661 8732
rect 3499 8678 3501 8730
rect 3563 8678 3575 8730
rect 3637 8678 3639 8730
rect 3477 8676 3501 8678
rect 3557 8676 3581 8678
rect 3637 8676 3661 8678
rect 3421 8656 3717 8676
rect 3421 7644 3717 7664
rect 3477 7642 3501 7644
rect 3557 7642 3581 7644
rect 3637 7642 3661 7644
rect 3499 7590 3501 7642
rect 3563 7590 3575 7642
rect 3637 7590 3639 7642
rect 3477 7588 3501 7590
rect 3557 7588 3581 7590
rect 3637 7588 3661 7590
rect 3421 7568 3717 7588
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 3068 5001 3096 7210
rect 3421 6556 3717 6576
rect 3477 6554 3501 6556
rect 3557 6554 3581 6556
rect 3637 6554 3661 6556
rect 3499 6502 3501 6554
rect 3563 6502 3575 6554
rect 3637 6502 3639 6554
rect 3477 6500 3501 6502
rect 3557 6500 3581 6502
rect 3637 6500 3661 6502
rect 3421 6480 3717 6500
rect 3804 5642 3832 9658
rect 3896 7206 3924 19520
rect 3974 18320 4030 18329
rect 3974 18255 4030 18264
rect 3988 13938 4016 18255
rect 4356 15910 4384 19520
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4724 15366 4752 19520
rect 4896 17944 4948 17950
rect 4896 17886 4948 17892
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4264 13530 4292 13806
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4344 12368 4396 12374
rect 4344 12310 4396 12316
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 3421 5468 3717 5488
rect 3477 5466 3501 5468
rect 3557 5466 3581 5468
rect 3637 5466 3661 5468
rect 3499 5414 3501 5466
rect 3563 5414 3575 5466
rect 3637 5414 3639 5466
rect 3477 5412 3501 5414
rect 3557 5412 3581 5414
rect 3637 5412 3661 5414
rect 3421 5392 3717 5412
rect 4080 5166 4108 11562
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4264 10810 4292 11222
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4356 5778 4384 12310
rect 4908 9518 4936 17886
rect 5184 15994 5212 19520
rect 5552 16522 5580 19520
rect 6012 17082 6040 19520
rect 6012 17054 6316 17082
rect 5886 16892 6182 16912
rect 5942 16890 5966 16892
rect 6022 16890 6046 16892
rect 6102 16890 6126 16892
rect 5964 16838 5966 16890
rect 6028 16838 6040 16890
rect 6102 16838 6104 16890
rect 5942 16836 5966 16838
rect 6022 16836 6046 16838
rect 6102 16836 6126 16838
rect 5886 16816 6182 16836
rect 6288 16590 6316 17054
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 6380 16454 6408 19520
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6840 16182 6868 19520
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 5184 15966 5488 15994
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5000 12442 5028 13330
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3884 5024 3936 5030
rect 3054 4992 3110 5001
rect 3884 4966 3936 4972
rect 3054 4927 3110 4936
rect 3421 4380 3717 4400
rect 3477 4378 3501 4380
rect 3557 4378 3581 4380
rect 3637 4378 3661 4380
rect 3499 4326 3501 4378
rect 3563 4326 3575 4378
rect 3637 4326 3639 4378
rect 3477 4324 3501 4326
rect 3557 4324 3581 4326
rect 3637 4324 3661 4326
rect 3421 4304 3717 4324
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 2962 1728 3018 1737
rect 2962 1663 3018 1672
rect 3160 480 3188 4014
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3421 3292 3717 3312
rect 3477 3290 3501 3292
rect 3557 3290 3581 3292
rect 3637 3290 3661 3292
rect 3499 3238 3501 3290
rect 3563 3238 3575 3290
rect 3637 3238 3639 3290
rect 3477 3236 3501 3238
rect 3557 3236 3581 3238
rect 3637 3236 3661 3238
rect 3421 3216 3717 3236
rect 3421 2204 3717 2224
rect 3477 2202 3501 2204
rect 3557 2202 3581 2204
rect 3637 2202 3661 2204
rect 3499 2150 3501 2202
rect 3563 2150 3575 2202
rect 3637 2150 3639 2202
rect 3477 2148 3501 2150
rect 3557 2148 3581 2150
rect 3637 2148 3661 2150
rect 3421 2128 3717 2148
rect 3804 1986 3832 3878
rect 3896 2854 3924 4966
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3620 1958 3832 1986
rect 3620 480 3648 1958
rect 3976 604 4028 610
rect 3976 546 4028 552
rect 3988 480 4016 546
rect 4448 480 4476 5850
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4540 2922 4568 5510
rect 4528 2916 4580 2922
rect 4528 2858 4580 2864
rect 4816 480 4844 5646
rect 5276 5166 5304 7346
rect 5368 5658 5396 15846
rect 5460 5794 5488 15966
rect 5886 15804 6182 15824
rect 5942 15802 5966 15804
rect 6022 15802 6046 15804
rect 6102 15802 6126 15804
rect 5964 15750 5966 15802
rect 6028 15750 6040 15802
rect 6102 15750 6104 15802
rect 5942 15748 5966 15750
rect 6022 15748 6046 15750
rect 6102 15748 6126 15750
rect 5886 15728 6182 15748
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 5886 14716 6182 14736
rect 5942 14714 5966 14716
rect 6022 14714 6046 14716
rect 6102 14714 6126 14716
rect 5964 14662 5966 14714
rect 6028 14662 6040 14714
rect 6102 14662 6104 14714
rect 5942 14660 5966 14662
rect 6022 14660 6046 14662
rect 6102 14660 6126 14662
rect 5886 14640 6182 14660
rect 5886 13628 6182 13648
rect 5942 13626 5966 13628
rect 6022 13626 6046 13628
rect 6102 13626 6126 13628
rect 5964 13574 5966 13626
rect 6028 13574 6040 13626
rect 6102 13574 6104 13626
rect 5942 13572 5966 13574
rect 6022 13572 6046 13574
rect 6102 13572 6126 13574
rect 5886 13552 6182 13572
rect 5886 12540 6182 12560
rect 5942 12538 5966 12540
rect 6022 12538 6046 12540
rect 6102 12538 6126 12540
rect 5964 12486 5966 12538
rect 6028 12486 6040 12538
rect 6102 12486 6104 12538
rect 5942 12484 5966 12486
rect 6022 12484 6046 12486
rect 6102 12484 6126 12486
rect 5886 12464 6182 12484
rect 6288 12238 6316 15574
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6840 15162 6868 15302
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 5886 11452 6182 11472
rect 5942 11450 5966 11452
rect 6022 11450 6046 11452
rect 6102 11450 6126 11452
rect 5964 11398 5966 11450
rect 6028 11398 6040 11450
rect 6102 11398 6104 11450
rect 5942 11396 5966 11398
rect 6022 11396 6046 11398
rect 6102 11396 6126 11398
rect 5886 11376 6182 11396
rect 5886 10364 6182 10384
rect 5942 10362 5966 10364
rect 6022 10362 6046 10364
rect 6102 10362 6126 10364
rect 5964 10310 5966 10362
rect 6028 10310 6040 10362
rect 6102 10310 6104 10362
rect 5942 10308 5966 10310
rect 6022 10308 6046 10310
rect 6102 10308 6126 10310
rect 5886 10288 6182 10308
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 7342 5580 9862
rect 5886 9276 6182 9296
rect 5942 9274 5966 9276
rect 6022 9274 6046 9276
rect 6102 9274 6126 9276
rect 5964 9222 5966 9274
rect 6028 9222 6040 9274
rect 6102 9222 6104 9274
rect 5942 9220 5966 9222
rect 6022 9220 6046 9222
rect 6102 9220 6126 9222
rect 5886 9200 6182 9220
rect 5886 8188 6182 8208
rect 5942 8186 5966 8188
rect 6022 8186 6046 8188
rect 6102 8186 6126 8188
rect 5964 8134 5966 8186
rect 6028 8134 6040 8186
rect 6102 8134 6104 8186
rect 5942 8132 5966 8134
rect 6022 8132 6046 8134
rect 6102 8132 6126 8134
rect 5886 8112 6182 8132
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5886 7100 6182 7120
rect 5942 7098 5966 7100
rect 6022 7098 6046 7100
rect 6102 7098 6126 7100
rect 5964 7046 5966 7098
rect 6028 7046 6040 7098
rect 6102 7046 6104 7098
rect 5942 7044 5966 7046
rect 6022 7044 6046 7046
rect 6102 7044 6126 7046
rect 5886 7024 6182 7044
rect 5886 6012 6182 6032
rect 5942 6010 5966 6012
rect 6022 6010 6046 6012
rect 6102 6010 6126 6012
rect 5964 5958 5966 6010
rect 6028 5958 6040 6010
rect 6102 5958 6104 6010
rect 5942 5956 5966 5958
rect 6022 5956 6046 5958
rect 6102 5956 6126 5958
rect 5886 5936 6182 5956
rect 5460 5766 5580 5794
rect 5368 5630 5488 5658
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5000 2990 5028 4966
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5276 480 5304 3402
rect 5368 3058 5396 5510
rect 5460 5370 5488 5630
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5552 5250 5580 5766
rect 5460 5222 5580 5250
rect 5460 4758 5488 5222
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5644 3738 5672 4626
rect 5736 4282 5764 5102
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 5736 480 5764 3946
rect 5828 3534 5856 4966
rect 5886 4924 6182 4944
rect 5942 4922 5966 4924
rect 6022 4922 6046 4924
rect 6102 4922 6126 4924
rect 5964 4870 5966 4922
rect 6028 4870 6040 4922
rect 6102 4870 6104 4922
rect 5942 4868 5966 4870
rect 6022 4868 6046 4870
rect 6102 4868 6126 4870
rect 5886 4848 6182 4868
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 5886 3836 6182 3856
rect 5942 3834 5966 3836
rect 6022 3834 6046 3836
rect 6102 3834 6126 3836
rect 5964 3782 5966 3834
rect 6028 3782 6040 3834
rect 6102 3782 6104 3834
rect 5942 3780 5966 3782
rect 6022 3780 6046 3782
rect 6102 3780 6126 3782
rect 5886 3760 6182 3780
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 5886 2748 6182 2768
rect 5942 2746 5966 2748
rect 6022 2746 6046 2748
rect 6102 2746 6126 2748
rect 5964 2694 5966 2746
rect 6028 2694 6040 2746
rect 6102 2694 6104 2746
rect 5942 2692 5966 2694
rect 6022 2692 6046 2694
rect 6102 2692 6126 2694
rect 5886 2672 6182 2692
rect 6288 1850 6316 2994
rect 6104 1822 6316 1850
rect 6104 480 6132 1822
rect 6380 610 6408 4490
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6368 604 6420 610
rect 6368 546 6420 552
rect 6564 480 6592 4082
rect 6656 2922 6684 12174
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6748 11354 6776 11494
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6932 11286 6960 12106
rect 7116 11558 7144 15642
rect 7208 15366 7236 19520
rect 7668 16402 7696 19520
rect 7668 16374 7788 16402
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7300 15178 7328 16050
rect 7208 15150 7328 15178
rect 7208 11626 7236 15150
rect 7668 12714 7696 16186
rect 7760 15502 7788 16374
rect 8036 15722 8064 19520
rect 8496 17626 8524 19520
rect 8496 17598 8708 17626
rect 8352 17436 8648 17456
rect 8408 17434 8432 17436
rect 8488 17434 8512 17436
rect 8568 17434 8592 17436
rect 8430 17382 8432 17434
rect 8494 17382 8506 17434
rect 8568 17382 8570 17434
rect 8408 17380 8432 17382
rect 8488 17380 8512 17382
rect 8568 17380 8592 17382
rect 8352 17360 8648 17380
rect 8352 16348 8648 16368
rect 8408 16346 8432 16348
rect 8488 16346 8512 16348
rect 8568 16346 8592 16348
rect 8430 16294 8432 16346
rect 8494 16294 8506 16346
rect 8568 16294 8570 16346
rect 8408 16292 8432 16294
rect 8488 16292 8512 16294
rect 8568 16292 8592 16294
rect 8352 16272 8648 16292
rect 8680 16046 8708 17598
rect 8864 16114 8892 19520
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8668 16040 8720 16046
rect 9324 16028 9352 19520
rect 8668 15982 8720 15988
rect 8956 16000 9352 16028
rect 9588 16040 9640 16046
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 8036 15694 8156 15722
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7852 12782 7880 15506
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 7300 11218 7328 11630
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6748 9602 6776 9658
rect 7116 9654 7144 10066
rect 7104 9648 7156 9654
rect 6748 9574 6960 9602
rect 7104 9590 7156 9596
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6748 4486 6776 9454
rect 6932 5166 6960 9574
rect 7208 9518 7236 11018
rect 7300 10810 7328 11154
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7300 10130 7328 10746
rect 7392 10606 7420 12378
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7576 11218 7604 11698
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7668 10690 7696 12650
rect 7576 10662 7696 10690
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7196 6180 7248 6186
rect 7196 6122 7248 6128
rect 7208 5778 7236 6122
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7392 5778 7420 6054
rect 7576 5846 7604 10662
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7668 10198 7696 10542
rect 7656 10192 7708 10198
rect 7708 10140 7788 10146
rect 7656 10134 7788 10140
rect 7668 10118 7788 10134
rect 7760 9586 7788 10118
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7852 7562 7880 12718
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7944 9926 7972 11562
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 8036 9722 8064 15506
rect 8128 15434 8156 15694
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 8128 12850 8156 13942
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8128 12170 8156 12786
rect 8220 12374 8248 15914
rect 8352 15260 8648 15280
rect 8408 15258 8432 15260
rect 8488 15258 8512 15260
rect 8568 15258 8592 15260
rect 8430 15206 8432 15258
rect 8494 15206 8506 15258
rect 8568 15206 8570 15258
rect 8408 15204 8432 15206
rect 8488 15204 8512 15206
rect 8568 15204 8592 15206
rect 8352 15184 8648 15204
rect 8352 14172 8648 14192
rect 8408 14170 8432 14172
rect 8488 14170 8512 14172
rect 8568 14170 8592 14172
rect 8430 14118 8432 14170
rect 8494 14118 8506 14170
rect 8568 14118 8570 14170
rect 8408 14116 8432 14118
rect 8488 14116 8512 14118
rect 8568 14116 8592 14118
rect 8352 14096 8648 14116
rect 8352 13084 8648 13104
rect 8408 13082 8432 13084
rect 8488 13082 8512 13084
rect 8568 13082 8592 13084
rect 8430 13030 8432 13082
rect 8494 13030 8506 13082
rect 8568 13030 8570 13082
rect 8408 13028 8432 13030
rect 8488 13028 8512 13030
rect 8568 13028 8592 13030
rect 8352 13008 8648 13028
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 8128 11898 8156 12106
rect 8352 11996 8648 12016
rect 8408 11994 8432 11996
rect 8488 11994 8512 11996
rect 8568 11994 8592 11996
rect 8430 11942 8432 11994
rect 8494 11942 8506 11994
rect 8568 11942 8570 11994
rect 8408 11940 8432 11942
rect 8488 11940 8512 11942
rect 8568 11940 8592 11942
rect 8352 11920 8648 11940
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7852 7534 7972 7562
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 7024 5114 7052 5510
rect 7024 5086 7144 5114
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6840 3466 6868 4762
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6932 3602 6960 4626
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 7024 3194 7052 4966
rect 7116 4078 7144 5086
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 7484 2666 7512 5578
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7576 3398 7604 4966
rect 7668 4758 7696 4966
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7852 4486 7880 7142
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7392 2638 7512 2666
rect 7012 2100 7064 2106
rect 7012 2042 7064 2048
rect 7024 480 7052 2042
rect 7392 480 7420 2638
rect 7852 480 7880 3606
rect 7944 3466 7972 7534
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 8036 2106 8064 5578
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8128 2990 8156 5034
rect 8220 3398 8248 11494
rect 8352 10908 8648 10928
rect 8408 10906 8432 10908
rect 8488 10906 8512 10908
rect 8568 10906 8592 10908
rect 8430 10854 8432 10906
rect 8494 10854 8506 10906
rect 8568 10854 8570 10906
rect 8408 10852 8432 10854
rect 8488 10852 8512 10854
rect 8568 10852 8592 10854
rect 8352 10832 8648 10852
rect 8352 9820 8648 9840
rect 8408 9818 8432 9820
rect 8488 9818 8512 9820
rect 8568 9818 8592 9820
rect 8430 9766 8432 9818
rect 8494 9766 8506 9818
rect 8568 9766 8570 9818
rect 8408 9764 8432 9766
rect 8488 9764 8512 9766
rect 8568 9764 8592 9766
rect 8352 9744 8648 9764
rect 8680 9586 8708 12854
rect 8956 12458 8984 16000
rect 9588 15982 9640 15988
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9140 12646 9168 13262
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 8864 12442 8984 12458
rect 8852 12436 8984 12442
rect 8904 12430 8984 12436
rect 9036 12436 9088 12442
rect 8852 12378 8904 12384
rect 9036 12378 9088 12384
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8772 10538 8800 10950
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8760 10532 8812 10538
rect 8760 10474 8812 10480
rect 8772 9586 8800 10474
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8352 8732 8648 8752
rect 8408 8730 8432 8732
rect 8488 8730 8512 8732
rect 8568 8730 8592 8732
rect 8430 8678 8432 8730
rect 8494 8678 8506 8730
rect 8568 8678 8570 8730
rect 8408 8676 8432 8678
rect 8488 8676 8512 8678
rect 8568 8676 8592 8678
rect 8352 8656 8648 8676
rect 8352 7644 8648 7664
rect 8408 7642 8432 7644
rect 8488 7642 8512 7644
rect 8568 7642 8592 7644
rect 8430 7590 8432 7642
rect 8494 7590 8506 7642
rect 8568 7590 8570 7642
rect 8408 7588 8432 7590
rect 8488 7588 8512 7590
rect 8568 7588 8592 7590
rect 8352 7568 8648 7588
rect 8352 6556 8648 6576
rect 8408 6554 8432 6556
rect 8488 6554 8512 6556
rect 8568 6554 8592 6556
rect 8430 6502 8432 6554
rect 8494 6502 8506 6554
rect 8568 6502 8570 6554
rect 8408 6500 8432 6502
rect 8488 6500 8512 6502
rect 8568 6500 8592 6502
rect 8352 6480 8648 6500
rect 8352 5468 8648 5488
rect 8408 5466 8432 5468
rect 8488 5466 8512 5468
rect 8568 5466 8592 5468
rect 8430 5414 8432 5466
rect 8494 5414 8506 5466
rect 8568 5414 8570 5466
rect 8408 5412 8432 5414
rect 8488 5412 8512 5414
rect 8568 5412 8592 5414
rect 8352 5392 8648 5412
rect 8300 4616 8352 4622
rect 8352 4564 8708 4570
rect 8300 4558 8708 4564
rect 8312 4542 8708 4558
rect 8352 4380 8648 4400
rect 8408 4378 8432 4380
rect 8488 4378 8512 4380
rect 8568 4378 8592 4380
rect 8430 4326 8432 4378
rect 8494 4326 8506 4378
rect 8568 4326 8570 4378
rect 8408 4324 8432 4326
rect 8488 4324 8512 4326
rect 8568 4324 8592 4326
rect 8352 4304 8648 4324
rect 8680 3534 8708 4542
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8772 3398 8800 9318
rect 8864 5778 8892 10746
rect 9048 7410 9076 12378
rect 9140 11898 9168 12582
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9232 10554 9260 15574
rect 9140 10526 9260 10554
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9140 5778 9168 10526
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9232 10266 9260 10406
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9324 4690 9352 15846
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9416 15162 9444 15302
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 9416 9382 9444 14826
rect 9508 10810 9536 15642
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9600 8650 9628 15982
rect 9692 15978 9720 19520
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 9772 16176 9824 16182
rect 9772 16118 9824 16124
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9692 10606 9720 10950
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9508 8622 9628 8650
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9416 4826 9444 5102
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9508 4214 9536 8622
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9588 4752 9640 4758
rect 9588 4694 9640 4700
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9600 3738 9628 4694
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8352 3292 8648 3312
rect 8408 3290 8432 3292
rect 8488 3290 8512 3292
rect 8568 3290 8592 3292
rect 8430 3238 8432 3290
rect 8494 3238 8506 3290
rect 8568 3238 8570 3290
rect 8408 3236 8432 3238
rect 8488 3236 8512 3238
rect 8568 3236 8592 3238
rect 8352 3216 8648 3236
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8024 2100 8076 2106
rect 8024 2042 8076 2048
rect 8220 480 8248 3062
rect 8352 2204 8648 2224
rect 8408 2202 8432 2204
rect 8488 2202 8512 2204
rect 8568 2202 8592 2204
rect 8430 2150 8432 2202
rect 8494 2150 8506 2202
rect 8568 2150 8570 2202
rect 8408 2148 8432 2150
rect 8488 2148 8512 2150
rect 8568 2148 8592 2150
rect 8352 2128 8648 2148
rect 8680 480 8708 3334
rect 9140 480 9168 3674
rect 9692 3058 9720 5510
rect 9784 5030 9812 16118
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9876 15638 9904 15846
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9968 15450 9996 16458
rect 9876 15422 9996 15450
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9876 4826 9904 15422
rect 10152 14634 10180 19520
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 9968 14606 10180 14634
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9968 4282 9996 14606
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10060 10266 10088 11154
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10152 5778 10180 11290
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10244 6186 10272 10746
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 10336 5370 10364 16390
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10152 5250 10180 5306
rect 10428 5302 10456 16526
rect 10520 16250 10548 19520
rect 10980 17082 11008 19520
rect 10612 17054 11008 17082
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10416 5296 10468 5302
rect 10152 5222 10272 5250
rect 10416 5238 10468 5244
rect 10244 5166 10272 5222
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10060 4434 10088 5102
rect 10060 4406 10272 4434
rect 10244 4282 10272 4406
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 9770 4176 9826 4185
rect 9770 4111 9826 4120
rect 9784 4078 9812 4111
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9508 480 9536 2858
rect 9968 480 9996 3538
rect 10336 3058 10364 5170
rect 10520 5166 10548 16050
rect 10612 15570 10640 17054
rect 10817 16892 11113 16912
rect 10873 16890 10897 16892
rect 10953 16890 10977 16892
rect 11033 16890 11057 16892
rect 10895 16838 10897 16890
rect 10959 16838 10971 16890
rect 11033 16838 11035 16890
rect 10873 16836 10897 16838
rect 10953 16836 10977 16838
rect 11033 16836 11057 16838
rect 10817 16816 11113 16836
rect 11348 16114 11376 19520
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11808 16046 11836 19520
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10612 10690 10640 14894
rect 10704 10810 10732 15982
rect 10817 15804 11113 15824
rect 10873 15802 10897 15804
rect 10953 15802 10977 15804
rect 11033 15802 11057 15804
rect 10895 15750 10897 15802
rect 10959 15750 10971 15802
rect 11033 15750 11035 15802
rect 10873 15748 10897 15750
rect 10953 15748 10977 15750
rect 11033 15748 11057 15750
rect 10817 15728 11113 15748
rect 12176 15552 12204 19520
rect 12084 15524 12204 15552
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 10817 14716 11113 14736
rect 10873 14714 10897 14716
rect 10953 14714 10977 14716
rect 11033 14714 11057 14716
rect 10895 14662 10897 14714
rect 10959 14662 10971 14714
rect 11033 14662 11035 14714
rect 10873 14660 10897 14662
rect 10953 14660 10977 14662
rect 11033 14660 11057 14662
rect 10817 14640 11113 14660
rect 10817 13628 11113 13648
rect 10873 13626 10897 13628
rect 10953 13626 10977 13628
rect 11033 13626 11057 13628
rect 10895 13574 10897 13626
rect 10959 13574 10971 13626
rect 11033 13574 11035 13626
rect 10873 13572 10897 13574
rect 10953 13572 10977 13574
rect 11033 13572 11057 13574
rect 10817 13552 11113 13572
rect 10817 12540 11113 12560
rect 10873 12538 10897 12540
rect 10953 12538 10977 12540
rect 11033 12538 11057 12540
rect 10895 12486 10897 12538
rect 10959 12486 10971 12538
rect 11033 12486 11035 12538
rect 10873 12484 10897 12486
rect 10953 12484 10977 12486
rect 11033 12484 11057 12486
rect 10817 12464 11113 12484
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 10817 11452 11113 11472
rect 10873 11450 10897 11452
rect 10953 11450 10977 11452
rect 11033 11450 11057 11452
rect 10895 11398 10897 11450
rect 10959 11398 10971 11450
rect 11033 11398 11035 11450
rect 10873 11396 10897 11398
rect 10953 11396 10977 11398
rect 11033 11396 11057 11398
rect 10817 11376 11113 11396
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10612 10662 10732 10690
rect 10704 10606 10732 10662
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10600 5092 10652 5098
rect 10600 5034 10652 5040
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10428 480 10456 3402
rect 10612 3398 10640 5034
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10520 2922 10548 3334
rect 10704 3194 10732 10542
rect 10817 10364 11113 10384
rect 10873 10362 10897 10364
rect 10953 10362 10977 10364
rect 11033 10362 11057 10364
rect 10895 10310 10897 10362
rect 10959 10310 10971 10362
rect 11033 10310 11035 10362
rect 10873 10308 10897 10310
rect 10953 10308 10977 10310
rect 11033 10308 11057 10310
rect 10817 10288 11113 10308
rect 10817 9276 11113 9296
rect 10873 9274 10897 9276
rect 10953 9274 10977 9276
rect 11033 9274 11057 9276
rect 10895 9222 10897 9274
rect 10959 9222 10971 9274
rect 11033 9222 11035 9274
rect 10873 9220 10897 9222
rect 10953 9220 10977 9222
rect 11033 9220 11057 9222
rect 10817 9200 11113 9220
rect 11164 8974 11192 12242
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11256 9602 11284 9658
rect 11256 9574 11376 9602
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 10817 8188 11113 8208
rect 10873 8186 10897 8188
rect 10953 8186 10977 8188
rect 11033 8186 11057 8188
rect 10895 8134 10897 8186
rect 10959 8134 10971 8186
rect 11033 8134 11035 8186
rect 10873 8132 10897 8134
rect 10953 8132 10977 8134
rect 11033 8132 11057 8134
rect 10817 8112 11113 8132
rect 10817 7100 11113 7120
rect 10873 7098 10897 7100
rect 10953 7098 10977 7100
rect 11033 7098 11057 7100
rect 10895 7046 10897 7098
rect 10959 7046 10971 7098
rect 11033 7046 11035 7098
rect 10873 7044 10897 7046
rect 10953 7044 10977 7046
rect 11033 7044 11057 7046
rect 10817 7024 11113 7044
rect 10817 6012 11113 6032
rect 10873 6010 10897 6012
rect 10953 6010 10977 6012
rect 11033 6010 11057 6012
rect 10895 5958 10897 6010
rect 10959 5958 10971 6010
rect 11033 5958 11035 6010
rect 10873 5956 10897 5958
rect 10953 5956 10977 5958
rect 11033 5956 11057 5958
rect 10817 5936 11113 5956
rect 10817 4924 11113 4944
rect 10873 4922 10897 4924
rect 10953 4922 10977 4924
rect 11033 4922 11057 4924
rect 10895 4870 10897 4922
rect 10959 4870 10971 4922
rect 11033 4870 11035 4922
rect 10873 4868 10897 4870
rect 10953 4868 10977 4870
rect 11033 4868 11057 4870
rect 10817 4848 11113 4868
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10888 4146 10916 4422
rect 11348 4185 11376 9574
rect 11440 5370 11468 15438
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11334 4176 11390 4185
rect 10876 4140 10928 4146
rect 11334 4111 11390 4120
rect 10876 4082 10928 4088
rect 10817 3836 11113 3856
rect 10873 3834 10897 3836
rect 10953 3834 10977 3836
rect 11033 3834 11057 3836
rect 10895 3782 10897 3834
rect 10959 3782 10971 3834
rect 11033 3782 11035 3834
rect 10873 3780 10897 3782
rect 10953 3780 10977 3782
rect 11033 3780 11057 3782
rect 10817 3760 11113 3780
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10692 2984 10744 2990
rect 10692 2926 10744 2932
rect 10508 2916 10560 2922
rect 10508 2858 10560 2864
rect 10704 2530 10732 2926
rect 10817 2748 11113 2768
rect 10873 2746 10897 2748
rect 10953 2746 10977 2748
rect 11033 2746 11057 2748
rect 10895 2694 10897 2746
rect 10959 2694 10971 2746
rect 11033 2694 11035 2746
rect 10873 2692 10897 2694
rect 10953 2692 10977 2694
rect 11033 2692 11057 2694
rect 10817 2672 11113 2692
rect 10704 2502 10824 2530
rect 10796 480 10824 2502
rect 11256 480 11284 3470
rect 11624 480 11652 6054
rect 11992 4758 12020 15438
rect 12084 9722 12112 15524
rect 12164 15428 12216 15434
rect 12164 15370 12216 15376
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 12176 5370 12204 15370
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12452 7449 12480 8978
rect 12438 7440 12494 7449
rect 12438 7375 12494 7384
rect 12636 5794 12664 19520
rect 13004 15706 13032 19520
rect 13464 17626 13492 19520
rect 13188 17598 13492 17626
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 12992 15428 13044 15434
rect 12992 15370 13044 15376
rect 12452 5766 12664 5794
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 11980 4752 12032 4758
rect 11980 4694 12032 4700
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 11980 3732 12032 3738
rect 11980 3674 12032 3680
rect 11992 2394 12020 3674
rect 12084 3670 12112 4422
rect 12176 4214 12204 4694
rect 12452 4554 12480 5766
rect 13004 5166 13032 15370
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12452 2666 12480 2994
rect 12544 2854 12572 4966
rect 12636 4758 12664 4966
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 13096 4690 13124 15982
rect 13188 15910 13216 17598
rect 13726 17504 13782 17513
rect 13282 17436 13578 17456
rect 13726 17439 13782 17448
rect 13338 17434 13362 17436
rect 13418 17434 13442 17436
rect 13498 17434 13522 17436
rect 13360 17382 13362 17434
rect 13424 17382 13436 17434
rect 13498 17382 13500 17434
rect 13338 17380 13362 17382
rect 13418 17380 13442 17382
rect 13498 17380 13522 17382
rect 13282 17360 13578 17380
rect 13282 16348 13578 16368
rect 13338 16346 13362 16348
rect 13418 16346 13442 16348
rect 13498 16346 13522 16348
rect 13360 16294 13362 16346
rect 13424 16294 13436 16346
rect 13498 16294 13500 16346
rect 13338 16292 13362 16294
rect 13418 16292 13442 16294
rect 13498 16292 13522 16294
rect 13282 16272 13578 16292
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13282 15260 13578 15280
rect 13338 15258 13362 15260
rect 13418 15258 13442 15260
rect 13498 15258 13522 15260
rect 13360 15206 13362 15258
rect 13424 15206 13436 15258
rect 13498 15206 13500 15258
rect 13338 15204 13362 15206
rect 13418 15204 13442 15206
rect 13498 15204 13522 15206
rect 13282 15184 13578 15204
rect 13282 14172 13578 14192
rect 13338 14170 13362 14172
rect 13418 14170 13442 14172
rect 13498 14170 13522 14172
rect 13360 14118 13362 14170
rect 13424 14118 13436 14170
rect 13498 14118 13500 14170
rect 13338 14116 13362 14118
rect 13418 14116 13442 14118
rect 13498 14116 13522 14118
rect 13282 14096 13578 14116
rect 13740 14074 13768 17439
rect 13832 15978 13860 19520
rect 14016 19502 14320 19520
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13282 13084 13578 13104
rect 13338 13082 13362 13084
rect 13418 13082 13442 13084
rect 13498 13082 13522 13084
rect 13360 13030 13362 13082
rect 13424 13030 13436 13082
rect 13498 13030 13500 13082
rect 13338 13028 13362 13030
rect 13418 13028 13442 13030
rect 13498 13028 13522 13030
rect 13282 13008 13578 13028
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13464 12481 13492 12582
rect 13450 12472 13506 12481
rect 13450 12407 13506 12416
rect 13282 11996 13578 12016
rect 13338 11994 13362 11996
rect 13418 11994 13442 11996
rect 13498 11994 13522 11996
rect 13360 11942 13362 11994
rect 13424 11942 13436 11994
rect 13498 11942 13500 11994
rect 13338 11940 13362 11942
rect 13418 11940 13442 11942
rect 13498 11940 13522 11942
rect 13282 11920 13578 11940
rect 13648 11286 13676 13806
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 13282 10908 13578 10928
rect 13338 10906 13362 10908
rect 13418 10906 13442 10908
rect 13498 10906 13522 10908
rect 13360 10854 13362 10906
rect 13424 10854 13436 10906
rect 13498 10854 13500 10906
rect 13338 10852 13362 10854
rect 13418 10852 13442 10854
rect 13498 10852 13522 10854
rect 13282 10832 13578 10852
rect 13282 9820 13578 9840
rect 13338 9818 13362 9820
rect 13418 9818 13442 9820
rect 13498 9818 13522 9820
rect 13360 9766 13362 9818
rect 13424 9766 13436 9818
rect 13498 9766 13500 9818
rect 13338 9764 13362 9766
rect 13418 9764 13442 9766
rect 13498 9764 13522 9766
rect 13282 9744 13578 9764
rect 13282 8732 13578 8752
rect 13338 8730 13362 8732
rect 13418 8730 13442 8732
rect 13498 8730 13522 8732
rect 13360 8678 13362 8730
rect 13424 8678 13436 8730
rect 13498 8678 13500 8730
rect 13338 8676 13362 8678
rect 13418 8676 13442 8678
rect 13498 8676 13522 8678
rect 13282 8656 13578 8676
rect 13282 7644 13578 7664
rect 13338 7642 13362 7644
rect 13418 7642 13442 7644
rect 13498 7642 13522 7644
rect 13360 7590 13362 7642
rect 13424 7590 13436 7642
rect 13498 7590 13500 7642
rect 13338 7588 13362 7590
rect 13418 7588 13442 7590
rect 13498 7588 13522 7590
rect 13282 7568 13578 7588
rect 13282 6556 13578 6576
rect 13338 6554 13362 6556
rect 13418 6554 13442 6556
rect 13498 6554 13522 6556
rect 13360 6502 13362 6554
rect 13424 6502 13436 6554
rect 13498 6502 13500 6554
rect 13338 6500 13362 6502
rect 13418 6500 13442 6502
rect 13498 6500 13522 6502
rect 13282 6480 13578 6500
rect 13282 5468 13578 5488
rect 13338 5466 13362 5468
rect 13418 5466 13442 5468
rect 13498 5466 13522 5468
rect 13360 5414 13362 5466
rect 13424 5414 13436 5466
rect 13498 5414 13500 5466
rect 13338 5412 13362 5414
rect 13418 5412 13442 5414
rect 13498 5412 13522 5414
rect 13282 5392 13578 5412
rect 13176 5024 13228 5030
rect 13176 4966 13228 4972
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 12452 2638 12572 2666
rect 11992 2366 12112 2394
rect 12084 480 12112 2366
rect 12544 480 12572 2638
rect 12912 480 12940 2858
rect 13096 1986 13124 3334
rect 13188 3126 13216 4966
rect 13282 4380 13578 4400
rect 13338 4378 13362 4380
rect 13418 4378 13442 4380
rect 13498 4378 13522 4380
rect 13360 4326 13362 4378
rect 13424 4326 13436 4378
rect 13498 4326 13500 4378
rect 13338 4324 13362 4326
rect 13418 4324 13442 4326
rect 13498 4324 13522 4326
rect 13282 4304 13578 4324
rect 13282 3292 13578 3312
rect 13338 3290 13362 3292
rect 13418 3290 13442 3292
rect 13498 3290 13522 3292
rect 13360 3238 13362 3290
rect 13424 3238 13436 3290
rect 13498 3238 13500 3290
rect 13338 3236 13362 3238
rect 13418 3236 13442 3238
rect 13498 3236 13522 3238
rect 13282 3216 13578 3236
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13648 2553 13676 11222
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13924 5846 13952 7142
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13740 2802 13768 4558
rect 14016 4078 14044 19502
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14476 5778 14504 15438
rect 14660 7206 14688 19520
rect 15120 15570 15148 19520
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 15488 11354 15516 19520
rect 15948 15502 15976 19520
rect 16316 16046 16344 19520
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 16776 15434 16804 19520
rect 16764 15428 16816 15434
rect 16764 15370 16816 15376
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 15936 5296 15988 5302
rect 15936 5238 15988 5244
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13740 2774 13860 2802
rect 13634 2544 13690 2553
rect 13634 2479 13690 2488
rect 13282 2204 13578 2224
rect 13338 2202 13362 2204
rect 13418 2202 13442 2204
rect 13498 2202 13522 2204
rect 13360 2150 13362 2202
rect 13424 2150 13436 2202
rect 13498 2150 13500 2202
rect 13338 2148 13362 2150
rect 13418 2148 13442 2150
rect 13498 2148 13522 2150
rect 13282 2128 13578 2148
rect 13096 1958 13400 1986
rect 13372 480 13400 1958
rect 13832 480 13860 2774
rect 14200 480 14228 4762
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14660 480 14688 4082
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15028 480 15056 2790
rect 15488 480 15516 3130
rect 15948 480 15976 5238
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16316 480 16344 5170
rect 16764 5092 16816 5098
rect 16764 5034 16816 5040
rect 16776 480 16804 5034
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1398 0 1454 480
rect 1858 0 1914 480
rect 2318 0 2374 480
rect 2686 0 2742 480
rect 3146 0 3202 480
rect 3606 0 3662 480
rect 3974 0 4030 480
rect 4434 0 4490 480
rect 4802 0 4858 480
rect 5262 0 5318 480
rect 5722 0 5778 480
rect 6090 0 6146 480
rect 6550 0 6606 480
rect 7010 0 7066 480
rect 7378 0 7434 480
rect 7838 0 7894 480
rect 8206 0 8262 480
rect 8666 0 8722 480
rect 9126 0 9182 480
rect 9494 0 9550 480
rect 9954 0 10010 480
rect 10414 0 10470 480
rect 10782 0 10838 480
rect 11242 0 11298 480
rect 11610 0 11666 480
rect 12070 0 12126 480
rect 12530 0 12586 480
rect 12898 0 12954 480
rect 13358 0 13414 480
rect 13818 0 13874 480
rect 14186 0 14242 480
rect 14646 0 14702 480
rect 15014 0 15070 480
rect 15474 0 15530 480
rect 15934 0 15990 480
rect 16302 0 16358 480
rect 16762 0 16818 480
<< via2 >>
rect 2778 15000 2834 15056
rect 3146 11600 3202 11656
rect 2778 8336 2834 8392
rect 3421 17434 3477 17436
rect 3501 17434 3557 17436
rect 3581 17434 3637 17436
rect 3661 17434 3717 17436
rect 3421 17382 3447 17434
rect 3447 17382 3477 17434
rect 3501 17382 3511 17434
rect 3511 17382 3557 17434
rect 3581 17382 3627 17434
rect 3627 17382 3637 17434
rect 3661 17382 3691 17434
rect 3691 17382 3717 17434
rect 3421 17380 3477 17382
rect 3501 17380 3557 17382
rect 3581 17380 3637 17382
rect 3661 17380 3717 17382
rect 3421 16346 3477 16348
rect 3501 16346 3557 16348
rect 3581 16346 3637 16348
rect 3661 16346 3717 16348
rect 3421 16294 3447 16346
rect 3447 16294 3477 16346
rect 3501 16294 3511 16346
rect 3511 16294 3557 16346
rect 3581 16294 3627 16346
rect 3627 16294 3637 16346
rect 3661 16294 3691 16346
rect 3691 16294 3717 16346
rect 3421 16292 3477 16294
rect 3501 16292 3557 16294
rect 3581 16292 3637 16294
rect 3661 16292 3717 16294
rect 3421 15258 3477 15260
rect 3501 15258 3557 15260
rect 3581 15258 3637 15260
rect 3661 15258 3717 15260
rect 3421 15206 3447 15258
rect 3447 15206 3477 15258
rect 3501 15206 3511 15258
rect 3511 15206 3557 15258
rect 3581 15206 3627 15258
rect 3627 15206 3637 15258
rect 3661 15206 3691 15258
rect 3691 15206 3717 15258
rect 3421 15204 3477 15206
rect 3501 15204 3557 15206
rect 3581 15204 3637 15206
rect 3661 15204 3717 15206
rect 3421 14170 3477 14172
rect 3501 14170 3557 14172
rect 3581 14170 3637 14172
rect 3661 14170 3717 14172
rect 3421 14118 3447 14170
rect 3447 14118 3477 14170
rect 3501 14118 3511 14170
rect 3511 14118 3557 14170
rect 3581 14118 3627 14170
rect 3627 14118 3637 14170
rect 3661 14118 3691 14170
rect 3691 14118 3717 14170
rect 3421 14116 3477 14118
rect 3501 14116 3557 14118
rect 3581 14116 3637 14118
rect 3661 14116 3717 14118
rect 3421 13082 3477 13084
rect 3501 13082 3557 13084
rect 3581 13082 3637 13084
rect 3661 13082 3717 13084
rect 3421 13030 3447 13082
rect 3447 13030 3477 13082
rect 3501 13030 3511 13082
rect 3511 13030 3557 13082
rect 3581 13030 3627 13082
rect 3627 13030 3637 13082
rect 3661 13030 3691 13082
rect 3691 13030 3717 13082
rect 3421 13028 3477 13030
rect 3501 13028 3557 13030
rect 3581 13028 3637 13030
rect 3661 13028 3717 13030
rect 3421 11994 3477 11996
rect 3501 11994 3557 11996
rect 3581 11994 3637 11996
rect 3661 11994 3717 11996
rect 3421 11942 3447 11994
rect 3447 11942 3477 11994
rect 3501 11942 3511 11994
rect 3511 11942 3557 11994
rect 3581 11942 3627 11994
rect 3627 11942 3637 11994
rect 3661 11942 3691 11994
rect 3691 11942 3717 11994
rect 3421 11940 3477 11942
rect 3501 11940 3557 11942
rect 3581 11940 3637 11942
rect 3661 11940 3717 11942
rect 3421 10906 3477 10908
rect 3501 10906 3557 10908
rect 3581 10906 3637 10908
rect 3661 10906 3717 10908
rect 3421 10854 3447 10906
rect 3447 10854 3477 10906
rect 3501 10854 3511 10906
rect 3511 10854 3557 10906
rect 3581 10854 3627 10906
rect 3627 10854 3637 10906
rect 3661 10854 3691 10906
rect 3691 10854 3717 10906
rect 3421 10852 3477 10854
rect 3501 10852 3557 10854
rect 3581 10852 3637 10854
rect 3661 10852 3717 10854
rect 3421 9818 3477 9820
rect 3501 9818 3557 9820
rect 3581 9818 3637 9820
rect 3661 9818 3717 9820
rect 3421 9766 3447 9818
rect 3447 9766 3477 9818
rect 3501 9766 3511 9818
rect 3511 9766 3557 9818
rect 3581 9766 3627 9818
rect 3627 9766 3637 9818
rect 3661 9766 3691 9818
rect 3691 9766 3717 9818
rect 3421 9764 3477 9766
rect 3501 9764 3557 9766
rect 3581 9764 3637 9766
rect 3661 9764 3717 9766
rect 3421 8730 3477 8732
rect 3501 8730 3557 8732
rect 3581 8730 3637 8732
rect 3661 8730 3717 8732
rect 3421 8678 3447 8730
rect 3447 8678 3477 8730
rect 3501 8678 3511 8730
rect 3511 8678 3557 8730
rect 3581 8678 3627 8730
rect 3627 8678 3637 8730
rect 3661 8678 3691 8730
rect 3691 8678 3717 8730
rect 3421 8676 3477 8678
rect 3501 8676 3557 8678
rect 3581 8676 3637 8678
rect 3661 8676 3717 8678
rect 3421 7642 3477 7644
rect 3501 7642 3557 7644
rect 3581 7642 3637 7644
rect 3661 7642 3717 7644
rect 3421 7590 3447 7642
rect 3447 7590 3477 7642
rect 3501 7590 3511 7642
rect 3511 7590 3557 7642
rect 3581 7590 3627 7642
rect 3627 7590 3637 7642
rect 3661 7590 3691 7642
rect 3691 7590 3717 7642
rect 3421 7588 3477 7590
rect 3501 7588 3557 7590
rect 3581 7588 3637 7590
rect 3661 7588 3717 7590
rect 3421 6554 3477 6556
rect 3501 6554 3557 6556
rect 3581 6554 3637 6556
rect 3661 6554 3717 6556
rect 3421 6502 3447 6554
rect 3447 6502 3477 6554
rect 3501 6502 3511 6554
rect 3511 6502 3557 6554
rect 3581 6502 3627 6554
rect 3627 6502 3637 6554
rect 3661 6502 3691 6554
rect 3691 6502 3717 6554
rect 3421 6500 3477 6502
rect 3501 6500 3557 6502
rect 3581 6500 3637 6502
rect 3661 6500 3717 6502
rect 3974 18264 4030 18320
rect 3421 5466 3477 5468
rect 3501 5466 3557 5468
rect 3581 5466 3637 5468
rect 3661 5466 3717 5468
rect 3421 5414 3447 5466
rect 3447 5414 3477 5466
rect 3501 5414 3511 5466
rect 3511 5414 3557 5466
rect 3581 5414 3627 5466
rect 3627 5414 3637 5466
rect 3661 5414 3691 5466
rect 3691 5414 3717 5466
rect 3421 5412 3477 5414
rect 3501 5412 3557 5414
rect 3581 5412 3637 5414
rect 3661 5412 3717 5414
rect 5886 16890 5942 16892
rect 5966 16890 6022 16892
rect 6046 16890 6102 16892
rect 6126 16890 6182 16892
rect 5886 16838 5912 16890
rect 5912 16838 5942 16890
rect 5966 16838 5976 16890
rect 5976 16838 6022 16890
rect 6046 16838 6092 16890
rect 6092 16838 6102 16890
rect 6126 16838 6156 16890
rect 6156 16838 6182 16890
rect 5886 16836 5942 16838
rect 5966 16836 6022 16838
rect 6046 16836 6102 16838
rect 6126 16836 6182 16838
rect 3054 4936 3110 4992
rect 3421 4378 3477 4380
rect 3501 4378 3557 4380
rect 3581 4378 3637 4380
rect 3661 4378 3717 4380
rect 3421 4326 3447 4378
rect 3447 4326 3477 4378
rect 3501 4326 3511 4378
rect 3511 4326 3557 4378
rect 3581 4326 3627 4378
rect 3627 4326 3637 4378
rect 3661 4326 3691 4378
rect 3691 4326 3717 4378
rect 3421 4324 3477 4326
rect 3501 4324 3557 4326
rect 3581 4324 3637 4326
rect 3661 4324 3717 4326
rect 2962 1672 3018 1728
rect 3421 3290 3477 3292
rect 3501 3290 3557 3292
rect 3581 3290 3637 3292
rect 3661 3290 3717 3292
rect 3421 3238 3447 3290
rect 3447 3238 3477 3290
rect 3501 3238 3511 3290
rect 3511 3238 3557 3290
rect 3581 3238 3627 3290
rect 3627 3238 3637 3290
rect 3661 3238 3691 3290
rect 3691 3238 3717 3290
rect 3421 3236 3477 3238
rect 3501 3236 3557 3238
rect 3581 3236 3637 3238
rect 3661 3236 3717 3238
rect 3421 2202 3477 2204
rect 3501 2202 3557 2204
rect 3581 2202 3637 2204
rect 3661 2202 3717 2204
rect 3421 2150 3447 2202
rect 3447 2150 3477 2202
rect 3501 2150 3511 2202
rect 3511 2150 3557 2202
rect 3581 2150 3627 2202
rect 3627 2150 3637 2202
rect 3661 2150 3691 2202
rect 3691 2150 3717 2202
rect 3421 2148 3477 2150
rect 3501 2148 3557 2150
rect 3581 2148 3637 2150
rect 3661 2148 3717 2150
rect 5886 15802 5942 15804
rect 5966 15802 6022 15804
rect 6046 15802 6102 15804
rect 6126 15802 6182 15804
rect 5886 15750 5912 15802
rect 5912 15750 5942 15802
rect 5966 15750 5976 15802
rect 5976 15750 6022 15802
rect 6046 15750 6092 15802
rect 6092 15750 6102 15802
rect 6126 15750 6156 15802
rect 6156 15750 6182 15802
rect 5886 15748 5942 15750
rect 5966 15748 6022 15750
rect 6046 15748 6102 15750
rect 6126 15748 6182 15750
rect 5886 14714 5942 14716
rect 5966 14714 6022 14716
rect 6046 14714 6102 14716
rect 6126 14714 6182 14716
rect 5886 14662 5912 14714
rect 5912 14662 5942 14714
rect 5966 14662 5976 14714
rect 5976 14662 6022 14714
rect 6046 14662 6092 14714
rect 6092 14662 6102 14714
rect 6126 14662 6156 14714
rect 6156 14662 6182 14714
rect 5886 14660 5942 14662
rect 5966 14660 6022 14662
rect 6046 14660 6102 14662
rect 6126 14660 6182 14662
rect 5886 13626 5942 13628
rect 5966 13626 6022 13628
rect 6046 13626 6102 13628
rect 6126 13626 6182 13628
rect 5886 13574 5912 13626
rect 5912 13574 5942 13626
rect 5966 13574 5976 13626
rect 5976 13574 6022 13626
rect 6046 13574 6092 13626
rect 6092 13574 6102 13626
rect 6126 13574 6156 13626
rect 6156 13574 6182 13626
rect 5886 13572 5942 13574
rect 5966 13572 6022 13574
rect 6046 13572 6102 13574
rect 6126 13572 6182 13574
rect 5886 12538 5942 12540
rect 5966 12538 6022 12540
rect 6046 12538 6102 12540
rect 6126 12538 6182 12540
rect 5886 12486 5912 12538
rect 5912 12486 5942 12538
rect 5966 12486 5976 12538
rect 5976 12486 6022 12538
rect 6046 12486 6092 12538
rect 6092 12486 6102 12538
rect 6126 12486 6156 12538
rect 6156 12486 6182 12538
rect 5886 12484 5942 12486
rect 5966 12484 6022 12486
rect 6046 12484 6102 12486
rect 6126 12484 6182 12486
rect 5886 11450 5942 11452
rect 5966 11450 6022 11452
rect 6046 11450 6102 11452
rect 6126 11450 6182 11452
rect 5886 11398 5912 11450
rect 5912 11398 5942 11450
rect 5966 11398 5976 11450
rect 5976 11398 6022 11450
rect 6046 11398 6092 11450
rect 6092 11398 6102 11450
rect 6126 11398 6156 11450
rect 6156 11398 6182 11450
rect 5886 11396 5942 11398
rect 5966 11396 6022 11398
rect 6046 11396 6102 11398
rect 6126 11396 6182 11398
rect 5886 10362 5942 10364
rect 5966 10362 6022 10364
rect 6046 10362 6102 10364
rect 6126 10362 6182 10364
rect 5886 10310 5912 10362
rect 5912 10310 5942 10362
rect 5966 10310 5976 10362
rect 5976 10310 6022 10362
rect 6046 10310 6092 10362
rect 6092 10310 6102 10362
rect 6126 10310 6156 10362
rect 6156 10310 6182 10362
rect 5886 10308 5942 10310
rect 5966 10308 6022 10310
rect 6046 10308 6102 10310
rect 6126 10308 6182 10310
rect 5886 9274 5942 9276
rect 5966 9274 6022 9276
rect 6046 9274 6102 9276
rect 6126 9274 6182 9276
rect 5886 9222 5912 9274
rect 5912 9222 5942 9274
rect 5966 9222 5976 9274
rect 5976 9222 6022 9274
rect 6046 9222 6092 9274
rect 6092 9222 6102 9274
rect 6126 9222 6156 9274
rect 6156 9222 6182 9274
rect 5886 9220 5942 9222
rect 5966 9220 6022 9222
rect 6046 9220 6102 9222
rect 6126 9220 6182 9222
rect 5886 8186 5942 8188
rect 5966 8186 6022 8188
rect 6046 8186 6102 8188
rect 6126 8186 6182 8188
rect 5886 8134 5912 8186
rect 5912 8134 5942 8186
rect 5966 8134 5976 8186
rect 5976 8134 6022 8186
rect 6046 8134 6092 8186
rect 6092 8134 6102 8186
rect 6126 8134 6156 8186
rect 6156 8134 6182 8186
rect 5886 8132 5942 8134
rect 5966 8132 6022 8134
rect 6046 8132 6102 8134
rect 6126 8132 6182 8134
rect 5886 7098 5942 7100
rect 5966 7098 6022 7100
rect 6046 7098 6102 7100
rect 6126 7098 6182 7100
rect 5886 7046 5912 7098
rect 5912 7046 5942 7098
rect 5966 7046 5976 7098
rect 5976 7046 6022 7098
rect 6046 7046 6092 7098
rect 6092 7046 6102 7098
rect 6126 7046 6156 7098
rect 6156 7046 6182 7098
rect 5886 7044 5942 7046
rect 5966 7044 6022 7046
rect 6046 7044 6102 7046
rect 6126 7044 6182 7046
rect 5886 6010 5942 6012
rect 5966 6010 6022 6012
rect 6046 6010 6102 6012
rect 6126 6010 6182 6012
rect 5886 5958 5912 6010
rect 5912 5958 5942 6010
rect 5966 5958 5976 6010
rect 5976 5958 6022 6010
rect 6046 5958 6092 6010
rect 6092 5958 6102 6010
rect 6126 5958 6156 6010
rect 6156 5958 6182 6010
rect 5886 5956 5942 5958
rect 5966 5956 6022 5958
rect 6046 5956 6102 5958
rect 6126 5956 6182 5958
rect 5886 4922 5942 4924
rect 5966 4922 6022 4924
rect 6046 4922 6102 4924
rect 6126 4922 6182 4924
rect 5886 4870 5912 4922
rect 5912 4870 5942 4922
rect 5966 4870 5976 4922
rect 5976 4870 6022 4922
rect 6046 4870 6092 4922
rect 6092 4870 6102 4922
rect 6126 4870 6156 4922
rect 6156 4870 6182 4922
rect 5886 4868 5942 4870
rect 5966 4868 6022 4870
rect 6046 4868 6102 4870
rect 6126 4868 6182 4870
rect 5886 3834 5942 3836
rect 5966 3834 6022 3836
rect 6046 3834 6102 3836
rect 6126 3834 6182 3836
rect 5886 3782 5912 3834
rect 5912 3782 5942 3834
rect 5966 3782 5976 3834
rect 5976 3782 6022 3834
rect 6046 3782 6092 3834
rect 6092 3782 6102 3834
rect 6126 3782 6156 3834
rect 6156 3782 6182 3834
rect 5886 3780 5942 3782
rect 5966 3780 6022 3782
rect 6046 3780 6102 3782
rect 6126 3780 6182 3782
rect 5886 2746 5942 2748
rect 5966 2746 6022 2748
rect 6046 2746 6102 2748
rect 6126 2746 6182 2748
rect 5886 2694 5912 2746
rect 5912 2694 5942 2746
rect 5966 2694 5976 2746
rect 5976 2694 6022 2746
rect 6046 2694 6092 2746
rect 6092 2694 6102 2746
rect 6126 2694 6156 2746
rect 6156 2694 6182 2746
rect 5886 2692 5942 2694
rect 5966 2692 6022 2694
rect 6046 2692 6102 2694
rect 6126 2692 6182 2694
rect 8352 17434 8408 17436
rect 8432 17434 8488 17436
rect 8512 17434 8568 17436
rect 8592 17434 8648 17436
rect 8352 17382 8378 17434
rect 8378 17382 8408 17434
rect 8432 17382 8442 17434
rect 8442 17382 8488 17434
rect 8512 17382 8558 17434
rect 8558 17382 8568 17434
rect 8592 17382 8622 17434
rect 8622 17382 8648 17434
rect 8352 17380 8408 17382
rect 8432 17380 8488 17382
rect 8512 17380 8568 17382
rect 8592 17380 8648 17382
rect 8352 16346 8408 16348
rect 8432 16346 8488 16348
rect 8512 16346 8568 16348
rect 8592 16346 8648 16348
rect 8352 16294 8378 16346
rect 8378 16294 8408 16346
rect 8432 16294 8442 16346
rect 8442 16294 8488 16346
rect 8512 16294 8558 16346
rect 8558 16294 8568 16346
rect 8592 16294 8622 16346
rect 8622 16294 8648 16346
rect 8352 16292 8408 16294
rect 8432 16292 8488 16294
rect 8512 16292 8568 16294
rect 8592 16292 8648 16294
rect 8352 15258 8408 15260
rect 8432 15258 8488 15260
rect 8512 15258 8568 15260
rect 8592 15258 8648 15260
rect 8352 15206 8378 15258
rect 8378 15206 8408 15258
rect 8432 15206 8442 15258
rect 8442 15206 8488 15258
rect 8512 15206 8558 15258
rect 8558 15206 8568 15258
rect 8592 15206 8622 15258
rect 8622 15206 8648 15258
rect 8352 15204 8408 15206
rect 8432 15204 8488 15206
rect 8512 15204 8568 15206
rect 8592 15204 8648 15206
rect 8352 14170 8408 14172
rect 8432 14170 8488 14172
rect 8512 14170 8568 14172
rect 8592 14170 8648 14172
rect 8352 14118 8378 14170
rect 8378 14118 8408 14170
rect 8432 14118 8442 14170
rect 8442 14118 8488 14170
rect 8512 14118 8558 14170
rect 8558 14118 8568 14170
rect 8592 14118 8622 14170
rect 8622 14118 8648 14170
rect 8352 14116 8408 14118
rect 8432 14116 8488 14118
rect 8512 14116 8568 14118
rect 8592 14116 8648 14118
rect 8352 13082 8408 13084
rect 8432 13082 8488 13084
rect 8512 13082 8568 13084
rect 8592 13082 8648 13084
rect 8352 13030 8378 13082
rect 8378 13030 8408 13082
rect 8432 13030 8442 13082
rect 8442 13030 8488 13082
rect 8512 13030 8558 13082
rect 8558 13030 8568 13082
rect 8592 13030 8622 13082
rect 8622 13030 8648 13082
rect 8352 13028 8408 13030
rect 8432 13028 8488 13030
rect 8512 13028 8568 13030
rect 8592 13028 8648 13030
rect 8352 11994 8408 11996
rect 8432 11994 8488 11996
rect 8512 11994 8568 11996
rect 8592 11994 8648 11996
rect 8352 11942 8378 11994
rect 8378 11942 8408 11994
rect 8432 11942 8442 11994
rect 8442 11942 8488 11994
rect 8512 11942 8558 11994
rect 8558 11942 8568 11994
rect 8592 11942 8622 11994
rect 8622 11942 8648 11994
rect 8352 11940 8408 11942
rect 8432 11940 8488 11942
rect 8512 11940 8568 11942
rect 8592 11940 8648 11942
rect 8352 10906 8408 10908
rect 8432 10906 8488 10908
rect 8512 10906 8568 10908
rect 8592 10906 8648 10908
rect 8352 10854 8378 10906
rect 8378 10854 8408 10906
rect 8432 10854 8442 10906
rect 8442 10854 8488 10906
rect 8512 10854 8558 10906
rect 8558 10854 8568 10906
rect 8592 10854 8622 10906
rect 8622 10854 8648 10906
rect 8352 10852 8408 10854
rect 8432 10852 8488 10854
rect 8512 10852 8568 10854
rect 8592 10852 8648 10854
rect 8352 9818 8408 9820
rect 8432 9818 8488 9820
rect 8512 9818 8568 9820
rect 8592 9818 8648 9820
rect 8352 9766 8378 9818
rect 8378 9766 8408 9818
rect 8432 9766 8442 9818
rect 8442 9766 8488 9818
rect 8512 9766 8558 9818
rect 8558 9766 8568 9818
rect 8592 9766 8622 9818
rect 8622 9766 8648 9818
rect 8352 9764 8408 9766
rect 8432 9764 8488 9766
rect 8512 9764 8568 9766
rect 8592 9764 8648 9766
rect 8352 8730 8408 8732
rect 8432 8730 8488 8732
rect 8512 8730 8568 8732
rect 8592 8730 8648 8732
rect 8352 8678 8378 8730
rect 8378 8678 8408 8730
rect 8432 8678 8442 8730
rect 8442 8678 8488 8730
rect 8512 8678 8558 8730
rect 8558 8678 8568 8730
rect 8592 8678 8622 8730
rect 8622 8678 8648 8730
rect 8352 8676 8408 8678
rect 8432 8676 8488 8678
rect 8512 8676 8568 8678
rect 8592 8676 8648 8678
rect 8352 7642 8408 7644
rect 8432 7642 8488 7644
rect 8512 7642 8568 7644
rect 8592 7642 8648 7644
rect 8352 7590 8378 7642
rect 8378 7590 8408 7642
rect 8432 7590 8442 7642
rect 8442 7590 8488 7642
rect 8512 7590 8558 7642
rect 8558 7590 8568 7642
rect 8592 7590 8622 7642
rect 8622 7590 8648 7642
rect 8352 7588 8408 7590
rect 8432 7588 8488 7590
rect 8512 7588 8568 7590
rect 8592 7588 8648 7590
rect 8352 6554 8408 6556
rect 8432 6554 8488 6556
rect 8512 6554 8568 6556
rect 8592 6554 8648 6556
rect 8352 6502 8378 6554
rect 8378 6502 8408 6554
rect 8432 6502 8442 6554
rect 8442 6502 8488 6554
rect 8512 6502 8558 6554
rect 8558 6502 8568 6554
rect 8592 6502 8622 6554
rect 8622 6502 8648 6554
rect 8352 6500 8408 6502
rect 8432 6500 8488 6502
rect 8512 6500 8568 6502
rect 8592 6500 8648 6502
rect 8352 5466 8408 5468
rect 8432 5466 8488 5468
rect 8512 5466 8568 5468
rect 8592 5466 8648 5468
rect 8352 5414 8378 5466
rect 8378 5414 8408 5466
rect 8432 5414 8442 5466
rect 8442 5414 8488 5466
rect 8512 5414 8558 5466
rect 8558 5414 8568 5466
rect 8592 5414 8622 5466
rect 8622 5414 8648 5466
rect 8352 5412 8408 5414
rect 8432 5412 8488 5414
rect 8512 5412 8568 5414
rect 8592 5412 8648 5414
rect 8352 4378 8408 4380
rect 8432 4378 8488 4380
rect 8512 4378 8568 4380
rect 8592 4378 8648 4380
rect 8352 4326 8378 4378
rect 8378 4326 8408 4378
rect 8432 4326 8442 4378
rect 8442 4326 8488 4378
rect 8512 4326 8558 4378
rect 8558 4326 8568 4378
rect 8592 4326 8622 4378
rect 8622 4326 8648 4378
rect 8352 4324 8408 4326
rect 8432 4324 8488 4326
rect 8512 4324 8568 4326
rect 8592 4324 8648 4326
rect 8352 3290 8408 3292
rect 8432 3290 8488 3292
rect 8512 3290 8568 3292
rect 8592 3290 8648 3292
rect 8352 3238 8378 3290
rect 8378 3238 8408 3290
rect 8432 3238 8442 3290
rect 8442 3238 8488 3290
rect 8512 3238 8558 3290
rect 8558 3238 8568 3290
rect 8592 3238 8622 3290
rect 8622 3238 8648 3290
rect 8352 3236 8408 3238
rect 8432 3236 8488 3238
rect 8512 3236 8568 3238
rect 8592 3236 8648 3238
rect 8352 2202 8408 2204
rect 8432 2202 8488 2204
rect 8512 2202 8568 2204
rect 8592 2202 8648 2204
rect 8352 2150 8378 2202
rect 8378 2150 8408 2202
rect 8432 2150 8442 2202
rect 8442 2150 8488 2202
rect 8512 2150 8558 2202
rect 8558 2150 8568 2202
rect 8592 2150 8622 2202
rect 8622 2150 8648 2202
rect 8352 2148 8408 2150
rect 8432 2148 8488 2150
rect 8512 2148 8568 2150
rect 8592 2148 8648 2150
rect 9770 4120 9826 4176
rect 10817 16890 10873 16892
rect 10897 16890 10953 16892
rect 10977 16890 11033 16892
rect 11057 16890 11113 16892
rect 10817 16838 10843 16890
rect 10843 16838 10873 16890
rect 10897 16838 10907 16890
rect 10907 16838 10953 16890
rect 10977 16838 11023 16890
rect 11023 16838 11033 16890
rect 11057 16838 11087 16890
rect 11087 16838 11113 16890
rect 10817 16836 10873 16838
rect 10897 16836 10953 16838
rect 10977 16836 11033 16838
rect 11057 16836 11113 16838
rect 10817 15802 10873 15804
rect 10897 15802 10953 15804
rect 10977 15802 11033 15804
rect 11057 15802 11113 15804
rect 10817 15750 10843 15802
rect 10843 15750 10873 15802
rect 10897 15750 10907 15802
rect 10907 15750 10953 15802
rect 10977 15750 11023 15802
rect 11023 15750 11033 15802
rect 11057 15750 11087 15802
rect 11087 15750 11113 15802
rect 10817 15748 10873 15750
rect 10897 15748 10953 15750
rect 10977 15748 11033 15750
rect 11057 15748 11113 15750
rect 10817 14714 10873 14716
rect 10897 14714 10953 14716
rect 10977 14714 11033 14716
rect 11057 14714 11113 14716
rect 10817 14662 10843 14714
rect 10843 14662 10873 14714
rect 10897 14662 10907 14714
rect 10907 14662 10953 14714
rect 10977 14662 11023 14714
rect 11023 14662 11033 14714
rect 11057 14662 11087 14714
rect 11087 14662 11113 14714
rect 10817 14660 10873 14662
rect 10897 14660 10953 14662
rect 10977 14660 11033 14662
rect 11057 14660 11113 14662
rect 10817 13626 10873 13628
rect 10897 13626 10953 13628
rect 10977 13626 11033 13628
rect 11057 13626 11113 13628
rect 10817 13574 10843 13626
rect 10843 13574 10873 13626
rect 10897 13574 10907 13626
rect 10907 13574 10953 13626
rect 10977 13574 11023 13626
rect 11023 13574 11033 13626
rect 11057 13574 11087 13626
rect 11087 13574 11113 13626
rect 10817 13572 10873 13574
rect 10897 13572 10953 13574
rect 10977 13572 11033 13574
rect 11057 13572 11113 13574
rect 10817 12538 10873 12540
rect 10897 12538 10953 12540
rect 10977 12538 11033 12540
rect 11057 12538 11113 12540
rect 10817 12486 10843 12538
rect 10843 12486 10873 12538
rect 10897 12486 10907 12538
rect 10907 12486 10953 12538
rect 10977 12486 11023 12538
rect 11023 12486 11033 12538
rect 11057 12486 11087 12538
rect 11087 12486 11113 12538
rect 10817 12484 10873 12486
rect 10897 12484 10953 12486
rect 10977 12484 11033 12486
rect 11057 12484 11113 12486
rect 10817 11450 10873 11452
rect 10897 11450 10953 11452
rect 10977 11450 11033 11452
rect 11057 11450 11113 11452
rect 10817 11398 10843 11450
rect 10843 11398 10873 11450
rect 10897 11398 10907 11450
rect 10907 11398 10953 11450
rect 10977 11398 11023 11450
rect 11023 11398 11033 11450
rect 11057 11398 11087 11450
rect 11087 11398 11113 11450
rect 10817 11396 10873 11398
rect 10897 11396 10953 11398
rect 10977 11396 11033 11398
rect 11057 11396 11113 11398
rect 10817 10362 10873 10364
rect 10897 10362 10953 10364
rect 10977 10362 11033 10364
rect 11057 10362 11113 10364
rect 10817 10310 10843 10362
rect 10843 10310 10873 10362
rect 10897 10310 10907 10362
rect 10907 10310 10953 10362
rect 10977 10310 11023 10362
rect 11023 10310 11033 10362
rect 11057 10310 11087 10362
rect 11087 10310 11113 10362
rect 10817 10308 10873 10310
rect 10897 10308 10953 10310
rect 10977 10308 11033 10310
rect 11057 10308 11113 10310
rect 10817 9274 10873 9276
rect 10897 9274 10953 9276
rect 10977 9274 11033 9276
rect 11057 9274 11113 9276
rect 10817 9222 10843 9274
rect 10843 9222 10873 9274
rect 10897 9222 10907 9274
rect 10907 9222 10953 9274
rect 10977 9222 11023 9274
rect 11023 9222 11033 9274
rect 11057 9222 11087 9274
rect 11087 9222 11113 9274
rect 10817 9220 10873 9222
rect 10897 9220 10953 9222
rect 10977 9220 11033 9222
rect 11057 9220 11113 9222
rect 10817 8186 10873 8188
rect 10897 8186 10953 8188
rect 10977 8186 11033 8188
rect 11057 8186 11113 8188
rect 10817 8134 10843 8186
rect 10843 8134 10873 8186
rect 10897 8134 10907 8186
rect 10907 8134 10953 8186
rect 10977 8134 11023 8186
rect 11023 8134 11033 8186
rect 11057 8134 11087 8186
rect 11087 8134 11113 8186
rect 10817 8132 10873 8134
rect 10897 8132 10953 8134
rect 10977 8132 11033 8134
rect 11057 8132 11113 8134
rect 10817 7098 10873 7100
rect 10897 7098 10953 7100
rect 10977 7098 11033 7100
rect 11057 7098 11113 7100
rect 10817 7046 10843 7098
rect 10843 7046 10873 7098
rect 10897 7046 10907 7098
rect 10907 7046 10953 7098
rect 10977 7046 11023 7098
rect 11023 7046 11033 7098
rect 11057 7046 11087 7098
rect 11087 7046 11113 7098
rect 10817 7044 10873 7046
rect 10897 7044 10953 7046
rect 10977 7044 11033 7046
rect 11057 7044 11113 7046
rect 10817 6010 10873 6012
rect 10897 6010 10953 6012
rect 10977 6010 11033 6012
rect 11057 6010 11113 6012
rect 10817 5958 10843 6010
rect 10843 5958 10873 6010
rect 10897 5958 10907 6010
rect 10907 5958 10953 6010
rect 10977 5958 11023 6010
rect 11023 5958 11033 6010
rect 11057 5958 11087 6010
rect 11087 5958 11113 6010
rect 10817 5956 10873 5958
rect 10897 5956 10953 5958
rect 10977 5956 11033 5958
rect 11057 5956 11113 5958
rect 10817 4922 10873 4924
rect 10897 4922 10953 4924
rect 10977 4922 11033 4924
rect 11057 4922 11113 4924
rect 10817 4870 10843 4922
rect 10843 4870 10873 4922
rect 10897 4870 10907 4922
rect 10907 4870 10953 4922
rect 10977 4870 11023 4922
rect 11023 4870 11033 4922
rect 11057 4870 11087 4922
rect 11087 4870 11113 4922
rect 10817 4868 10873 4870
rect 10897 4868 10953 4870
rect 10977 4868 11033 4870
rect 11057 4868 11113 4870
rect 11334 4120 11390 4176
rect 10817 3834 10873 3836
rect 10897 3834 10953 3836
rect 10977 3834 11033 3836
rect 11057 3834 11113 3836
rect 10817 3782 10843 3834
rect 10843 3782 10873 3834
rect 10897 3782 10907 3834
rect 10907 3782 10953 3834
rect 10977 3782 11023 3834
rect 11023 3782 11033 3834
rect 11057 3782 11087 3834
rect 11087 3782 11113 3834
rect 10817 3780 10873 3782
rect 10897 3780 10953 3782
rect 10977 3780 11033 3782
rect 11057 3780 11113 3782
rect 10817 2746 10873 2748
rect 10897 2746 10953 2748
rect 10977 2746 11033 2748
rect 11057 2746 11113 2748
rect 10817 2694 10843 2746
rect 10843 2694 10873 2746
rect 10897 2694 10907 2746
rect 10907 2694 10953 2746
rect 10977 2694 11023 2746
rect 11023 2694 11033 2746
rect 11057 2694 11087 2746
rect 11087 2694 11113 2746
rect 10817 2692 10873 2694
rect 10897 2692 10953 2694
rect 10977 2692 11033 2694
rect 11057 2692 11113 2694
rect 12438 7384 12494 7440
rect 13726 17448 13782 17504
rect 13282 17434 13338 17436
rect 13362 17434 13418 17436
rect 13442 17434 13498 17436
rect 13522 17434 13578 17436
rect 13282 17382 13308 17434
rect 13308 17382 13338 17434
rect 13362 17382 13372 17434
rect 13372 17382 13418 17434
rect 13442 17382 13488 17434
rect 13488 17382 13498 17434
rect 13522 17382 13552 17434
rect 13552 17382 13578 17434
rect 13282 17380 13338 17382
rect 13362 17380 13418 17382
rect 13442 17380 13498 17382
rect 13522 17380 13578 17382
rect 13282 16346 13338 16348
rect 13362 16346 13418 16348
rect 13442 16346 13498 16348
rect 13522 16346 13578 16348
rect 13282 16294 13308 16346
rect 13308 16294 13338 16346
rect 13362 16294 13372 16346
rect 13372 16294 13418 16346
rect 13442 16294 13488 16346
rect 13488 16294 13498 16346
rect 13522 16294 13552 16346
rect 13552 16294 13578 16346
rect 13282 16292 13338 16294
rect 13362 16292 13418 16294
rect 13442 16292 13498 16294
rect 13522 16292 13578 16294
rect 13282 15258 13338 15260
rect 13362 15258 13418 15260
rect 13442 15258 13498 15260
rect 13522 15258 13578 15260
rect 13282 15206 13308 15258
rect 13308 15206 13338 15258
rect 13362 15206 13372 15258
rect 13372 15206 13418 15258
rect 13442 15206 13488 15258
rect 13488 15206 13498 15258
rect 13522 15206 13552 15258
rect 13552 15206 13578 15258
rect 13282 15204 13338 15206
rect 13362 15204 13418 15206
rect 13442 15204 13498 15206
rect 13522 15204 13578 15206
rect 13282 14170 13338 14172
rect 13362 14170 13418 14172
rect 13442 14170 13498 14172
rect 13522 14170 13578 14172
rect 13282 14118 13308 14170
rect 13308 14118 13338 14170
rect 13362 14118 13372 14170
rect 13372 14118 13418 14170
rect 13442 14118 13488 14170
rect 13488 14118 13498 14170
rect 13522 14118 13552 14170
rect 13552 14118 13578 14170
rect 13282 14116 13338 14118
rect 13362 14116 13418 14118
rect 13442 14116 13498 14118
rect 13522 14116 13578 14118
rect 13282 13082 13338 13084
rect 13362 13082 13418 13084
rect 13442 13082 13498 13084
rect 13522 13082 13578 13084
rect 13282 13030 13308 13082
rect 13308 13030 13338 13082
rect 13362 13030 13372 13082
rect 13372 13030 13418 13082
rect 13442 13030 13488 13082
rect 13488 13030 13498 13082
rect 13522 13030 13552 13082
rect 13552 13030 13578 13082
rect 13282 13028 13338 13030
rect 13362 13028 13418 13030
rect 13442 13028 13498 13030
rect 13522 13028 13578 13030
rect 13450 12416 13506 12472
rect 13282 11994 13338 11996
rect 13362 11994 13418 11996
rect 13442 11994 13498 11996
rect 13522 11994 13578 11996
rect 13282 11942 13308 11994
rect 13308 11942 13338 11994
rect 13362 11942 13372 11994
rect 13372 11942 13418 11994
rect 13442 11942 13488 11994
rect 13488 11942 13498 11994
rect 13522 11942 13552 11994
rect 13552 11942 13578 11994
rect 13282 11940 13338 11942
rect 13362 11940 13418 11942
rect 13442 11940 13498 11942
rect 13522 11940 13578 11942
rect 13282 10906 13338 10908
rect 13362 10906 13418 10908
rect 13442 10906 13498 10908
rect 13522 10906 13578 10908
rect 13282 10854 13308 10906
rect 13308 10854 13338 10906
rect 13362 10854 13372 10906
rect 13372 10854 13418 10906
rect 13442 10854 13488 10906
rect 13488 10854 13498 10906
rect 13522 10854 13552 10906
rect 13552 10854 13578 10906
rect 13282 10852 13338 10854
rect 13362 10852 13418 10854
rect 13442 10852 13498 10854
rect 13522 10852 13578 10854
rect 13282 9818 13338 9820
rect 13362 9818 13418 9820
rect 13442 9818 13498 9820
rect 13522 9818 13578 9820
rect 13282 9766 13308 9818
rect 13308 9766 13338 9818
rect 13362 9766 13372 9818
rect 13372 9766 13418 9818
rect 13442 9766 13488 9818
rect 13488 9766 13498 9818
rect 13522 9766 13552 9818
rect 13552 9766 13578 9818
rect 13282 9764 13338 9766
rect 13362 9764 13418 9766
rect 13442 9764 13498 9766
rect 13522 9764 13578 9766
rect 13282 8730 13338 8732
rect 13362 8730 13418 8732
rect 13442 8730 13498 8732
rect 13522 8730 13578 8732
rect 13282 8678 13308 8730
rect 13308 8678 13338 8730
rect 13362 8678 13372 8730
rect 13372 8678 13418 8730
rect 13442 8678 13488 8730
rect 13488 8678 13498 8730
rect 13522 8678 13552 8730
rect 13552 8678 13578 8730
rect 13282 8676 13338 8678
rect 13362 8676 13418 8678
rect 13442 8676 13498 8678
rect 13522 8676 13578 8678
rect 13282 7642 13338 7644
rect 13362 7642 13418 7644
rect 13442 7642 13498 7644
rect 13522 7642 13578 7644
rect 13282 7590 13308 7642
rect 13308 7590 13338 7642
rect 13362 7590 13372 7642
rect 13372 7590 13418 7642
rect 13442 7590 13488 7642
rect 13488 7590 13498 7642
rect 13522 7590 13552 7642
rect 13552 7590 13578 7642
rect 13282 7588 13338 7590
rect 13362 7588 13418 7590
rect 13442 7588 13498 7590
rect 13522 7588 13578 7590
rect 13282 6554 13338 6556
rect 13362 6554 13418 6556
rect 13442 6554 13498 6556
rect 13522 6554 13578 6556
rect 13282 6502 13308 6554
rect 13308 6502 13338 6554
rect 13362 6502 13372 6554
rect 13372 6502 13418 6554
rect 13442 6502 13488 6554
rect 13488 6502 13498 6554
rect 13522 6502 13552 6554
rect 13552 6502 13578 6554
rect 13282 6500 13338 6502
rect 13362 6500 13418 6502
rect 13442 6500 13498 6502
rect 13522 6500 13578 6502
rect 13282 5466 13338 5468
rect 13362 5466 13418 5468
rect 13442 5466 13498 5468
rect 13522 5466 13578 5468
rect 13282 5414 13308 5466
rect 13308 5414 13338 5466
rect 13362 5414 13372 5466
rect 13372 5414 13418 5466
rect 13442 5414 13488 5466
rect 13488 5414 13498 5466
rect 13522 5414 13552 5466
rect 13552 5414 13578 5466
rect 13282 5412 13338 5414
rect 13362 5412 13418 5414
rect 13442 5412 13498 5414
rect 13522 5412 13578 5414
rect 13282 4378 13338 4380
rect 13362 4378 13418 4380
rect 13442 4378 13498 4380
rect 13522 4378 13578 4380
rect 13282 4326 13308 4378
rect 13308 4326 13338 4378
rect 13362 4326 13372 4378
rect 13372 4326 13418 4378
rect 13442 4326 13488 4378
rect 13488 4326 13498 4378
rect 13522 4326 13552 4378
rect 13552 4326 13578 4378
rect 13282 4324 13338 4326
rect 13362 4324 13418 4326
rect 13442 4324 13498 4326
rect 13522 4324 13578 4326
rect 13282 3290 13338 3292
rect 13362 3290 13418 3292
rect 13442 3290 13498 3292
rect 13522 3290 13578 3292
rect 13282 3238 13308 3290
rect 13308 3238 13338 3290
rect 13362 3238 13372 3290
rect 13372 3238 13418 3290
rect 13442 3238 13488 3290
rect 13488 3238 13498 3290
rect 13522 3238 13552 3290
rect 13552 3238 13578 3290
rect 13282 3236 13338 3238
rect 13362 3236 13418 3238
rect 13442 3236 13498 3238
rect 13522 3236 13578 3238
rect 13634 2488 13690 2544
rect 13282 2202 13338 2204
rect 13362 2202 13418 2204
rect 13442 2202 13498 2204
rect 13522 2202 13578 2204
rect 13282 2150 13308 2202
rect 13308 2150 13338 2202
rect 13362 2150 13372 2202
rect 13372 2150 13418 2202
rect 13442 2150 13488 2202
rect 13488 2150 13498 2202
rect 13522 2150 13552 2202
rect 13552 2150 13578 2202
rect 13282 2148 13338 2150
rect 13362 2148 13418 2150
rect 13442 2148 13498 2150
rect 13522 2148 13578 2150
<< metal3 >>
rect 0 18322 480 18352
rect 3969 18322 4035 18325
rect 0 18320 4035 18322
rect 0 18264 3974 18320
rect 4030 18264 4035 18320
rect 0 18262 4035 18264
rect 0 18232 480 18262
rect 3969 18259 4035 18262
rect 13721 17506 13787 17509
rect 16520 17506 17000 17536
rect 13721 17504 17000 17506
rect 13721 17448 13726 17504
rect 13782 17448 17000 17504
rect 13721 17446 17000 17448
rect 13721 17443 13787 17446
rect 3409 17440 3729 17441
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 17375 3729 17376
rect 8340 17440 8660 17441
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 17375 8660 17376
rect 13270 17440 13590 17441
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 16520 17416 17000 17446
rect 13270 17375 13590 17376
rect 5874 16896 6194 16897
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6194 16896
rect 5874 16831 6194 16832
rect 10805 16896 11125 16897
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 16831 11125 16832
rect 3409 16352 3729 16353
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 16287 3729 16288
rect 8340 16352 8660 16353
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 16287 8660 16288
rect 13270 16352 13590 16353
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 16287 13590 16288
rect 5874 15808 6194 15809
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6194 15808
rect 5874 15743 6194 15744
rect 10805 15808 11125 15809
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 15743 11125 15744
rect 3409 15264 3729 15265
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 15199 3729 15200
rect 8340 15264 8660 15265
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 15199 8660 15200
rect 13270 15264 13590 15265
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 15199 13590 15200
rect 0 15058 480 15088
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14968 480 14998
rect 2773 14995 2839 14998
rect 5874 14720 6194 14721
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6194 14720
rect 5874 14655 6194 14656
rect 10805 14720 11125 14721
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 14655 11125 14656
rect 3409 14176 3729 14177
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 14111 3729 14112
rect 8340 14176 8660 14177
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 14111 8660 14112
rect 13270 14176 13590 14177
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 14111 13590 14112
rect 5874 13632 6194 13633
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6194 13632
rect 5874 13567 6194 13568
rect 10805 13632 11125 13633
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 13567 11125 13568
rect 3409 13088 3729 13089
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 13023 3729 13024
rect 8340 13088 8660 13089
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 13023 8660 13024
rect 13270 13088 13590 13089
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 13023 13590 13024
rect 5874 12544 6194 12545
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6194 12544
rect 5874 12479 6194 12480
rect 10805 12544 11125 12545
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 12479 11125 12480
rect 13445 12474 13511 12477
rect 16520 12474 17000 12504
rect 13445 12472 17000 12474
rect 13445 12416 13450 12472
rect 13506 12416 17000 12472
rect 13445 12414 17000 12416
rect 13445 12411 13511 12414
rect 16520 12384 17000 12414
rect 3409 12000 3729 12001
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 11935 3729 11936
rect 8340 12000 8660 12001
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 11935 8660 11936
rect 13270 12000 13590 12001
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 11935 13590 11936
rect 0 11658 480 11688
rect 3141 11658 3207 11661
rect 0 11656 3207 11658
rect 0 11600 3146 11656
rect 3202 11600 3207 11656
rect 0 11598 3207 11600
rect 0 11568 480 11598
rect 3141 11595 3207 11598
rect 5874 11456 6194 11457
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6194 11456
rect 5874 11391 6194 11392
rect 10805 11456 11125 11457
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 11391 11125 11392
rect 3409 10912 3729 10913
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 10847 3729 10848
rect 8340 10912 8660 10913
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 10847 8660 10848
rect 13270 10912 13590 10913
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 10847 13590 10848
rect 5874 10368 6194 10369
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6194 10368
rect 5874 10303 6194 10304
rect 10805 10368 11125 10369
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 10303 11125 10304
rect 3409 9824 3729 9825
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 9759 3729 9760
rect 8340 9824 8660 9825
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 9759 8660 9760
rect 13270 9824 13590 9825
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 9759 13590 9760
rect 5874 9280 6194 9281
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6194 9280
rect 5874 9215 6194 9216
rect 10805 9280 11125 9281
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 9215 11125 9216
rect 3409 8736 3729 8737
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 8671 3729 8672
rect 8340 8736 8660 8737
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 8671 8660 8672
rect 13270 8736 13590 8737
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 8671 13590 8672
rect 0 8394 480 8424
rect 2773 8394 2839 8397
rect 0 8392 2839 8394
rect 0 8336 2778 8392
rect 2834 8336 2839 8392
rect 0 8334 2839 8336
rect 0 8304 480 8334
rect 2773 8331 2839 8334
rect 5874 8192 6194 8193
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6194 8192
rect 5874 8127 6194 8128
rect 10805 8192 11125 8193
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 8127 11125 8128
rect 3409 7648 3729 7649
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 7583 3729 7584
rect 8340 7648 8660 7649
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 7583 8660 7584
rect 13270 7648 13590 7649
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 7583 13590 7584
rect 12433 7442 12499 7445
rect 16520 7442 17000 7472
rect 12433 7440 17000 7442
rect 12433 7384 12438 7440
rect 12494 7384 17000 7440
rect 12433 7382 17000 7384
rect 12433 7379 12499 7382
rect 16520 7352 17000 7382
rect 5874 7104 6194 7105
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6194 7104
rect 5874 7039 6194 7040
rect 10805 7104 11125 7105
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 7039 11125 7040
rect 3409 6560 3729 6561
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 6495 3729 6496
rect 8340 6560 8660 6561
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 6495 8660 6496
rect 13270 6560 13590 6561
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 6495 13590 6496
rect 5874 6016 6194 6017
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6194 6016
rect 5874 5951 6194 5952
rect 10805 6016 11125 6017
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 5951 11125 5952
rect 3409 5472 3729 5473
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 5407 3729 5408
rect 8340 5472 8660 5473
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 5407 8660 5408
rect 13270 5472 13590 5473
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 5407 13590 5408
rect 0 4994 480 5024
rect 3049 4994 3115 4997
rect 0 4992 3115 4994
rect 0 4936 3054 4992
rect 3110 4936 3115 4992
rect 0 4934 3115 4936
rect 0 4904 480 4934
rect 3049 4931 3115 4934
rect 5874 4928 6194 4929
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6194 4928
rect 5874 4863 6194 4864
rect 10805 4928 11125 4929
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 4863 11125 4864
rect 3409 4384 3729 4385
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 4319 3729 4320
rect 8340 4384 8660 4385
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 4319 8660 4320
rect 13270 4384 13590 4385
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 4319 13590 4320
rect 9765 4178 9831 4181
rect 11329 4178 11395 4181
rect 9765 4176 11395 4178
rect 9765 4120 9770 4176
rect 9826 4120 11334 4176
rect 11390 4120 11395 4176
rect 9765 4118 11395 4120
rect 9765 4115 9831 4118
rect 11329 4115 11395 4118
rect 5874 3840 6194 3841
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6194 3840
rect 5874 3775 6194 3776
rect 10805 3840 11125 3841
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 3775 11125 3776
rect 3409 3296 3729 3297
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 3231 3729 3232
rect 8340 3296 8660 3297
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 3231 8660 3232
rect 13270 3296 13590 3297
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 3231 13590 3232
rect 5874 2752 6194 2753
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6194 2752
rect 5874 2687 6194 2688
rect 10805 2752 11125 2753
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2687 11125 2688
rect 13629 2546 13695 2549
rect 16520 2546 17000 2576
rect 13629 2544 17000 2546
rect 13629 2488 13634 2544
rect 13690 2488 17000 2544
rect 13629 2486 17000 2488
rect 13629 2483 13695 2486
rect 16520 2456 17000 2486
rect 3409 2208 3729 2209
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2143 3729 2144
rect 8340 2208 8660 2209
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2143 8660 2144
rect 13270 2208 13590 2209
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2143 13590 2144
rect 0 1730 480 1760
rect 2957 1730 3023 1733
rect 0 1728 3023 1730
rect 0 1672 2962 1728
rect 3018 1672 3023 1728
rect 0 1670 3023 1672
rect 0 1640 480 1670
rect 2957 1667 3023 1670
<< via3 >>
rect 3417 17436 3481 17440
rect 3417 17380 3421 17436
rect 3421 17380 3477 17436
rect 3477 17380 3481 17436
rect 3417 17376 3481 17380
rect 3497 17436 3561 17440
rect 3497 17380 3501 17436
rect 3501 17380 3557 17436
rect 3557 17380 3561 17436
rect 3497 17376 3561 17380
rect 3577 17436 3641 17440
rect 3577 17380 3581 17436
rect 3581 17380 3637 17436
rect 3637 17380 3641 17436
rect 3577 17376 3641 17380
rect 3657 17436 3721 17440
rect 3657 17380 3661 17436
rect 3661 17380 3717 17436
rect 3717 17380 3721 17436
rect 3657 17376 3721 17380
rect 8348 17436 8412 17440
rect 8348 17380 8352 17436
rect 8352 17380 8408 17436
rect 8408 17380 8412 17436
rect 8348 17376 8412 17380
rect 8428 17436 8492 17440
rect 8428 17380 8432 17436
rect 8432 17380 8488 17436
rect 8488 17380 8492 17436
rect 8428 17376 8492 17380
rect 8508 17436 8572 17440
rect 8508 17380 8512 17436
rect 8512 17380 8568 17436
rect 8568 17380 8572 17436
rect 8508 17376 8572 17380
rect 8588 17436 8652 17440
rect 8588 17380 8592 17436
rect 8592 17380 8648 17436
rect 8648 17380 8652 17436
rect 8588 17376 8652 17380
rect 13278 17436 13342 17440
rect 13278 17380 13282 17436
rect 13282 17380 13338 17436
rect 13338 17380 13342 17436
rect 13278 17376 13342 17380
rect 13358 17436 13422 17440
rect 13358 17380 13362 17436
rect 13362 17380 13418 17436
rect 13418 17380 13422 17436
rect 13358 17376 13422 17380
rect 13438 17436 13502 17440
rect 13438 17380 13442 17436
rect 13442 17380 13498 17436
rect 13498 17380 13502 17436
rect 13438 17376 13502 17380
rect 13518 17436 13582 17440
rect 13518 17380 13522 17436
rect 13522 17380 13578 17436
rect 13578 17380 13582 17436
rect 13518 17376 13582 17380
rect 5882 16892 5946 16896
rect 5882 16836 5886 16892
rect 5886 16836 5942 16892
rect 5942 16836 5946 16892
rect 5882 16832 5946 16836
rect 5962 16892 6026 16896
rect 5962 16836 5966 16892
rect 5966 16836 6022 16892
rect 6022 16836 6026 16892
rect 5962 16832 6026 16836
rect 6042 16892 6106 16896
rect 6042 16836 6046 16892
rect 6046 16836 6102 16892
rect 6102 16836 6106 16892
rect 6042 16832 6106 16836
rect 6122 16892 6186 16896
rect 6122 16836 6126 16892
rect 6126 16836 6182 16892
rect 6182 16836 6186 16892
rect 6122 16832 6186 16836
rect 10813 16892 10877 16896
rect 10813 16836 10817 16892
rect 10817 16836 10873 16892
rect 10873 16836 10877 16892
rect 10813 16832 10877 16836
rect 10893 16892 10957 16896
rect 10893 16836 10897 16892
rect 10897 16836 10953 16892
rect 10953 16836 10957 16892
rect 10893 16832 10957 16836
rect 10973 16892 11037 16896
rect 10973 16836 10977 16892
rect 10977 16836 11033 16892
rect 11033 16836 11037 16892
rect 10973 16832 11037 16836
rect 11053 16892 11117 16896
rect 11053 16836 11057 16892
rect 11057 16836 11113 16892
rect 11113 16836 11117 16892
rect 11053 16832 11117 16836
rect 3417 16348 3481 16352
rect 3417 16292 3421 16348
rect 3421 16292 3477 16348
rect 3477 16292 3481 16348
rect 3417 16288 3481 16292
rect 3497 16348 3561 16352
rect 3497 16292 3501 16348
rect 3501 16292 3557 16348
rect 3557 16292 3561 16348
rect 3497 16288 3561 16292
rect 3577 16348 3641 16352
rect 3577 16292 3581 16348
rect 3581 16292 3637 16348
rect 3637 16292 3641 16348
rect 3577 16288 3641 16292
rect 3657 16348 3721 16352
rect 3657 16292 3661 16348
rect 3661 16292 3717 16348
rect 3717 16292 3721 16348
rect 3657 16288 3721 16292
rect 8348 16348 8412 16352
rect 8348 16292 8352 16348
rect 8352 16292 8408 16348
rect 8408 16292 8412 16348
rect 8348 16288 8412 16292
rect 8428 16348 8492 16352
rect 8428 16292 8432 16348
rect 8432 16292 8488 16348
rect 8488 16292 8492 16348
rect 8428 16288 8492 16292
rect 8508 16348 8572 16352
rect 8508 16292 8512 16348
rect 8512 16292 8568 16348
rect 8568 16292 8572 16348
rect 8508 16288 8572 16292
rect 8588 16348 8652 16352
rect 8588 16292 8592 16348
rect 8592 16292 8648 16348
rect 8648 16292 8652 16348
rect 8588 16288 8652 16292
rect 13278 16348 13342 16352
rect 13278 16292 13282 16348
rect 13282 16292 13338 16348
rect 13338 16292 13342 16348
rect 13278 16288 13342 16292
rect 13358 16348 13422 16352
rect 13358 16292 13362 16348
rect 13362 16292 13418 16348
rect 13418 16292 13422 16348
rect 13358 16288 13422 16292
rect 13438 16348 13502 16352
rect 13438 16292 13442 16348
rect 13442 16292 13498 16348
rect 13498 16292 13502 16348
rect 13438 16288 13502 16292
rect 13518 16348 13582 16352
rect 13518 16292 13522 16348
rect 13522 16292 13578 16348
rect 13578 16292 13582 16348
rect 13518 16288 13582 16292
rect 5882 15804 5946 15808
rect 5882 15748 5886 15804
rect 5886 15748 5942 15804
rect 5942 15748 5946 15804
rect 5882 15744 5946 15748
rect 5962 15804 6026 15808
rect 5962 15748 5966 15804
rect 5966 15748 6022 15804
rect 6022 15748 6026 15804
rect 5962 15744 6026 15748
rect 6042 15804 6106 15808
rect 6042 15748 6046 15804
rect 6046 15748 6102 15804
rect 6102 15748 6106 15804
rect 6042 15744 6106 15748
rect 6122 15804 6186 15808
rect 6122 15748 6126 15804
rect 6126 15748 6182 15804
rect 6182 15748 6186 15804
rect 6122 15744 6186 15748
rect 10813 15804 10877 15808
rect 10813 15748 10817 15804
rect 10817 15748 10873 15804
rect 10873 15748 10877 15804
rect 10813 15744 10877 15748
rect 10893 15804 10957 15808
rect 10893 15748 10897 15804
rect 10897 15748 10953 15804
rect 10953 15748 10957 15804
rect 10893 15744 10957 15748
rect 10973 15804 11037 15808
rect 10973 15748 10977 15804
rect 10977 15748 11033 15804
rect 11033 15748 11037 15804
rect 10973 15744 11037 15748
rect 11053 15804 11117 15808
rect 11053 15748 11057 15804
rect 11057 15748 11113 15804
rect 11113 15748 11117 15804
rect 11053 15744 11117 15748
rect 3417 15260 3481 15264
rect 3417 15204 3421 15260
rect 3421 15204 3477 15260
rect 3477 15204 3481 15260
rect 3417 15200 3481 15204
rect 3497 15260 3561 15264
rect 3497 15204 3501 15260
rect 3501 15204 3557 15260
rect 3557 15204 3561 15260
rect 3497 15200 3561 15204
rect 3577 15260 3641 15264
rect 3577 15204 3581 15260
rect 3581 15204 3637 15260
rect 3637 15204 3641 15260
rect 3577 15200 3641 15204
rect 3657 15260 3721 15264
rect 3657 15204 3661 15260
rect 3661 15204 3717 15260
rect 3717 15204 3721 15260
rect 3657 15200 3721 15204
rect 8348 15260 8412 15264
rect 8348 15204 8352 15260
rect 8352 15204 8408 15260
rect 8408 15204 8412 15260
rect 8348 15200 8412 15204
rect 8428 15260 8492 15264
rect 8428 15204 8432 15260
rect 8432 15204 8488 15260
rect 8488 15204 8492 15260
rect 8428 15200 8492 15204
rect 8508 15260 8572 15264
rect 8508 15204 8512 15260
rect 8512 15204 8568 15260
rect 8568 15204 8572 15260
rect 8508 15200 8572 15204
rect 8588 15260 8652 15264
rect 8588 15204 8592 15260
rect 8592 15204 8648 15260
rect 8648 15204 8652 15260
rect 8588 15200 8652 15204
rect 13278 15260 13342 15264
rect 13278 15204 13282 15260
rect 13282 15204 13338 15260
rect 13338 15204 13342 15260
rect 13278 15200 13342 15204
rect 13358 15260 13422 15264
rect 13358 15204 13362 15260
rect 13362 15204 13418 15260
rect 13418 15204 13422 15260
rect 13358 15200 13422 15204
rect 13438 15260 13502 15264
rect 13438 15204 13442 15260
rect 13442 15204 13498 15260
rect 13498 15204 13502 15260
rect 13438 15200 13502 15204
rect 13518 15260 13582 15264
rect 13518 15204 13522 15260
rect 13522 15204 13578 15260
rect 13578 15204 13582 15260
rect 13518 15200 13582 15204
rect 5882 14716 5946 14720
rect 5882 14660 5886 14716
rect 5886 14660 5942 14716
rect 5942 14660 5946 14716
rect 5882 14656 5946 14660
rect 5962 14716 6026 14720
rect 5962 14660 5966 14716
rect 5966 14660 6022 14716
rect 6022 14660 6026 14716
rect 5962 14656 6026 14660
rect 6042 14716 6106 14720
rect 6042 14660 6046 14716
rect 6046 14660 6102 14716
rect 6102 14660 6106 14716
rect 6042 14656 6106 14660
rect 6122 14716 6186 14720
rect 6122 14660 6126 14716
rect 6126 14660 6182 14716
rect 6182 14660 6186 14716
rect 6122 14656 6186 14660
rect 10813 14716 10877 14720
rect 10813 14660 10817 14716
rect 10817 14660 10873 14716
rect 10873 14660 10877 14716
rect 10813 14656 10877 14660
rect 10893 14716 10957 14720
rect 10893 14660 10897 14716
rect 10897 14660 10953 14716
rect 10953 14660 10957 14716
rect 10893 14656 10957 14660
rect 10973 14716 11037 14720
rect 10973 14660 10977 14716
rect 10977 14660 11033 14716
rect 11033 14660 11037 14716
rect 10973 14656 11037 14660
rect 11053 14716 11117 14720
rect 11053 14660 11057 14716
rect 11057 14660 11113 14716
rect 11113 14660 11117 14716
rect 11053 14656 11117 14660
rect 3417 14172 3481 14176
rect 3417 14116 3421 14172
rect 3421 14116 3477 14172
rect 3477 14116 3481 14172
rect 3417 14112 3481 14116
rect 3497 14172 3561 14176
rect 3497 14116 3501 14172
rect 3501 14116 3557 14172
rect 3557 14116 3561 14172
rect 3497 14112 3561 14116
rect 3577 14172 3641 14176
rect 3577 14116 3581 14172
rect 3581 14116 3637 14172
rect 3637 14116 3641 14172
rect 3577 14112 3641 14116
rect 3657 14172 3721 14176
rect 3657 14116 3661 14172
rect 3661 14116 3717 14172
rect 3717 14116 3721 14172
rect 3657 14112 3721 14116
rect 8348 14172 8412 14176
rect 8348 14116 8352 14172
rect 8352 14116 8408 14172
rect 8408 14116 8412 14172
rect 8348 14112 8412 14116
rect 8428 14172 8492 14176
rect 8428 14116 8432 14172
rect 8432 14116 8488 14172
rect 8488 14116 8492 14172
rect 8428 14112 8492 14116
rect 8508 14172 8572 14176
rect 8508 14116 8512 14172
rect 8512 14116 8568 14172
rect 8568 14116 8572 14172
rect 8508 14112 8572 14116
rect 8588 14172 8652 14176
rect 8588 14116 8592 14172
rect 8592 14116 8648 14172
rect 8648 14116 8652 14172
rect 8588 14112 8652 14116
rect 13278 14172 13342 14176
rect 13278 14116 13282 14172
rect 13282 14116 13338 14172
rect 13338 14116 13342 14172
rect 13278 14112 13342 14116
rect 13358 14172 13422 14176
rect 13358 14116 13362 14172
rect 13362 14116 13418 14172
rect 13418 14116 13422 14172
rect 13358 14112 13422 14116
rect 13438 14172 13502 14176
rect 13438 14116 13442 14172
rect 13442 14116 13498 14172
rect 13498 14116 13502 14172
rect 13438 14112 13502 14116
rect 13518 14172 13582 14176
rect 13518 14116 13522 14172
rect 13522 14116 13578 14172
rect 13578 14116 13582 14172
rect 13518 14112 13582 14116
rect 5882 13628 5946 13632
rect 5882 13572 5886 13628
rect 5886 13572 5942 13628
rect 5942 13572 5946 13628
rect 5882 13568 5946 13572
rect 5962 13628 6026 13632
rect 5962 13572 5966 13628
rect 5966 13572 6022 13628
rect 6022 13572 6026 13628
rect 5962 13568 6026 13572
rect 6042 13628 6106 13632
rect 6042 13572 6046 13628
rect 6046 13572 6102 13628
rect 6102 13572 6106 13628
rect 6042 13568 6106 13572
rect 6122 13628 6186 13632
rect 6122 13572 6126 13628
rect 6126 13572 6182 13628
rect 6182 13572 6186 13628
rect 6122 13568 6186 13572
rect 10813 13628 10877 13632
rect 10813 13572 10817 13628
rect 10817 13572 10873 13628
rect 10873 13572 10877 13628
rect 10813 13568 10877 13572
rect 10893 13628 10957 13632
rect 10893 13572 10897 13628
rect 10897 13572 10953 13628
rect 10953 13572 10957 13628
rect 10893 13568 10957 13572
rect 10973 13628 11037 13632
rect 10973 13572 10977 13628
rect 10977 13572 11033 13628
rect 11033 13572 11037 13628
rect 10973 13568 11037 13572
rect 11053 13628 11117 13632
rect 11053 13572 11057 13628
rect 11057 13572 11113 13628
rect 11113 13572 11117 13628
rect 11053 13568 11117 13572
rect 3417 13084 3481 13088
rect 3417 13028 3421 13084
rect 3421 13028 3477 13084
rect 3477 13028 3481 13084
rect 3417 13024 3481 13028
rect 3497 13084 3561 13088
rect 3497 13028 3501 13084
rect 3501 13028 3557 13084
rect 3557 13028 3561 13084
rect 3497 13024 3561 13028
rect 3577 13084 3641 13088
rect 3577 13028 3581 13084
rect 3581 13028 3637 13084
rect 3637 13028 3641 13084
rect 3577 13024 3641 13028
rect 3657 13084 3721 13088
rect 3657 13028 3661 13084
rect 3661 13028 3717 13084
rect 3717 13028 3721 13084
rect 3657 13024 3721 13028
rect 8348 13084 8412 13088
rect 8348 13028 8352 13084
rect 8352 13028 8408 13084
rect 8408 13028 8412 13084
rect 8348 13024 8412 13028
rect 8428 13084 8492 13088
rect 8428 13028 8432 13084
rect 8432 13028 8488 13084
rect 8488 13028 8492 13084
rect 8428 13024 8492 13028
rect 8508 13084 8572 13088
rect 8508 13028 8512 13084
rect 8512 13028 8568 13084
rect 8568 13028 8572 13084
rect 8508 13024 8572 13028
rect 8588 13084 8652 13088
rect 8588 13028 8592 13084
rect 8592 13028 8648 13084
rect 8648 13028 8652 13084
rect 8588 13024 8652 13028
rect 13278 13084 13342 13088
rect 13278 13028 13282 13084
rect 13282 13028 13338 13084
rect 13338 13028 13342 13084
rect 13278 13024 13342 13028
rect 13358 13084 13422 13088
rect 13358 13028 13362 13084
rect 13362 13028 13418 13084
rect 13418 13028 13422 13084
rect 13358 13024 13422 13028
rect 13438 13084 13502 13088
rect 13438 13028 13442 13084
rect 13442 13028 13498 13084
rect 13498 13028 13502 13084
rect 13438 13024 13502 13028
rect 13518 13084 13582 13088
rect 13518 13028 13522 13084
rect 13522 13028 13578 13084
rect 13578 13028 13582 13084
rect 13518 13024 13582 13028
rect 5882 12540 5946 12544
rect 5882 12484 5886 12540
rect 5886 12484 5942 12540
rect 5942 12484 5946 12540
rect 5882 12480 5946 12484
rect 5962 12540 6026 12544
rect 5962 12484 5966 12540
rect 5966 12484 6022 12540
rect 6022 12484 6026 12540
rect 5962 12480 6026 12484
rect 6042 12540 6106 12544
rect 6042 12484 6046 12540
rect 6046 12484 6102 12540
rect 6102 12484 6106 12540
rect 6042 12480 6106 12484
rect 6122 12540 6186 12544
rect 6122 12484 6126 12540
rect 6126 12484 6182 12540
rect 6182 12484 6186 12540
rect 6122 12480 6186 12484
rect 10813 12540 10877 12544
rect 10813 12484 10817 12540
rect 10817 12484 10873 12540
rect 10873 12484 10877 12540
rect 10813 12480 10877 12484
rect 10893 12540 10957 12544
rect 10893 12484 10897 12540
rect 10897 12484 10953 12540
rect 10953 12484 10957 12540
rect 10893 12480 10957 12484
rect 10973 12540 11037 12544
rect 10973 12484 10977 12540
rect 10977 12484 11033 12540
rect 11033 12484 11037 12540
rect 10973 12480 11037 12484
rect 11053 12540 11117 12544
rect 11053 12484 11057 12540
rect 11057 12484 11113 12540
rect 11113 12484 11117 12540
rect 11053 12480 11117 12484
rect 3417 11996 3481 12000
rect 3417 11940 3421 11996
rect 3421 11940 3477 11996
rect 3477 11940 3481 11996
rect 3417 11936 3481 11940
rect 3497 11996 3561 12000
rect 3497 11940 3501 11996
rect 3501 11940 3557 11996
rect 3557 11940 3561 11996
rect 3497 11936 3561 11940
rect 3577 11996 3641 12000
rect 3577 11940 3581 11996
rect 3581 11940 3637 11996
rect 3637 11940 3641 11996
rect 3577 11936 3641 11940
rect 3657 11996 3721 12000
rect 3657 11940 3661 11996
rect 3661 11940 3717 11996
rect 3717 11940 3721 11996
rect 3657 11936 3721 11940
rect 8348 11996 8412 12000
rect 8348 11940 8352 11996
rect 8352 11940 8408 11996
rect 8408 11940 8412 11996
rect 8348 11936 8412 11940
rect 8428 11996 8492 12000
rect 8428 11940 8432 11996
rect 8432 11940 8488 11996
rect 8488 11940 8492 11996
rect 8428 11936 8492 11940
rect 8508 11996 8572 12000
rect 8508 11940 8512 11996
rect 8512 11940 8568 11996
rect 8568 11940 8572 11996
rect 8508 11936 8572 11940
rect 8588 11996 8652 12000
rect 8588 11940 8592 11996
rect 8592 11940 8648 11996
rect 8648 11940 8652 11996
rect 8588 11936 8652 11940
rect 13278 11996 13342 12000
rect 13278 11940 13282 11996
rect 13282 11940 13338 11996
rect 13338 11940 13342 11996
rect 13278 11936 13342 11940
rect 13358 11996 13422 12000
rect 13358 11940 13362 11996
rect 13362 11940 13418 11996
rect 13418 11940 13422 11996
rect 13358 11936 13422 11940
rect 13438 11996 13502 12000
rect 13438 11940 13442 11996
rect 13442 11940 13498 11996
rect 13498 11940 13502 11996
rect 13438 11936 13502 11940
rect 13518 11996 13582 12000
rect 13518 11940 13522 11996
rect 13522 11940 13578 11996
rect 13578 11940 13582 11996
rect 13518 11936 13582 11940
rect 5882 11452 5946 11456
rect 5882 11396 5886 11452
rect 5886 11396 5942 11452
rect 5942 11396 5946 11452
rect 5882 11392 5946 11396
rect 5962 11452 6026 11456
rect 5962 11396 5966 11452
rect 5966 11396 6022 11452
rect 6022 11396 6026 11452
rect 5962 11392 6026 11396
rect 6042 11452 6106 11456
rect 6042 11396 6046 11452
rect 6046 11396 6102 11452
rect 6102 11396 6106 11452
rect 6042 11392 6106 11396
rect 6122 11452 6186 11456
rect 6122 11396 6126 11452
rect 6126 11396 6182 11452
rect 6182 11396 6186 11452
rect 6122 11392 6186 11396
rect 10813 11452 10877 11456
rect 10813 11396 10817 11452
rect 10817 11396 10873 11452
rect 10873 11396 10877 11452
rect 10813 11392 10877 11396
rect 10893 11452 10957 11456
rect 10893 11396 10897 11452
rect 10897 11396 10953 11452
rect 10953 11396 10957 11452
rect 10893 11392 10957 11396
rect 10973 11452 11037 11456
rect 10973 11396 10977 11452
rect 10977 11396 11033 11452
rect 11033 11396 11037 11452
rect 10973 11392 11037 11396
rect 11053 11452 11117 11456
rect 11053 11396 11057 11452
rect 11057 11396 11113 11452
rect 11113 11396 11117 11452
rect 11053 11392 11117 11396
rect 3417 10908 3481 10912
rect 3417 10852 3421 10908
rect 3421 10852 3477 10908
rect 3477 10852 3481 10908
rect 3417 10848 3481 10852
rect 3497 10908 3561 10912
rect 3497 10852 3501 10908
rect 3501 10852 3557 10908
rect 3557 10852 3561 10908
rect 3497 10848 3561 10852
rect 3577 10908 3641 10912
rect 3577 10852 3581 10908
rect 3581 10852 3637 10908
rect 3637 10852 3641 10908
rect 3577 10848 3641 10852
rect 3657 10908 3721 10912
rect 3657 10852 3661 10908
rect 3661 10852 3717 10908
rect 3717 10852 3721 10908
rect 3657 10848 3721 10852
rect 8348 10908 8412 10912
rect 8348 10852 8352 10908
rect 8352 10852 8408 10908
rect 8408 10852 8412 10908
rect 8348 10848 8412 10852
rect 8428 10908 8492 10912
rect 8428 10852 8432 10908
rect 8432 10852 8488 10908
rect 8488 10852 8492 10908
rect 8428 10848 8492 10852
rect 8508 10908 8572 10912
rect 8508 10852 8512 10908
rect 8512 10852 8568 10908
rect 8568 10852 8572 10908
rect 8508 10848 8572 10852
rect 8588 10908 8652 10912
rect 8588 10852 8592 10908
rect 8592 10852 8648 10908
rect 8648 10852 8652 10908
rect 8588 10848 8652 10852
rect 13278 10908 13342 10912
rect 13278 10852 13282 10908
rect 13282 10852 13338 10908
rect 13338 10852 13342 10908
rect 13278 10848 13342 10852
rect 13358 10908 13422 10912
rect 13358 10852 13362 10908
rect 13362 10852 13418 10908
rect 13418 10852 13422 10908
rect 13358 10848 13422 10852
rect 13438 10908 13502 10912
rect 13438 10852 13442 10908
rect 13442 10852 13498 10908
rect 13498 10852 13502 10908
rect 13438 10848 13502 10852
rect 13518 10908 13582 10912
rect 13518 10852 13522 10908
rect 13522 10852 13578 10908
rect 13578 10852 13582 10908
rect 13518 10848 13582 10852
rect 5882 10364 5946 10368
rect 5882 10308 5886 10364
rect 5886 10308 5942 10364
rect 5942 10308 5946 10364
rect 5882 10304 5946 10308
rect 5962 10364 6026 10368
rect 5962 10308 5966 10364
rect 5966 10308 6022 10364
rect 6022 10308 6026 10364
rect 5962 10304 6026 10308
rect 6042 10364 6106 10368
rect 6042 10308 6046 10364
rect 6046 10308 6102 10364
rect 6102 10308 6106 10364
rect 6042 10304 6106 10308
rect 6122 10364 6186 10368
rect 6122 10308 6126 10364
rect 6126 10308 6182 10364
rect 6182 10308 6186 10364
rect 6122 10304 6186 10308
rect 10813 10364 10877 10368
rect 10813 10308 10817 10364
rect 10817 10308 10873 10364
rect 10873 10308 10877 10364
rect 10813 10304 10877 10308
rect 10893 10364 10957 10368
rect 10893 10308 10897 10364
rect 10897 10308 10953 10364
rect 10953 10308 10957 10364
rect 10893 10304 10957 10308
rect 10973 10364 11037 10368
rect 10973 10308 10977 10364
rect 10977 10308 11033 10364
rect 11033 10308 11037 10364
rect 10973 10304 11037 10308
rect 11053 10364 11117 10368
rect 11053 10308 11057 10364
rect 11057 10308 11113 10364
rect 11113 10308 11117 10364
rect 11053 10304 11117 10308
rect 3417 9820 3481 9824
rect 3417 9764 3421 9820
rect 3421 9764 3477 9820
rect 3477 9764 3481 9820
rect 3417 9760 3481 9764
rect 3497 9820 3561 9824
rect 3497 9764 3501 9820
rect 3501 9764 3557 9820
rect 3557 9764 3561 9820
rect 3497 9760 3561 9764
rect 3577 9820 3641 9824
rect 3577 9764 3581 9820
rect 3581 9764 3637 9820
rect 3637 9764 3641 9820
rect 3577 9760 3641 9764
rect 3657 9820 3721 9824
rect 3657 9764 3661 9820
rect 3661 9764 3717 9820
rect 3717 9764 3721 9820
rect 3657 9760 3721 9764
rect 8348 9820 8412 9824
rect 8348 9764 8352 9820
rect 8352 9764 8408 9820
rect 8408 9764 8412 9820
rect 8348 9760 8412 9764
rect 8428 9820 8492 9824
rect 8428 9764 8432 9820
rect 8432 9764 8488 9820
rect 8488 9764 8492 9820
rect 8428 9760 8492 9764
rect 8508 9820 8572 9824
rect 8508 9764 8512 9820
rect 8512 9764 8568 9820
rect 8568 9764 8572 9820
rect 8508 9760 8572 9764
rect 8588 9820 8652 9824
rect 8588 9764 8592 9820
rect 8592 9764 8648 9820
rect 8648 9764 8652 9820
rect 8588 9760 8652 9764
rect 13278 9820 13342 9824
rect 13278 9764 13282 9820
rect 13282 9764 13338 9820
rect 13338 9764 13342 9820
rect 13278 9760 13342 9764
rect 13358 9820 13422 9824
rect 13358 9764 13362 9820
rect 13362 9764 13418 9820
rect 13418 9764 13422 9820
rect 13358 9760 13422 9764
rect 13438 9820 13502 9824
rect 13438 9764 13442 9820
rect 13442 9764 13498 9820
rect 13498 9764 13502 9820
rect 13438 9760 13502 9764
rect 13518 9820 13582 9824
rect 13518 9764 13522 9820
rect 13522 9764 13578 9820
rect 13578 9764 13582 9820
rect 13518 9760 13582 9764
rect 5882 9276 5946 9280
rect 5882 9220 5886 9276
rect 5886 9220 5942 9276
rect 5942 9220 5946 9276
rect 5882 9216 5946 9220
rect 5962 9276 6026 9280
rect 5962 9220 5966 9276
rect 5966 9220 6022 9276
rect 6022 9220 6026 9276
rect 5962 9216 6026 9220
rect 6042 9276 6106 9280
rect 6042 9220 6046 9276
rect 6046 9220 6102 9276
rect 6102 9220 6106 9276
rect 6042 9216 6106 9220
rect 6122 9276 6186 9280
rect 6122 9220 6126 9276
rect 6126 9220 6182 9276
rect 6182 9220 6186 9276
rect 6122 9216 6186 9220
rect 10813 9276 10877 9280
rect 10813 9220 10817 9276
rect 10817 9220 10873 9276
rect 10873 9220 10877 9276
rect 10813 9216 10877 9220
rect 10893 9276 10957 9280
rect 10893 9220 10897 9276
rect 10897 9220 10953 9276
rect 10953 9220 10957 9276
rect 10893 9216 10957 9220
rect 10973 9276 11037 9280
rect 10973 9220 10977 9276
rect 10977 9220 11033 9276
rect 11033 9220 11037 9276
rect 10973 9216 11037 9220
rect 11053 9276 11117 9280
rect 11053 9220 11057 9276
rect 11057 9220 11113 9276
rect 11113 9220 11117 9276
rect 11053 9216 11117 9220
rect 3417 8732 3481 8736
rect 3417 8676 3421 8732
rect 3421 8676 3477 8732
rect 3477 8676 3481 8732
rect 3417 8672 3481 8676
rect 3497 8732 3561 8736
rect 3497 8676 3501 8732
rect 3501 8676 3557 8732
rect 3557 8676 3561 8732
rect 3497 8672 3561 8676
rect 3577 8732 3641 8736
rect 3577 8676 3581 8732
rect 3581 8676 3637 8732
rect 3637 8676 3641 8732
rect 3577 8672 3641 8676
rect 3657 8732 3721 8736
rect 3657 8676 3661 8732
rect 3661 8676 3717 8732
rect 3717 8676 3721 8732
rect 3657 8672 3721 8676
rect 8348 8732 8412 8736
rect 8348 8676 8352 8732
rect 8352 8676 8408 8732
rect 8408 8676 8412 8732
rect 8348 8672 8412 8676
rect 8428 8732 8492 8736
rect 8428 8676 8432 8732
rect 8432 8676 8488 8732
rect 8488 8676 8492 8732
rect 8428 8672 8492 8676
rect 8508 8732 8572 8736
rect 8508 8676 8512 8732
rect 8512 8676 8568 8732
rect 8568 8676 8572 8732
rect 8508 8672 8572 8676
rect 8588 8732 8652 8736
rect 8588 8676 8592 8732
rect 8592 8676 8648 8732
rect 8648 8676 8652 8732
rect 8588 8672 8652 8676
rect 13278 8732 13342 8736
rect 13278 8676 13282 8732
rect 13282 8676 13338 8732
rect 13338 8676 13342 8732
rect 13278 8672 13342 8676
rect 13358 8732 13422 8736
rect 13358 8676 13362 8732
rect 13362 8676 13418 8732
rect 13418 8676 13422 8732
rect 13358 8672 13422 8676
rect 13438 8732 13502 8736
rect 13438 8676 13442 8732
rect 13442 8676 13498 8732
rect 13498 8676 13502 8732
rect 13438 8672 13502 8676
rect 13518 8732 13582 8736
rect 13518 8676 13522 8732
rect 13522 8676 13578 8732
rect 13578 8676 13582 8732
rect 13518 8672 13582 8676
rect 5882 8188 5946 8192
rect 5882 8132 5886 8188
rect 5886 8132 5942 8188
rect 5942 8132 5946 8188
rect 5882 8128 5946 8132
rect 5962 8188 6026 8192
rect 5962 8132 5966 8188
rect 5966 8132 6022 8188
rect 6022 8132 6026 8188
rect 5962 8128 6026 8132
rect 6042 8188 6106 8192
rect 6042 8132 6046 8188
rect 6046 8132 6102 8188
rect 6102 8132 6106 8188
rect 6042 8128 6106 8132
rect 6122 8188 6186 8192
rect 6122 8132 6126 8188
rect 6126 8132 6182 8188
rect 6182 8132 6186 8188
rect 6122 8128 6186 8132
rect 10813 8188 10877 8192
rect 10813 8132 10817 8188
rect 10817 8132 10873 8188
rect 10873 8132 10877 8188
rect 10813 8128 10877 8132
rect 10893 8188 10957 8192
rect 10893 8132 10897 8188
rect 10897 8132 10953 8188
rect 10953 8132 10957 8188
rect 10893 8128 10957 8132
rect 10973 8188 11037 8192
rect 10973 8132 10977 8188
rect 10977 8132 11033 8188
rect 11033 8132 11037 8188
rect 10973 8128 11037 8132
rect 11053 8188 11117 8192
rect 11053 8132 11057 8188
rect 11057 8132 11113 8188
rect 11113 8132 11117 8188
rect 11053 8128 11117 8132
rect 3417 7644 3481 7648
rect 3417 7588 3421 7644
rect 3421 7588 3477 7644
rect 3477 7588 3481 7644
rect 3417 7584 3481 7588
rect 3497 7644 3561 7648
rect 3497 7588 3501 7644
rect 3501 7588 3557 7644
rect 3557 7588 3561 7644
rect 3497 7584 3561 7588
rect 3577 7644 3641 7648
rect 3577 7588 3581 7644
rect 3581 7588 3637 7644
rect 3637 7588 3641 7644
rect 3577 7584 3641 7588
rect 3657 7644 3721 7648
rect 3657 7588 3661 7644
rect 3661 7588 3717 7644
rect 3717 7588 3721 7644
rect 3657 7584 3721 7588
rect 8348 7644 8412 7648
rect 8348 7588 8352 7644
rect 8352 7588 8408 7644
rect 8408 7588 8412 7644
rect 8348 7584 8412 7588
rect 8428 7644 8492 7648
rect 8428 7588 8432 7644
rect 8432 7588 8488 7644
rect 8488 7588 8492 7644
rect 8428 7584 8492 7588
rect 8508 7644 8572 7648
rect 8508 7588 8512 7644
rect 8512 7588 8568 7644
rect 8568 7588 8572 7644
rect 8508 7584 8572 7588
rect 8588 7644 8652 7648
rect 8588 7588 8592 7644
rect 8592 7588 8648 7644
rect 8648 7588 8652 7644
rect 8588 7584 8652 7588
rect 13278 7644 13342 7648
rect 13278 7588 13282 7644
rect 13282 7588 13338 7644
rect 13338 7588 13342 7644
rect 13278 7584 13342 7588
rect 13358 7644 13422 7648
rect 13358 7588 13362 7644
rect 13362 7588 13418 7644
rect 13418 7588 13422 7644
rect 13358 7584 13422 7588
rect 13438 7644 13502 7648
rect 13438 7588 13442 7644
rect 13442 7588 13498 7644
rect 13498 7588 13502 7644
rect 13438 7584 13502 7588
rect 13518 7644 13582 7648
rect 13518 7588 13522 7644
rect 13522 7588 13578 7644
rect 13578 7588 13582 7644
rect 13518 7584 13582 7588
rect 5882 7100 5946 7104
rect 5882 7044 5886 7100
rect 5886 7044 5942 7100
rect 5942 7044 5946 7100
rect 5882 7040 5946 7044
rect 5962 7100 6026 7104
rect 5962 7044 5966 7100
rect 5966 7044 6022 7100
rect 6022 7044 6026 7100
rect 5962 7040 6026 7044
rect 6042 7100 6106 7104
rect 6042 7044 6046 7100
rect 6046 7044 6102 7100
rect 6102 7044 6106 7100
rect 6042 7040 6106 7044
rect 6122 7100 6186 7104
rect 6122 7044 6126 7100
rect 6126 7044 6182 7100
rect 6182 7044 6186 7100
rect 6122 7040 6186 7044
rect 10813 7100 10877 7104
rect 10813 7044 10817 7100
rect 10817 7044 10873 7100
rect 10873 7044 10877 7100
rect 10813 7040 10877 7044
rect 10893 7100 10957 7104
rect 10893 7044 10897 7100
rect 10897 7044 10953 7100
rect 10953 7044 10957 7100
rect 10893 7040 10957 7044
rect 10973 7100 11037 7104
rect 10973 7044 10977 7100
rect 10977 7044 11033 7100
rect 11033 7044 11037 7100
rect 10973 7040 11037 7044
rect 11053 7100 11117 7104
rect 11053 7044 11057 7100
rect 11057 7044 11113 7100
rect 11113 7044 11117 7100
rect 11053 7040 11117 7044
rect 3417 6556 3481 6560
rect 3417 6500 3421 6556
rect 3421 6500 3477 6556
rect 3477 6500 3481 6556
rect 3417 6496 3481 6500
rect 3497 6556 3561 6560
rect 3497 6500 3501 6556
rect 3501 6500 3557 6556
rect 3557 6500 3561 6556
rect 3497 6496 3561 6500
rect 3577 6556 3641 6560
rect 3577 6500 3581 6556
rect 3581 6500 3637 6556
rect 3637 6500 3641 6556
rect 3577 6496 3641 6500
rect 3657 6556 3721 6560
rect 3657 6500 3661 6556
rect 3661 6500 3717 6556
rect 3717 6500 3721 6556
rect 3657 6496 3721 6500
rect 8348 6556 8412 6560
rect 8348 6500 8352 6556
rect 8352 6500 8408 6556
rect 8408 6500 8412 6556
rect 8348 6496 8412 6500
rect 8428 6556 8492 6560
rect 8428 6500 8432 6556
rect 8432 6500 8488 6556
rect 8488 6500 8492 6556
rect 8428 6496 8492 6500
rect 8508 6556 8572 6560
rect 8508 6500 8512 6556
rect 8512 6500 8568 6556
rect 8568 6500 8572 6556
rect 8508 6496 8572 6500
rect 8588 6556 8652 6560
rect 8588 6500 8592 6556
rect 8592 6500 8648 6556
rect 8648 6500 8652 6556
rect 8588 6496 8652 6500
rect 13278 6556 13342 6560
rect 13278 6500 13282 6556
rect 13282 6500 13338 6556
rect 13338 6500 13342 6556
rect 13278 6496 13342 6500
rect 13358 6556 13422 6560
rect 13358 6500 13362 6556
rect 13362 6500 13418 6556
rect 13418 6500 13422 6556
rect 13358 6496 13422 6500
rect 13438 6556 13502 6560
rect 13438 6500 13442 6556
rect 13442 6500 13498 6556
rect 13498 6500 13502 6556
rect 13438 6496 13502 6500
rect 13518 6556 13582 6560
rect 13518 6500 13522 6556
rect 13522 6500 13578 6556
rect 13578 6500 13582 6556
rect 13518 6496 13582 6500
rect 5882 6012 5946 6016
rect 5882 5956 5886 6012
rect 5886 5956 5942 6012
rect 5942 5956 5946 6012
rect 5882 5952 5946 5956
rect 5962 6012 6026 6016
rect 5962 5956 5966 6012
rect 5966 5956 6022 6012
rect 6022 5956 6026 6012
rect 5962 5952 6026 5956
rect 6042 6012 6106 6016
rect 6042 5956 6046 6012
rect 6046 5956 6102 6012
rect 6102 5956 6106 6012
rect 6042 5952 6106 5956
rect 6122 6012 6186 6016
rect 6122 5956 6126 6012
rect 6126 5956 6182 6012
rect 6182 5956 6186 6012
rect 6122 5952 6186 5956
rect 10813 6012 10877 6016
rect 10813 5956 10817 6012
rect 10817 5956 10873 6012
rect 10873 5956 10877 6012
rect 10813 5952 10877 5956
rect 10893 6012 10957 6016
rect 10893 5956 10897 6012
rect 10897 5956 10953 6012
rect 10953 5956 10957 6012
rect 10893 5952 10957 5956
rect 10973 6012 11037 6016
rect 10973 5956 10977 6012
rect 10977 5956 11033 6012
rect 11033 5956 11037 6012
rect 10973 5952 11037 5956
rect 11053 6012 11117 6016
rect 11053 5956 11057 6012
rect 11057 5956 11113 6012
rect 11113 5956 11117 6012
rect 11053 5952 11117 5956
rect 3417 5468 3481 5472
rect 3417 5412 3421 5468
rect 3421 5412 3477 5468
rect 3477 5412 3481 5468
rect 3417 5408 3481 5412
rect 3497 5468 3561 5472
rect 3497 5412 3501 5468
rect 3501 5412 3557 5468
rect 3557 5412 3561 5468
rect 3497 5408 3561 5412
rect 3577 5468 3641 5472
rect 3577 5412 3581 5468
rect 3581 5412 3637 5468
rect 3637 5412 3641 5468
rect 3577 5408 3641 5412
rect 3657 5468 3721 5472
rect 3657 5412 3661 5468
rect 3661 5412 3717 5468
rect 3717 5412 3721 5468
rect 3657 5408 3721 5412
rect 8348 5468 8412 5472
rect 8348 5412 8352 5468
rect 8352 5412 8408 5468
rect 8408 5412 8412 5468
rect 8348 5408 8412 5412
rect 8428 5468 8492 5472
rect 8428 5412 8432 5468
rect 8432 5412 8488 5468
rect 8488 5412 8492 5468
rect 8428 5408 8492 5412
rect 8508 5468 8572 5472
rect 8508 5412 8512 5468
rect 8512 5412 8568 5468
rect 8568 5412 8572 5468
rect 8508 5408 8572 5412
rect 8588 5468 8652 5472
rect 8588 5412 8592 5468
rect 8592 5412 8648 5468
rect 8648 5412 8652 5468
rect 8588 5408 8652 5412
rect 13278 5468 13342 5472
rect 13278 5412 13282 5468
rect 13282 5412 13338 5468
rect 13338 5412 13342 5468
rect 13278 5408 13342 5412
rect 13358 5468 13422 5472
rect 13358 5412 13362 5468
rect 13362 5412 13418 5468
rect 13418 5412 13422 5468
rect 13358 5408 13422 5412
rect 13438 5468 13502 5472
rect 13438 5412 13442 5468
rect 13442 5412 13498 5468
rect 13498 5412 13502 5468
rect 13438 5408 13502 5412
rect 13518 5468 13582 5472
rect 13518 5412 13522 5468
rect 13522 5412 13578 5468
rect 13578 5412 13582 5468
rect 13518 5408 13582 5412
rect 5882 4924 5946 4928
rect 5882 4868 5886 4924
rect 5886 4868 5942 4924
rect 5942 4868 5946 4924
rect 5882 4864 5946 4868
rect 5962 4924 6026 4928
rect 5962 4868 5966 4924
rect 5966 4868 6022 4924
rect 6022 4868 6026 4924
rect 5962 4864 6026 4868
rect 6042 4924 6106 4928
rect 6042 4868 6046 4924
rect 6046 4868 6102 4924
rect 6102 4868 6106 4924
rect 6042 4864 6106 4868
rect 6122 4924 6186 4928
rect 6122 4868 6126 4924
rect 6126 4868 6182 4924
rect 6182 4868 6186 4924
rect 6122 4864 6186 4868
rect 10813 4924 10877 4928
rect 10813 4868 10817 4924
rect 10817 4868 10873 4924
rect 10873 4868 10877 4924
rect 10813 4864 10877 4868
rect 10893 4924 10957 4928
rect 10893 4868 10897 4924
rect 10897 4868 10953 4924
rect 10953 4868 10957 4924
rect 10893 4864 10957 4868
rect 10973 4924 11037 4928
rect 10973 4868 10977 4924
rect 10977 4868 11033 4924
rect 11033 4868 11037 4924
rect 10973 4864 11037 4868
rect 11053 4924 11117 4928
rect 11053 4868 11057 4924
rect 11057 4868 11113 4924
rect 11113 4868 11117 4924
rect 11053 4864 11117 4868
rect 3417 4380 3481 4384
rect 3417 4324 3421 4380
rect 3421 4324 3477 4380
rect 3477 4324 3481 4380
rect 3417 4320 3481 4324
rect 3497 4380 3561 4384
rect 3497 4324 3501 4380
rect 3501 4324 3557 4380
rect 3557 4324 3561 4380
rect 3497 4320 3561 4324
rect 3577 4380 3641 4384
rect 3577 4324 3581 4380
rect 3581 4324 3637 4380
rect 3637 4324 3641 4380
rect 3577 4320 3641 4324
rect 3657 4380 3721 4384
rect 3657 4324 3661 4380
rect 3661 4324 3717 4380
rect 3717 4324 3721 4380
rect 3657 4320 3721 4324
rect 8348 4380 8412 4384
rect 8348 4324 8352 4380
rect 8352 4324 8408 4380
rect 8408 4324 8412 4380
rect 8348 4320 8412 4324
rect 8428 4380 8492 4384
rect 8428 4324 8432 4380
rect 8432 4324 8488 4380
rect 8488 4324 8492 4380
rect 8428 4320 8492 4324
rect 8508 4380 8572 4384
rect 8508 4324 8512 4380
rect 8512 4324 8568 4380
rect 8568 4324 8572 4380
rect 8508 4320 8572 4324
rect 8588 4380 8652 4384
rect 8588 4324 8592 4380
rect 8592 4324 8648 4380
rect 8648 4324 8652 4380
rect 8588 4320 8652 4324
rect 13278 4380 13342 4384
rect 13278 4324 13282 4380
rect 13282 4324 13338 4380
rect 13338 4324 13342 4380
rect 13278 4320 13342 4324
rect 13358 4380 13422 4384
rect 13358 4324 13362 4380
rect 13362 4324 13418 4380
rect 13418 4324 13422 4380
rect 13358 4320 13422 4324
rect 13438 4380 13502 4384
rect 13438 4324 13442 4380
rect 13442 4324 13498 4380
rect 13498 4324 13502 4380
rect 13438 4320 13502 4324
rect 13518 4380 13582 4384
rect 13518 4324 13522 4380
rect 13522 4324 13578 4380
rect 13578 4324 13582 4380
rect 13518 4320 13582 4324
rect 5882 3836 5946 3840
rect 5882 3780 5886 3836
rect 5886 3780 5942 3836
rect 5942 3780 5946 3836
rect 5882 3776 5946 3780
rect 5962 3836 6026 3840
rect 5962 3780 5966 3836
rect 5966 3780 6022 3836
rect 6022 3780 6026 3836
rect 5962 3776 6026 3780
rect 6042 3836 6106 3840
rect 6042 3780 6046 3836
rect 6046 3780 6102 3836
rect 6102 3780 6106 3836
rect 6042 3776 6106 3780
rect 6122 3836 6186 3840
rect 6122 3780 6126 3836
rect 6126 3780 6182 3836
rect 6182 3780 6186 3836
rect 6122 3776 6186 3780
rect 10813 3836 10877 3840
rect 10813 3780 10817 3836
rect 10817 3780 10873 3836
rect 10873 3780 10877 3836
rect 10813 3776 10877 3780
rect 10893 3836 10957 3840
rect 10893 3780 10897 3836
rect 10897 3780 10953 3836
rect 10953 3780 10957 3836
rect 10893 3776 10957 3780
rect 10973 3836 11037 3840
rect 10973 3780 10977 3836
rect 10977 3780 11033 3836
rect 11033 3780 11037 3836
rect 10973 3776 11037 3780
rect 11053 3836 11117 3840
rect 11053 3780 11057 3836
rect 11057 3780 11113 3836
rect 11113 3780 11117 3836
rect 11053 3776 11117 3780
rect 3417 3292 3481 3296
rect 3417 3236 3421 3292
rect 3421 3236 3477 3292
rect 3477 3236 3481 3292
rect 3417 3232 3481 3236
rect 3497 3292 3561 3296
rect 3497 3236 3501 3292
rect 3501 3236 3557 3292
rect 3557 3236 3561 3292
rect 3497 3232 3561 3236
rect 3577 3292 3641 3296
rect 3577 3236 3581 3292
rect 3581 3236 3637 3292
rect 3637 3236 3641 3292
rect 3577 3232 3641 3236
rect 3657 3292 3721 3296
rect 3657 3236 3661 3292
rect 3661 3236 3717 3292
rect 3717 3236 3721 3292
rect 3657 3232 3721 3236
rect 8348 3292 8412 3296
rect 8348 3236 8352 3292
rect 8352 3236 8408 3292
rect 8408 3236 8412 3292
rect 8348 3232 8412 3236
rect 8428 3292 8492 3296
rect 8428 3236 8432 3292
rect 8432 3236 8488 3292
rect 8488 3236 8492 3292
rect 8428 3232 8492 3236
rect 8508 3292 8572 3296
rect 8508 3236 8512 3292
rect 8512 3236 8568 3292
rect 8568 3236 8572 3292
rect 8508 3232 8572 3236
rect 8588 3292 8652 3296
rect 8588 3236 8592 3292
rect 8592 3236 8648 3292
rect 8648 3236 8652 3292
rect 8588 3232 8652 3236
rect 13278 3292 13342 3296
rect 13278 3236 13282 3292
rect 13282 3236 13338 3292
rect 13338 3236 13342 3292
rect 13278 3232 13342 3236
rect 13358 3292 13422 3296
rect 13358 3236 13362 3292
rect 13362 3236 13418 3292
rect 13418 3236 13422 3292
rect 13358 3232 13422 3236
rect 13438 3292 13502 3296
rect 13438 3236 13442 3292
rect 13442 3236 13498 3292
rect 13498 3236 13502 3292
rect 13438 3232 13502 3236
rect 13518 3292 13582 3296
rect 13518 3236 13522 3292
rect 13522 3236 13578 3292
rect 13578 3236 13582 3292
rect 13518 3232 13582 3236
rect 5882 2748 5946 2752
rect 5882 2692 5886 2748
rect 5886 2692 5942 2748
rect 5942 2692 5946 2748
rect 5882 2688 5946 2692
rect 5962 2748 6026 2752
rect 5962 2692 5966 2748
rect 5966 2692 6022 2748
rect 6022 2692 6026 2748
rect 5962 2688 6026 2692
rect 6042 2748 6106 2752
rect 6042 2692 6046 2748
rect 6046 2692 6102 2748
rect 6102 2692 6106 2748
rect 6042 2688 6106 2692
rect 6122 2748 6186 2752
rect 6122 2692 6126 2748
rect 6126 2692 6182 2748
rect 6182 2692 6186 2748
rect 6122 2688 6186 2692
rect 10813 2748 10877 2752
rect 10813 2692 10817 2748
rect 10817 2692 10873 2748
rect 10873 2692 10877 2748
rect 10813 2688 10877 2692
rect 10893 2748 10957 2752
rect 10893 2692 10897 2748
rect 10897 2692 10953 2748
rect 10953 2692 10957 2748
rect 10893 2688 10957 2692
rect 10973 2748 11037 2752
rect 10973 2692 10977 2748
rect 10977 2692 11033 2748
rect 11033 2692 11037 2748
rect 10973 2688 11037 2692
rect 11053 2748 11117 2752
rect 11053 2692 11057 2748
rect 11057 2692 11113 2748
rect 11113 2692 11117 2748
rect 11053 2688 11117 2692
rect 3417 2204 3481 2208
rect 3417 2148 3421 2204
rect 3421 2148 3477 2204
rect 3477 2148 3481 2204
rect 3417 2144 3481 2148
rect 3497 2204 3561 2208
rect 3497 2148 3501 2204
rect 3501 2148 3557 2204
rect 3557 2148 3561 2204
rect 3497 2144 3561 2148
rect 3577 2204 3641 2208
rect 3577 2148 3581 2204
rect 3581 2148 3637 2204
rect 3637 2148 3641 2204
rect 3577 2144 3641 2148
rect 3657 2204 3721 2208
rect 3657 2148 3661 2204
rect 3661 2148 3717 2204
rect 3717 2148 3721 2204
rect 3657 2144 3721 2148
rect 8348 2204 8412 2208
rect 8348 2148 8352 2204
rect 8352 2148 8408 2204
rect 8408 2148 8412 2204
rect 8348 2144 8412 2148
rect 8428 2204 8492 2208
rect 8428 2148 8432 2204
rect 8432 2148 8488 2204
rect 8488 2148 8492 2204
rect 8428 2144 8492 2148
rect 8508 2204 8572 2208
rect 8508 2148 8512 2204
rect 8512 2148 8568 2204
rect 8568 2148 8572 2204
rect 8508 2144 8572 2148
rect 8588 2204 8652 2208
rect 8588 2148 8592 2204
rect 8592 2148 8648 2204
rect 8648 2148 8652 2204
rect 8588 2144 8652 2148
rect 13278 2204 13342 2208
rect 13278 2148 13282 2204
rect 13282 2148 13338 2204
rect 13338 2148 13342 2204
rect 13278 2144 13342 2148
rect 13358 2204 13422 2208
rect 13358 2148 13362 2204
rect 13362 2148 13418 2204
rect 13418 2148 13422 2204
rect 13358 2144 13422 2148
rect 13438 2204 13502 2208
rect 13438 2148 13442 2204
rect 13442 2148 13498 2204
rect 13498 2148 13502 2204
rect 13438 2144 13502 2148
rect 13518 2204 13582 2208
rect 13518 2148 13522 2204
rect 13522 2148 13578 2204
rect 13578 2148 13582 2204
rect 13518 2144 13582 2148
<< metal4 >>
rect 3409 17440 3729 17456
rect 3409 17376 3417 17440
rect 3481 17376 3497 17440
rect 3561 17376 3577 17440
rect 3641 17376 3657 17440
rect 3721 17376 3729 17440
rect 3409 16352 3729 17376
rect 3409 16288 3417 16352
rect 3481 16288 3497 16352
rect 3561 16288 3577 16352
rect 3641 16288 3657 16352
rect 3721 16288 3729 16352
rect 3409 15264 3729 16288
rect 3409 15200 3417 15264
rect 3481 15200 3497 15264
rect 3561 15200 3577 15264
rect 3641 15200 3657 15264
rect 3721 15200 3729 15264
rect 3409 14176 3729 15200
rect 3409 14112 3417 14176
rect 3481 14112 3497 14176
rect 3561 14112 3577 14176
rect 3641 14112 3657 14176
rect 3721 14112 3729 14176
rect 3409 13088 3729 14112
rect 3409 13024 3417 13088
rect 3481 13024 3497 13088
rect 3561 13024 3577 13088
rect 3641 13024 3657 13088
rect 3721 13024 3729 13088
rect 3409 12000 3729 13024
rect 3409 11936 3417 12000
rect 3481 11936 3497 12000
rect 3561 11936 3577 12000
rect 3641 11936 3657 12000
rect 3721 11936 3729 12000
rect 3409 10912 3729 11936
rect 3409 10848 3417 10912
rect 3481 10848 3497 10912
rect 3561 10848 3577 10912
rect 3641 10848 3657 10912
rect 3721 10848 3729 10912
rect 3409 9824 3729 10848
rect 3409 9760 3417 9824
rect 3481 9760 3497 9824
rect 3561 9760 3577 9824
rect 3641 9760 3657 9824
rect 3721 9760 3729 9824
rect 3409 8736 3729 9760
rect 3409 8672 3417 8736
rect 3481 8672 3497 8736
rect 3561 8672 3577 8736
rect 3641 8672 3657 8736
rect 3721 8672 3729 8736
rect 3409 7648 3729 8672
rect 3409 7584 3417 7648
rect 3481 7584 3497 7648
rect 3561 7584 3577 7648
rect 3641 7584 3657 7648
rect 3721 7584 3729 7648
rect 3409 6560 3729 7584
rect 3409 6496 3417 6560
rect 3481 6496 3497 6560
rect 3561 6496 3577 6560
rect 3641 6496 3657 6560
rect 3721 6496 3729 6560
rect 3409 5472 3729 6496
rect 3409 5408 3417 5472
rect 3481 5408 3497 5472
rect 3561 5408 3577 5472
rect 3641 5408 3657 5472
rect 3721 5408 3729 5472
rect 3409 4384 3729 5408
rect 3409 4320 3417 4384
rect 3481 4320 3497 4384
rect 3561 4320 3577 4384
rect 3641 4320 3657 4384
rect 3721 4320 3729 4384
rect 3409 3296 3729 4320
rect 3409 3232 3417 3296
rect 3481 3232 3497 3296
rect 3561 3232 3577 3296
rect 3641 3232 3657 3296
rect 3721 3232 3729 3296
rect 3409 2208 3729 3232
rect 3409 2144 3417 2208
rect 3481 2144 3497 2208
rect 3561 2144 3577 2208
rect 3641 2144 3657 2208
rect 3721 2144 3729 2208
rect 3409 2128 3729 2144
rect 5874 16896 6195 17456
rect 5874 16832 5882 16896
rect 5946 16832 5962 16896
rect 6026 16832 6042 16896
rect 6106 16832 6122 16896
rect 6186 16832 6195 16896
rect 5874 15808 6195 16832
rect 5874 15744 5882 15808
rect 5946 15744 5962 15808
rect 6026 15744 6042 15808
rect 6106 15744 6122 15808
rect 6186 15744 6195 15808
rect 5874 14720 6195 15744
rect 5874 14656 5882 14720
rect 5946 14656 5962 14720
rect 6026 14656 6042 14720
rect 6106 14656 6122 14720
rect 6186 14656 6195 14720
rect 5874 13632 6195 14656
rect 5874 13568 5882 13632
rect 5946 13568 5962 13632
rect 6026 13568 6042 13632
rect 6106 13568 6122 13632
rect 6186 13568 6195 13632
rect 5874 12544 6195 13568
rect 5874 12480 5882 12544
rect 5946 12480 5962 12544
rect 6026 12480 6042 12544
rect 6106 12480 6122 12544
rect 6186 12480 6195 12544
rect 5874 11456 6195 12480
rect 5874 11392 5882 11456
rect 5946 11392 5962 11456
rect 6026 11392 6042 11456
rect 6106 11392 6122 11456
rect 6186 11392 6195 11456
rect 5874 10368 6195 11392
rect 5874 10304 5882 10368
rect 5946 10304 5962 10368
rect 6026 10304 6042 10368
rect 6106 10304 6122 10368
rect 6186 10304 6195 10368
rect 5874 9280 6195 10304
rect 5874 9216 5882 9280
rect 5946 9216 5962 9280
rect 6026 9216 6042 9280
rect 6106 9216 6122 9280
rect 6186 9216 6195 9280
rect 5874 8192 6195 9216
rect 5874 8128 5882 8192
rect 5946 8128 5962 8192
rect 6026 8128 6042 8192
rect 6106 8128 6122 8192
rect 6186 8128 6195 8192
rect 5874 7104 6195 8128
rect 5874 7040 5882 7104
rect 5946 7040 5962 7104
rect 6026 7040 6042 7104
rect 6106 7040 6122 7104
rect 6186 7040 6195 7104
rect 5874 6016 6195 7040
rect 5874 5952 5882 6016
rect 5946 5952 5962 6016
rect 6026 5952 6042 6016
rect 6106 5952 6122 6016
rect 6186 5952 6195 6016
rect 5874 4928 6195 5952
rect 5874 4864 5882 4928
rect 5946 4864 5962 4928
rect 6026 4864 6042 4928
rect 6106 4864 6122 4928
rect 6186 4864 6195 4928
rect 5874 3840 6195 4864
rect 5874 3776 5882 3840
rect 5946 3776 5962 3840
rect 6026 3776 6042 3840
rect 6106 3776 6122 3840
rect 6186 3776 6195 3840
rect 5874 2752 6195 3776
rect 5874 2688 5882 2752
rect 5946 2688 5962 2752
rect 6026 2688 6042 2752
rect 6106 2688 6122 2752
rect 6186 2688 6195 2752
rect 5874 2128 6195 2688
rect 8340 17440 8660 17456
rect 8340 17376 8348 17440
rect 8412 17376 8428 17440
rect 8492 17376 8508 17440
rect 8572 17376 8588 17440
rect 8652 17376 8660 17440
rect 8340 16352 8660 17376
rect 8340 16288 8348 16352
rect 8412 16288 8428 16352
rect 8492 16288 8508 16352
rect 8572 16288 8588 16352
rect 8652 16288 8660 16352
rect 8340 15264 8660 16288
rect 8340 15200 8348 15264
rect 8412 15200 8428 15264
rect 8492 15200 8508 15264
rect 8572 15200 8588 15264
rect 8652 15200 8660 15264
rect 8340 14176 8660 15200
rect 8340 14112 8348 14176
rect 8412 14112 8428 14176
rect 8492 14112 8508 14176
rect 8572 14112 8588 14176
rect 8652 14112 8660 14176
rect 8340 13088 8660 14112
rect 8340 13024 8348 13088
rect 8412 13024 8428 13088
rect 8492 13024 8508 13088
rect 8572 13024 8588 13088
rect 8652 13024 8660 13088
rect 8340 12000 8660 13024
rect 8340 11936 8348 12000
rect 8412 11936 8428 12000
rect 8492 11936 8508 12000
rect 8572 11936 8588 12000
rect 8652 11936 8660 12000
rect 8340 10912 8660 11936
rect 8340 10848 8348 10912
rect 8412 10848 8428 10912
rect 8492 10848 8508 10912
rect 8572 10848 8588 10912
rect 8652 10848 8660 10912
rect 8340 9824 8660 10848
rect 8340 9760 8348 9824
rect 8412 9760 8428 9824
rect 8492 9760 8508 9824
rect 8572 9760 8588 9824
rect 8652 9760 8660 9824
rect 8340 8736 8660 9760
rect 8340 8672 8348 8736
rect 8412 8672 8428 8736
rect 8492 8672 8508 8736
rect 8572 8672 8588 8736
rect 8652 8672 8660 8736
rect 8340 7648 8660 8672
rect 8340 7584 8348 7648
rect 8412 7584 8428 7648
rect 8492 7584 8508 7648
rect 8572 7584 8588 7648
rect 8652 7584 8660 7648
rect 8340 6560 8660 7584
rect 8340 6496 8348 6560
rect 8412 6496 8428 6560
rect 8492 6496 8508 6560
rect 8572 6496 8588 6560
rect 8652 6496 8660 6560
rect 8340 5472 8660 6496
rect 8340 5408 8348 5472
rect 8412 5408 8428 5472
rect 8492 5408 8508 5472
rect 8572 5408 8588 5472
rect 8652 5408 8660 5472
rect 8340 4384 8660 5408
rect 8340 4320 8348 4384
rect 8412 4320 8428 4384
rect 8492 4320 8508 4384
rect 8572 4320 8588 4384
rect 8652 4320 8660 4384
rect 8340 3296 8660 4320
rect 8340 3232 8348 3296
rect 8412 3232 8428 3296
rect 8492 3232 8508 3296
rect 8572 3232 8588 3296
rect 8652 3232 8660 3296
rect 8340 2208 8660 3232
rect 8340 2144 8348 2208
rect 8412 2144 8428 2208
rect 8492 2144 8508 2208
rect 8572 2144 8588 2208
rect 8652 2144 8660 2208
rect 8340 2128 8660 2144
rect 10805 16896 11125 17456
rect 10805 16832 10813 16896
rect 10877 16832 10893 16896
rect 10957 16832 10973 16896
rect 11037 16832 11053 16896
rect 11117 16832 11125 16896
rect 10805 15808 11125 16832
rect 10805 15744 10813 15808
rect 10877 15744 10893 15808
rect 10957 15744 10973 15808
rect 11037 15744 11053 15808
rect 11117 15744 11125 15808
rect 10805 14720 11125 15744
rect 10805 14656 10813 14720
rect 10877 14656 10893 14720
rect 10957 14656 10973 14720
rect 11037 14656 11053 14720
rect 11117 14656 11125 14720
rect 10805 13632 11125 14656
rect 10805 13568 10813 13632
rect 10877 13568 10893 13632
rect 10957 13568 10973 13632
rect 11037 13568 11053 13632
rect 11117 13568 11125 13632
rect 10805 12544 11125 13568
rect 10805 12480 10813 12544
rect 10877 12480 10893 12544
rect 10957 12480 10973 12544
rect 11037 12480 11053 12544
rect 11117 12480 11125 12544
rect 10805 11456 11125 12480
rect 10805 11392 10813 11456
rect 10877 11392 10893 11456
rect 10957 11392 10973 11456
rect 11037 11392 11053 11456
rect 11117 11392 11125 11456
rect 10805 10368 11125 11392
rect 10805 10304 10813 10368
rect 10877 10304 10893 10368
rect 10957 10304 10973 10368
rect 11037 10304 11053 10368
rect 11117 10304 11125 10368
rect 10805 9280 11125 10304
rect 10805 9216 10813 9280
rect 10877 9216 10893 9280
rect 10957 9216 10973 9280
rect 11037 9216 11053 9280
rect 11117 9216 11125 9280
rect 10805 8192 11125 9216
rect 10805 8128 10813 8192
rect 10877 8128 10893 8192
rect 10957 8128 10973 8192
rect 11037 8128 11053 8192
rect 11117 8128 11125 8192
rect 10805 7104 11125 8128
rect 10805 7040 10813 7104
rect 10877 7040 10893 7104
rect 10957 7040 10973 7104
rect 11037 7040 11053 7104
rect 11117 7040 11125 7104
rect 10805 6016 11125 7040
rect 10805 5952 10813 6016
rect 10877 5952 10893 6016
rect 10957 5952 10973 6016
rect 11037 5952 11053 6016
rect 11117 5952 11125 6016
rect 10805 4928 11125 5952
rect 10805 4864 10813 4928
rect 10877 4864 10893 4928
rect 10957 4864 10973 4928
rect 11037 4864 11053 4928
rect 11117 4864 11125 4928
rect 10805 3840 11125 4864
rect 10805 3776 10813 3840
rect 10877 3776 10893 3840
rect 10957 3776 10973 3840
rect 11037 3776 11053 3840
rect 11117 3776 11125 3840
rect 10805 2752 11125 3776
rect 10805 2688 10813 2752
rect 10877 2688 10893 2752
rect 10957 2688 10973 2752
rect 11037 2688 11053 2752
rect 11117 2688 11125 2752
rect 10805 2128 11125 2688
rect 13270 17440 13590 17456
rect 13270 17376 13278 17440
rect 13342 17376 13358 17440
rect 13422 17376 13438 17440
rect 13502 17376 13518 17440
rect 13582 17376 13590 17440
rect 13270 16352 13590 17376
rect 13270 16288 13278 16352
rect 13342 16288 13358 16352
rect 13422 16288 13438 16352
rect 13502 16288 13518 16352
rect 13582 16288 13590 16352
rect 13270 15264 13590 16288
rect 13270 15200 13278 15264
rect 13342 15200 13358 15264
rect 13422 15200 13438 15264
rect 13502 15200 13518 15264
rect 13582 15200 13590 15264
rect 13270 14176 13590 15200
rect 13270 14112 13278 14176
rect 13342 14112 13358 14176
rect 13422 14112 13438 14176
rect 13502 14112 13518 14176
rect 13582 14112 13590 14176
rect 13270 13088 13590 14112
rect 13270 13024 13278 13088
rect 13342 13024 13358 13088
rect 13422 13024 13438 13088
rect 13502 13024 13518 13088
rect 13582 13024 13590 13088
rect 13270 12000 13590 13024
rect 13270 11936 13278 12000
rect 13342 11936 13358 12000
rect 13422 11936 13438 12000
rect 13502 11936 13518 12000
rect 13582 11936 13590 12000
rect 13270 10912 13590 11936
rect 13270 10848 13278 10912
rect 13342 10848 13358 10912
rect 13422 10848 13438 10912
rect 13502 10848 13518 10912
rect 13582 10848 13590 10912
rect 13270 9824 13590 10848
rect 13270 9760 13278 9824
rect 13342 9760 13358 9824
rect 13422 9760 13438 9824
rect 13502 9760 13518 9824
rect 13582 9760 13590 9824
rect 13270 8736 13590 9760
rect 13270 8672 13278 8736
rect 13342 8672 13358 8736
rect 13422 8672 13438 8736
rect 13502 8672 13518 8736
rect 13582 8672 13590 8736
rect 13270 7648 13590 8672
rect 13270 7584 13278 7648
rect 13342 7584 13358 7648
rect 13422 7584 13438 7648
rect 13502 7584 13518 7648
rect 13582 7584 13590 7648
rect 13270 6560 13590 7584
rect 13270 6496 13278 6560
rect 13342 6496 13358 6560
rect 13422 6496 13438 6560
rect 13502 6496 13518 6560
rect 13582 6496 13590 6560
rect 13270 5472 13590 6496
rect 13270 5408 13278 5472
rect 13342 5408 13358 5472
rect 13422 5408 13438 5472
rect 13502 5408 13518 5472
rect 13582 5408 13590 5472
rect 13270 4384 13590 5408
rect 13270 4320 13278 4384
rect 13342 4320 13358 4384
rect 13422 4320 13438 4384
rect 13502 4320 13518 4384
rect 13582 4320 13590 4384
rect 13270 3296 13590 4320
rect 13270 3232 13278 3296
rect 13342 3232 13358 3296
rect 13422 3232 13438 3296
rect 13502 3232 13518 3296
rect 13582 3232 13590 3296
rect 13270 2208 13590 3232
rect 13270 2144 13278 2208
rect 13342 2144 13358 2208
rect 13422 2144 13438 2208
rect 13502 2144 13518 2208
rect 13582 2144 13590 2208
rect 13270 2128 13590 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606256979
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606256979
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1606256979
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1606256979
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606256979
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606256979
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1606256979
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606256979
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1606256979
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1606256979
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1606256979
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1606256979
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1606256979
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1606256979
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1606256979
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 15824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 15824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1606256979
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_147
timestamp 1606256979
transform 1 0 14628 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1606256979
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606256979
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606256979
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606256979
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1606256979
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1606256979
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1606256979
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1606256979
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1606256979
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1606256979
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1606256979
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 15824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606256979
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606256979
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606256979
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606256979
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606256979
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _30_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7728 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1606256979
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_76
timestamp 1606256979
transform 1 0 8096 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1606256979
transform 1 0 9844 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_88
timestamp 1606256979
transform 1 0 9200 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_94
timestamp 1606256979
transform 1 0 9752 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_99
timestamp 1606256979
transform 1 0 10212 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_111
timestamp 1606256979
transform 1 0 11316 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1606256979
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1606256979
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 15824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_147
timestamp 1606256979
transform 1 0 14628 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_155
timestamp 1606256979
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606256979
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1606256979
transform 1 0 4876 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606256979
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_32
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_40
timestamp 1606256979
transform 1 0 4784 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1606256979
transform 1 0 5704 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_45
timestamp 1606256979
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_49
timestamp 1606256979
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_54
timestamp 1606256979
transform 1 0 6072 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_62
timestamp 1606256979
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _09_
timestamp 1606256979
transform 1 0 7820 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _11_
timestamp 1606256979
transform 1 0 6992 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1606256979
transform 1 0 8372 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_68
timestamp 1606256979
transform 1 0 7360 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_72
timestamp 1606256979
transform 1 0 7728 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 1606256979
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_83
timestamp 1606256979
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _05_
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1606256979
transform 1 0 10672 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1606256979
transform 1 0 9016 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1606256979
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_97
timestamp 1606256979
transform 1 0 10028 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_103
timestamp 1606256979
transform 1 0 10580 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1606256979
transform 1 0 11868 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_108
timestamp 1606256979
transform 1 0 11040 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_116
timestamp 1606256979
transform 1 0 11776 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1606256979
transform 1 0 12236 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_133
timestamp 1606256979
transform 1 0 13340 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_145
timestamp 1606256979
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606256979
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1606256979
transform 1 0 4784 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1606256979
transform 1 0 3680 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_27
timestamp 1606256979
transform 1 0 3588 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_32
timestamp 1606256979
transform 1 0 4048 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1606256979
transform 1 0 6164 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1606256979
transform 1 0 5612 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_44
timestamp 1606256979
transform 1 0 5152 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_48
timestamp 1606256979
transform 1 0 5520 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1606256979
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606256979
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1606256979
transform 1 0 8280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1606256979
transform 1 0 7360 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1606256979
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_72
timestamp 1606256979
transform 1 0 7728 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_82
timestamp 1606256979
transform 1 0 8648 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _02_
timestamp 1606256979
transform 1 0 10672 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _03_
timestamp 1606256979
transform 1 0 10120 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _04_
timestamp 1606256979
transform 1 0 9568 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _06_
timestamp 1606256979
transform 1 0 9016 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_90
timestamp 1606256979
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_96
timestamp 1606256979
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_102
timestamp 1606256979
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1606256979
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1606256979
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_108
timestamp 1606256979
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1606256979
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1606256979
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1606256979
transform 1 0 12972 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1606256979
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_133
timestamp 1606256979
transform 1 0 13340 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_145
timestamp 1606256979
transform 1 0 14444 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 15824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606256979
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606256979
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1606256979
transform 1 0 4324 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606256979
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_32
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_39
timestamp 1606256979
transform 1 0 4692 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1606256979
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1606256979
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1606256979
transform 1 0 6808 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1606256979
transform 1 0 5152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_43
timestamp 1606256979
transform 1 0 5060 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_48
timestamp 1606256979
transform 1 0 5520 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_60
timestamp 1606256979
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606256979
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606256979
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _10_
timestamp 1606256979
transform 1 0 7360 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1606256979
transform 1 0 7912 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_66
timestamp 1606256979
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_72
timestamp 1606256979
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78
timestamp 1606256979
transform 1 0 8280 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1606256979
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1606256979
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_84
timestamp 1606256979
transform 1 0 8832 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1606256979
transform 1 0 8924 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_103
timestamp 1606256979
transform 1 0 10580 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_97
timestamp 1606256979
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1606256979
transform 1 0 10212 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1606256979
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1606256979
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1606256979
transform 1 0 11500 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_111
timestamp 1606256979
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1606256979
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1606256979
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1606256979
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1606256979
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1606256979
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 15824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 15824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_147
timestamp 1606256979
transform 1 0 14628 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1606256979
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606256979
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606256979
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1606256979
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1606256979
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1606256979
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1606256979
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1606256979
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1606256979
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1606256979
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1606256979
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1606256979
transform 1 0 2484 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3220 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_29
timestamp 1606256979
transform 1 0 3772 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_41
timestamp 1606256979
transform 1 0 4876 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_53
timestamp 1606256979
transform 1 0 5980 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1606256979
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1606256979
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1606256979
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1606256979
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1606256979
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_147
timestamp 1606256979
transform 1 0 14628 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_155
timestamp 1606256979
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606256979
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606256979
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1606256979
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1606256979
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1606256979
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1606256979
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1606256979
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1606256979
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1606256979
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1606256979
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 15824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1606256979
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1606256979
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1606256979
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1606256979
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606256979
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1606256979
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1606256979
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1606256979
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1606256979
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1606256979
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 15824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_147
timestamp 1606256979
transform 1 0 14628 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1606256979
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1606256979
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1606256979
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1606256979
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1606256979
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1606256979
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1606256979
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 12236 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1606256979
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_117
timestamp 1606256979
transform 1 0 11868 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_133
timestamp 1606256979
transform 1 0 13340 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1606256979
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1606256979
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1606256979
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1606256979
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1606256979
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606256979
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6164 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1606256979
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606256979
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_44
timestamp 1606256979
transform 1 0 5152 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_52
timestamp 1606256979
transform 1 0 5888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7176 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 8188 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 7176 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_75
timestamp 1606256979
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_64
timestamp 1606256979
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_82
timestamp 1606256979
transform 1 0 8648 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _01_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9752 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1606256979
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1606256979
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606256979
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1606256979
transform 1 0 10028 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1606256979
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1606256979
transform 1 0 11132 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1606256979
transform 1 0 12236 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1606256979
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_133
timestamp 1606256979
transform 1 0 13340 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1606256979
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 15824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_147
timestamp 1606256979
transform 1 0 14628 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1606256979
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2760 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_16
timestamp 1606256979
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_21
timestamp 1606256979
transform 1 0 3036 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_33
timestamp 1606256979
transform 1 0 4140 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_45
timestamp 1606256979
transform 1 0 5244 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1606256979
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7544 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7268 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1606256979
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 10212 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 9200 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_86
timestamp 1606256979
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_97
timestamp 1606256979
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_108
timestamp 1606256979
transform 1 0 11040 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606256979
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1606256979
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 15824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_147
timestamp 1606256979
transform 1 0 14628 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1606256979
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1606256979
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606256979
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6256 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_45
timestamp 1606256979
transform 1 0 5244 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_53
timestamp 1606256979
transform 1 0 5980 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7268 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_65
timestamp 1606256979
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_83
timestamp 1606256979
transform 1 0 8740 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1606256979
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_102
timestamp 1606256979
transform 1 0 10488 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_114
timestamp 1606256979
transform 1 0 11592 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_126
timestamp 1606256979
transform 1 0 12696 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_138
timestamp 1606256979
transform 1 0 13800 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 15824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1606256979
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1606256979
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1606256979
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1606256979
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1606256979
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606256979
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7728 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_71
timestamp 1606256979
transform 1 0 7636 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_88
timestamp 1606256979
transform 1 0 9200 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_100
timestamp 1606256979
transform 1 0 10304 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_112
timestamp 1606256979
transform 1 0 11408 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1606256979
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1606256979
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 15824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_147
timestamp 1606256979
transform 1 0 14628 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1606256979
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606256979
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606256979
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5980 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_18_44
timestamp 1606256979
transform 1 0 5152 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_52
timestamp 1606256979
transform 1 0 5888 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 7820 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_82
timestamp 1606256979
transform 1 0 8648 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1606256979
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1606256979
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1606256979
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1606256979
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1606256979
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 15824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2668 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1606256979
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1606256979
transform 1 0 2484 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1606256979
transform 1 0 4784 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1606256979
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1606256979
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_26
timestamp 1606256979
transform 1 0 3496 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1606256979
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_32
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1606256979
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606256979
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_62
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_43
timestamp 1606256979
transform 1 0 5060 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_55
timestamp 1606256979
transform 1 0 6164 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 7544 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_19_79
timestamp 1606256979
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_67
timestamp 1606256979
transform 1 0 7268 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_79
timestamp 1606256979
transform 1 0 8372 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_91
timestamp 1606256979
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_103
timestamp 1606256979
transform 1 0 10580 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606256979
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_115
timestamp 1606256979
transform 1 0 11684 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1606256979
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1606256979
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1606256979
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1606256979
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1606256979
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1606256979
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 15824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_147
timestamp 1606256979
transform 1 0 14628 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1606256979
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1606256979
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4232 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_21_27
timestamp 1606256979
transform 1 0 3588 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_33
timestamp 1606256979
transform 1 0 4140 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_50
timestamp 1606256979
transform 1 0 5704 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_58
timestamp 1606256979
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1606256979
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1606256979
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1606256979
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1606256979
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1606256979
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1606256979
transform 1 0 14996 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 15824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_147
timestamp 1606256979
transform 1 0 14628 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_155
timestamp 1606256979
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1606256979
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606256979
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1606256979
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1606256979
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1606256979
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1606256979
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1606256979
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1606256979
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1606256979
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1606256979
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1606256979
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1606256979
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1606256979
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1606256979
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1606256979
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1606256979
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606256979
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_62
timestamp 1606256979
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _07_
timestamp 1606256979
transform 1 0 7084 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1606256979
transform 1 0 7452 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_81
timestamp 1606256979
transform 1 0 8556 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1606256979
transform 1 0 9200 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_87
timestamp 1606256979
transform 1 0 9108 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_92
timestamp 1606256979
transform 1 0 9568 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_104
timestamp 1606256979
transform 1 0 10672 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_116
timestamp 1606256979
transform 1 0 11776 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1606256979
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1606256979
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp 1606256979
transform 1 0 14628 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1606256979
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1606256979
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1606256979
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _15_
timestamp 1606256979
transform 1 0 4600 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1606256979
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1606256979
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_36
timestamp 1606256979
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1606256979
transform 1 0 5336 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_42
timestamp 1606256979
transform 1 0 4968 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_50
timestamp 1606256979
transform 1 0 5704 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_62
timestamp 1606256979
transform 1 0 6808 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_74
timestamp 1606256979
transform 1 0 7912 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_86
timestamp 1606256979
transform 1 0 9016 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1606256979
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1606256979
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1606256979
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1606256979
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1606256979
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1606256979
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1606256979
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1606256979
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1606256979
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1606256979
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1606256979
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606256979
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1606256979
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1606256979
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1606256979
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1606256979
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1606256979
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1606256979
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1606256979
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_147
timestamp 1606256979
transform 1 0 14628 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1606256979
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1606256979
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1606256979
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1606256979
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1606256979
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1606256979
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1606256979
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1606256979
transform 1 0 3588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1606256979
transform 1 0 4048 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1606256979
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1606256979
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1606256979
transform 1 0 5152 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_56
timestamp 1606256979
transform 1 0 6256 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1606256979
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1606256979
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_63
timestamp 1606256979
transform 1 0 6900 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_75
timestamp 1606256979
transform 1 0 8004 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1606256979
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_87
timestamp 1606256979
transform 1 0 9108 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1606256979
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1606256979
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1606256979
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_106
timestamp 1606256979
transform 1 0 10856 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_118
timestamp 1606256979
transform 1 0 11960 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1606256979
transform 1 0 12604 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1606256979
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1606256979
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1606256979
transform 1 0 13708 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 15824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 15824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1606256979
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_149
timestamp 1606256979
transform 1 0 14812 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1606256979
transform 1 0 15456 0 1 16864
box -38 -48 130 592
<< labels >>
rlabel metal2 s 202 19520 258 20000 6 IO_ISOL_N
port 0 nsew default input
rlabel metal3 s 0 18232 480 18352 6 ccff_head
port 1 nsew default input
rlabel metal3 s 16520 12384 17000 12504 6 ccff_tail
port 2 nsew default tristate
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[0]
port 3 nsew default input
rlabel metal2 s 12898 0 12954 480 6 chany_bottom_in[10]
port 4 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[11]
port 5 nsew default input
rlabel metal2 s 13818 0 13874 480 6 chany_bottom_in[12]
port 6 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[13]
port 7 nsew default input
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_in[14]
port 8 nsew default input
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_in[15]
port 9 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_in[16]
port 10 nsew default input
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_in[17]
port 11 nsew default input
rlabel metal2 s 16302 0 16358 480 6 chany_bottom_in[18]
port 12 nsew default input
rlabel metal2 s 16762 0 16818 480 6 chany_bottom_in[19]
port 13 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[1]
port 14 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[2]
port 15 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[3]
port 16 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[4]
port 17 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_in[5]
port 18 nsew default input
rlabel metal2 s 11242 0 11298 480 6 chany_bottom_in[6]
port 19 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_in[7]
port 20 nsew default input
rlabel metal2 s 12070 0 12126 480 6 chany_bottom_in[8]
port 21 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[9]
port 22 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 23 nsew default tristate
rlabel metal2 s 4434 0 4490 480 6 chany_bottom_out[10]
port 24 nsew default tristate
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_out[11]
port 25 nsew default tristate
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_out[12]
port 26 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[13]
port 27 nsew default tristate
rlabel metal2 s 6090 0 6146 480 6 chany_bottom_out[14]
port 28 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[15]
port 29 nsew default tristate
rlabel metal2 s 7010 0 7066 480 6 chany_bottom_out[16]
port 30 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[17]
port 31 nsew default tristate
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_out[18]
port 32 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_out[19]
port 33 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 34 nsew default tristate
rlabel metal2 s 1030 0 1086 480 6 chany_bottom_out[2]
port 35 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 36 nsew default tristate
rlabel metal2 s 1858 0 1914 480 6 chany_bottom_out[4]
port 37 nsew default tristate
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_out[5]
port 38 nsew default tristate
rlabel metal2 s 2686 0 2742 480 6 chany_bottom_out[6]
port 39 nsew default tristate
rlabel metal2 s 3146 0 3202 480 6 chany_bottom_out[7]
port 40 nsew default tristate
rlabel metal2 s 3606 0 3662 480 6 chany_bottom_out[8]
port 41 nsew default tristate
rlabel metal2 s 3974 0 4030 480 6 chany_bottom_out[9]
port 42 nsew default tristate
rlabel metal2 s 8850 19520 8906 20000 6 chany_top_in[0]
port 43 nsew default input
rlabel metal2 s 12990 19520 13046 20000 6 chany_top_in[10]
port 44 nsew default input
rlabel metal2 s 13450 19520 13506 20000 6 chany_top_in[11]
port 45 nsew default input
rlabel metal2 s 13818 19520 13874 20000 6 chany_top_in[12]
port 46 nsew default input
rlabel metal2 s 14278 19520 14334 20000 6 chany_top_in[13]
port 47 nsew default input
rlabel metal2 s 14646 19520 14702 20000 6 chany_top_in[14]
port 48 nsew default input
rlabel metal2 s 15106 19520 15162 20000 6 chany_top_in[15]
port 49 nsew default input
rlabel metal2 s 15474 19520 15530 20000 6 chany_top_in[16]
port 50 nsew default input
rlabel metal2 s 15934 19520 15990 20000 6 chany_top_in[17]
port 51 nsew default input
rlabel metal2 s 16302 19520 16358 20000 6 chany_top_in[18]
port 52 nsew default input
rlabel metal2 s 16762 19520 16818 20000 6 chany_top_in[19]
port 53 nsew default input
rlabel metal2 s 9310 19520 9366 20000 6 chany_top_in[1]
port 54 nsew default input
rlabel metal2 s 9678 19520 9734 20000 6 chany_top_in[2]
port 55 nsew default input
rlabel metal2 s 10138 19520 10194 20000 6 chany_top_in[3]
port 56 nsew default input
rlabel metal2 s 10506 19520 10562 20000 6 chany_top_in[4]
port 57 nsew default input
rlabel metal2 s 10966 19520 11022 20000 6 chany_top_in[5]
port 58 nsew default input
rlabel metal2 s 11334 19520 11390 20000 6 chany_top_in[6]
port 59 nsew default input
rlabel metal2 s 11794 19520 11850 20000 6 chany_top_in[7]
port 60 nsew default input
rlabel metal2 s 12162 19520 12218 20000 6 chany_top_in[8]
port 61 nsew default input
rlabel metal2 s 12622 19520 12678 20000 6 chany_top_in[9]
port 62 nsew default input
rlabel metal2 s 570 19520 626 20000 6 chany_top_out[0]
port 63 nsew default tristate
rlabel metal2 s 4710 19520 4766 20000 6 chany_top_out[10]
port 64 nsew default tristate
rlabel metal2 s 5170 19520 5226 20000 6 chany_top_out[11]
port 65 nsew default tristate
rlabel metal2 s 5538 19520 5594 20000 6 chany_top_out[12]
port 66 nsew default tristate
rlabel metal2 s 5998 19520 6054 20000 6 chany_top_out[13]
port 67 nsew default tristate
rlabel metal2 s 6366 19520 6422 20000 6 chany_top_out[14]
port 68 nsew default tristate
rlabel metal2 s 6826 19520 6882 20000 6 chany_top_out[15]
port 69 nsew default tristate
rlabel metal2 s 7194 19520 7250 20000 6 chany_top_out[16]
port 70 nsew default tristate
rlabel metal2 s 7654 19520 7710 20000 6 chany_top_out[17]
port 71 nsew default tristate
rlabel metal2 s 8022 19520 8078 20000 6 chany_top_out[18]
port 72 nsew default tristate
rlabel metal2 s 8482 19520 8538 20000 6 chany_top_out[19]
port 73 nsew default tristate
rlabel metal2 s 1030 19520 1086 20000 6 chany_top_out[1]
port 74 nsew default tristate
rlabel metal2 s 1398 19520 1454 20000 6 chany_top_out[2]
port 75 nsew default tristate
rlabel metal2 s 1858 19520 1914 20000 6 chany_top_out[3]
port 76 nsew default tristate
rlabel metal2 s 2226 19520 2282 20000 6 chany_top_out[4]
port 77 nsew default tristate
rlabel metal2 s 2686 19520 2742 20000 6 chany_top_out[5]
port 78 nsew default tristate
rlabel metal2 s 3054 19520 3110 20000 6 chany_top_out[6]
port 79 nsew default tristate
rlabel metal2 s 3514 19520 3570 20000 6 chany_top_out[7]
port 80 nsew default tristate
rlabel metal2 s 3882 19520 3938 20000 6 chany_top_out[8]
port 81 nsew default tristate
rlabel metal2 s 4342 19520 4398 20000 6 chany_top_out[9]
port 82 nsew default tristate
rlabel metal3 s 0 8304 480 8424 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 83 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 84 nsew default input
rlabel metal3 s 0 14968 480 15088 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 85 nsew default tristate
rlabel metal3 s 0 4904 480 5024 6 left_grid_pin_0_
port 86 nsew default tristate
rlabel metal3 s 16520 7352 17000 7472 6 prog_clk_0_E_in
port 87 nsew default input
rlabel metal3 s 0 1640 480 1760 6 right_width_0_height_0__pin_0_
port 88 nsew default input
rlabel metal3 s 16520 2456 17000 2576 6 right_width_0_height_0__pin_1_lower
port 89 nsew default tristate
rlabel metal3 s 16520 17416 17000 17536 6 right_width_0_height_0__pin_1_upper
port 90 nsew default tristate
rlabel metal4 s 3409 2128 3729 17456 6 VPWR
port 91 nsew default input
rlabel metal4 s 5875 2128 6195 17456 6 VGND
port 92 nsew default input
<< properties >>
string FIXED_BBOX 0 0 17000 20000
<< end >>
