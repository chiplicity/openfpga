magic
tech sky130A
magscale 1 2
timestamp 1609018614
<< locali >>
rect 4445 18207 4479 18377
rect 12817 18139 12851 18377
rect 16129 15351 16163 15521
rect 4353 13719 4387 13889
rect 9045 11067 9079 11305
rect 13921 10455 13955 10557
rect 4537 8823 4571 8993
rect 9321 8415 9355 8585
<< viali >>
rect 1961 20553 1995 20587
rect 2513 20553 2547 20587
rect 9137 20553 9171 20587
rect 14289 20553 14323 20587
rect 8585 20417 8619 20451
rect 8769 20417 8803 20451
rect 1777 20349 1811 20383
rect 2329 20349 2363 20383
rect 12817 20349 12851 20383
rect 14105 20349 14139 20383
rect 7849 20281 7883 20315
rect 8493 20281 8527 20315
rect 13093 20281 13127 20315
rect 3157 20213 3191 20247
rect 4905 20213 4939 20247
rect 8125 20213 8159 20247
rect 4169 20009 4203 20043
rect 4905 20009 4939 20043
rect 9045 20009 9079 20043
rect 9689 20009 9723 20043
rect 11529 20009 11563 20043
rect 14197 20009 14231 20043
rect 14749 20009 14783 20043
rect 15485 20009 15519 20043
rect 16037 20009 16071 20043
rect 16589 20009 16623 20043
rect 17141 20009 17175 20043
rect 19165 20009 19199 20043
rect 1593 19873 1627 19907
rect 1869 19873 1903 19907
rect 2596 19873 2630 19907
rect 4997 19873 5031 19907
rect 5908 19873 5942 19907
rect 8953 19873 8987 19907
rect 10405 19873 10439 19907
rect 11989 19873 12023 19907
rect 12265 19873 12299 19907
rect 12725 19873 12759 19907
rect 13277 19873 13311 19907
rect 13553 19873 13587 19907
rect 14013 19873 14047 19907
rect 14565 19873 14599 19907
rect 15301 19873 15335 19907
rect 15853 19873 15887 19907
rect 16405 19873 16439 19907
rect 16957 19873 16991 19907
rect 17693 19873 17727 19907
rect 18429 19873 18463 19907
rect 18981 19873 19015 19907
rect 2329 19805 2363 19839
rect 5181 19805 5215 19839
rect 5641 19805 5675 19839
rect 9229 19805 9263 19839
rect 10149 19805 10183 19839
rect 17969 19805 18003 19839
rect 12909 19737 12943 19771
rect 18613 19737 18647 19771
rect 3709 19669 3743 19703
rect 4537 19669 4571 19703
rect 7021 19669 7055 19703
rect 8309 19669 8343 19703
rect 8585 19669 8619 19703
rect 1593 19465 1627 19499
rect 4445 19465 4479 19499
rect 6469 19465 6503 19499
rect 2145 19329 2179 19363
rect 9781 19329 9815 19363
rect 11805 19329 11839 19363
rect 15853 19329 15887 19363
rect 16589 19329 16623 19363
rect 1409 19261 1443 19295
rect 1961 19261 1995 19295
rect 3065 19261 3099 19295
rect 5089 19261 5123 19295
rect 7389 19261 7423 19295
rect 7656 19261 7690 19295
rect 11529 19261 11563 19295
rect 12572 19261 12606 19295
rect 13369 19261 13403 19295
rect 13645 19261 13679 19295
rect 14105 19261 14139 19295
rect 14749 19261 14783 19295
rect 15025 19261 15059 19295
rect 15577 19261 15611 19295
rect 16313 19261 16347 19295
rect 17049 19261 17083 19295
rect 18061 19261 18095 19295
rect 18337 19261 18371 19295
rect 18797 19261 18831 19295
rect 20545 19261 20579 19295
rect 3332 19193 3366 19227
rect 5356 19193 5390 19227
rect 10048 19193 10082 19227
rect 12817 19193 12851 19227
rect 17325 19193 17359 19227
rect 21189 19193 21223 19227
rect 4813 19125 4847 19159
rect 6837 19125 6871 19159
rect 8769 19125 8803 19159
rect 9321 19125 9355 19159
rect 11161 19125 11195 19159
rect 14289 19125 14323 19159
rect 18981 19125 19015 19159
rect 2881 18921 2915 18955
rect 3249 18921 3283 18955
rect 3341 18921 3375 18955
rect 4077 18921 4111 18955
rect 4445 18921 4479 18955
rect 6101 18921 6135 18955
rect 6469 18921 6503 18955
rect 7481 18921 7515 18955
rect 7941 18921 7975 18955
rect 8953 18921 8987 18955
rect 9045 18921 9079 18955
rect 11069 18921 11103 18955
rect 13185 18921 13219 18955
rect 14565 18921 14599 18955
rect 15669 18921 15703 18955
rect 16681 18921 16715 18955
rect 18429 18921 18463 18955
rect 18981 18921 19015 18955
rect 21373 18921 21407 18955
rect 2237 18853 2271 18887
rect 6561 18853 6595 18887
rect 7113 18853 7147 18887
rect 11612 18853 11646 18887
rect 1971 18785 2005 18819
rect 4537 18785 4571 18819
rect 5457 18785 5491 18819
rect 7849 18785 7883 18819
rect 9956 18785 9990 18819
rect 11345 18785 11379 18819
rect 13553 18785 13587 18819
rect 17509 18785 17543 18819
rect 18245 18785 18279 18819
rect 18797 18785 18831 18819
rect 3525 18717 3559 18751
rect 4629 18717 4663 18751
rect 5549 18717 5583 18751
rect 5733 18717 5767 18751
rect 6653 18717 6687 18751
rect 8033 18717 8067 18751
rect 9229 18717 9263 18751
rect 9689 18717 9723 18751
rect 13645 18717 13679 18751
rect 13737 18717 13771 18751
rect 14657 18717 14691 18751
rect 14749 18717 14783 18751
rect 15761 18717 15795 18751
rect 15945 18717 15979 18751
rect 16773 18717 16807 18751
rect 16865 18717 16899 18751
rect 17785 18717 17819 18751
rect 5089 18649 5123 18683
rect 14197 18649 14231 18683
rect 8585 18581 8619 18615
rect 12725 18581 12759 18615
rect 15301 18581 15335 18615
rect 16313 18581 16347 18615
rect 4353 18377 4387 18411
rect 4445 18377 4479 18411
rect 2973 18241 3007 18275
rect 12817 18377 12851 18411
rect 14289 18377 14323 18411
rect 14841 18377 14875 18411
rect 17233 18377 17267 18411
rect 6469 18309 6503 18343
rect 12541 18309 12575 18343
rect 7205 18241 7239 18275
rect 7849 18241 7883 18275
rect 8585 18241 8619 18275
rect 1777 18173 1811 18207
rect 2329 18173 2363 18207
rect 4445 18173 4479 18207
rect 4629 18173 4663 18207
rect 5089 18173 5123 18207
rect 7021 18173 7055 18207
rect 8309 18173 8343 18207
rect 15301 18241 15335 18275
rect 15393 18241 15427 18275
rect 18245 18241 18279 18275
rect 12909 18173 12943 18207
rect 13176 18173 13210 18207
rect 15209 18173 15243 18207
rect 15853 18173 15887 18207
rect 18061 18173 18095 18207
rect 3240 18105 3274 18139
rect 5356 18105 5390 18139
rect 12817 18105 12851 18139
rect 16120 18105 16154 18139
rect 1961 18037 1995 18071
rect 2513 18037 2547 18071
rect 17509 18037 17543 18071
rect 1777 17833 1811 17867
rect 3065 17833 3099 17867
rect 4537 17833 4571 17867
rect 5089 17833 5123 17867
rect 5641 17833 5675 17867
rect 6101 17833 6135 17867
rect 6653 17833 6687 17867
rect 8585 17833 8619 17867
rect 11345 17833 11379 17867
rect 13553 17833 13587 17867
rect 14565 17833 14599 17867
rect 16681 17833 16715 17867
rect 18153 17833 18187 17867
rect 9956 17765 9990 17799
rect 12357 17765 12391 17799
rect 14841 17765 14875 17799
rect 1593 17697 1627 17731
rect 2145 17697 2179 17731
rect 2421 17697 2455 17731
rect 2881 17697 2915 17731
rect 4445 17697 4479 17731
rect 6009 17697 6043 17731
rect 8309 17697 8343 17731
rect 8953 17697 8987 17731
rect 9689 17697 9723 17731
rect 11713 17697 11747 17731
rect 15557 17697 15591 17731
rect 18521 17697 18555 17731
rect 19165 17697 19199 17731
rect 4629 17629 4663 17663
rect 6193 17629 6227 17663
rect 7205 17629 7239 17663
rect 9045 17629 9079 17663
rect 9229 17629 9263 17663
rect 11805 17629 11839 17663
rect 11989 17629 12023 17663
rect 15301 17629 15335 17663
rect 18613 17629 18647 17663
rect 18797 17629 18831 17663
rect 8125 17561 8159 17595
rect 3617 17493 3651 17527
rect 4077 17493 4111 17527
rect 11069 17493 11103 17527
rect 12817 17493 12851 17527
rect 14105 17493 14139 17527
rect 16957 17493 16991 17527
rect 8769 17289 8803 17323
rect 9137 17289 9171 17323
rect 11345 17289 11379 17323
rect 13461 17289 13495 17323
rect 16957 17289 16991 17323
rect 2237 17153 2271 17187
rect 2973 17153 3007 17187
rect 3525 17153 3559 17187
rect 7113 17153 7147 17187
rect 9781 17153 9815 17187
rect 10149 17153 10183 17187
rect 11989 17153 12023 17187
rect 13001 17153 13035 17187
rect 14197 17153 14231 17187
rect 17601 17153 17635 17187
rect 1501 17085 1535 17119
rect 2053 17085 2087 17119
rect 2789 17085 2823 17119
rect 3792 17085 3826 17119
rect 7380 17085 7414 17119
rect 9597 17085 9631 17119
rect 10609 17085 10643 17119
rect 11069 17085 11103 17119
rect 13645 17085 13679 17119
rect 18153 17085 18187 17119
rect 11713 17017 11747 17051
rect 12909 17017 12943 17051
rect 14464 17017 14498 17051
rect 18420 17017 18454 17051
rect 1685 16949 1719 16983
rect 4905 16949 4939 16983
rect 5549 16949 5583 16983
rect 8493 16949 8527 16983
rect 9505 16949 9539 16983
rect 11805 16949 11839 16983
rect 12449 16949 12483 16983
rect 12817 16949 12851 16983
rect 15577 16949 15611 16983
rect 17325 16949 17359 16983
rect 17417 16949 17451 16983
rect 19533 16949 19567 16983
rect 1961 16745 1995 16779
rect 2973 16745 3007 16779
rect 3433 16745 3467 16779
rect 6285 16745 6319 16779
rect 8953 16745 8987 16779
rect 10241 16745 10275 16779
rect 12357 16745 12391 16779
rect 12909 16745 12943 16779
rect 14381 16745 14415 16779
rect 15301 16745 15335 16779
rect 17785 16745 17819 16779
rect 19441 16745 19475 16779
rect 11244 16677 11278 16711
rect 13277 16677 13311 16711
rect 16672 16677 16706 16711
rect 18306 16677 18340 16711
rect 1777 16609 1811 16643
rect 3341 16609 3375 16643
rect 4077 16609 4111 16643
rect 5172 16609 5206 16643
rect 6929 16609 6963 16643
rect 7196 16609 7230 16643
rect 9689 16609 9723 16643
rect 10609 16609 10643 16643
rect 10977 16609 11011 16643
rect 13369 16609 13403 16643
rect 14289 16609 14323 16643
rect 16405 16609 16439 16643
rect 18061 16609 18095 16643
rect 3617 16541 3651 16575
rect 4905 16541 4939 16575
rect 9045 16541 9079 16575
rect 9137 16541 9171 16575
rect 13553 16541 13587 16575
rect 14565 16541 14599 16575
rect 8585 16473 8619 16507
rect 8309 16405 8343 16439
rect 13921 16405 13955 16439
rect 15669 16405 15703 16439
rect 1685 16201 1719 16235
rect 7389 16201 7423 16235
rect 10057 16201 10091 16235
rect 10333 16201 10367 16235
rect 12449 16201 12483 16235
rect 15025 16201 15059 16235
rect 18061 16201 18095 16235
rect 4905 16133 4939 16167
rect 16589 16133 16623 16167
rect 2237 16065 2271 16099
rect 5457 16065 5491 16099
rect 8033 16065 8067 16099
rect 8677 16065 8711 16099
rect 10977 16065 11011 16099
rect 11989 16065 12023 16099
rect 13001 16065 13035 16099
rect 15761 16065 15795 16099
rect 15945 16065 15979 16099
rect 17049 16065 17083 16099
rect 18613 16065 18647 16099
rect 1501 15997 1535 16031
rect 2053 15997 2087 16031
rect 6377 15997 6411 16031
rect 7021 15997 7055 16031
rect 12817 15997 12851 16031
rect 13645 15997 13679 16031
rect 16773 15997 16807 16031
rect 5273 15929 5307 15963
rect 5917 15929 5951 15963
rect 7757 15929 7791 15963
rect 7849 15929 7883 15963
rect 8944 15929 8978 15963
rect 11713 15929 11747 15963
rect 13912 15929 13946 15963
rect 15669 15929 15703 15963
rect 5365 15861 5399 15895
rect 6837 15861 6871 15895
rect 10701 15861 10735 15895
rect 10793 15861 10827 15895
rect 11345 15861 11379 15895
rect 11805 15861 11839 15895
rect 12909 15861 12943 15895
rect 15301 15861 15335 15895
rect 17601 15861 17635 15895
rect 18429 15861 18463 15895
rect 18521 15861 18555 15895
rect 1685 15657 1719 15691
rect 2973 15657 3007 15691
rect 6377 15657 6411 15691
rect 6837 15657 6871 15691
rect 7389 15657 7423 15691
rect 8585 15657 8619 15691
rect 9045 15657 9079 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 12541 15657 12575 15691
rect 14013 15657 14047 15691
rect 14381 15657 14415 15691
rect 16221 15657 16255 15691
rect 11152 15589 11186 15623
rect 14473 15589 14507 15623
rect 17233 15589 17267 15623
rect 18788 15589 18822 15623
rect 1501 15521 1535 15555
rect 2053 15521 2087 15555
rect 2789 15521 2823 15555
rect 4721 15521 4755 15555
rect 4988 15521 5022 15555
rect 6745 15521 6779 15555
rect 7573 15521 7607 15555
rect 8125 15521 8159 15555
rect 8953 15521 8987 15555
rect 10057 15521 10091 15555
rect 10885 15521 10919 15555
rect 13277 15521 13311 15555
rect 15669 15521 15703 15555
rect 16129 15521 16163 15555
rect 16589 15521 16623 15555
rect 17601 15521 17635 15555
rect 18521 15521 18555 15555
rect 2237 15453 2271 15487
rect 6929 15453 6963 15487
rect 9229 15453 9263 15487
rect 10241 15453 10275 15487
rect 13553 15453 13587 15487
rect 14657 15453 14691 15487
rect 13093 15385 13127 15419
rect 15485 15385 15519 15419
rect 16681 15453 16715 15487
rect 16773 15453 16807 15487
rect 17969 15385 18003 15419
rect 3341 15317 3375 15351
rect 6101 15317 6135 15351
rect 12265 15317 12299 15351
rect 16129 15317 16163 15351
rect 19901 15317 19935 15351
rect 1685 15113 1719 15147
rect 4537 15113 4571 15147
rect 6285 15113 6319 15147
rect 7205 15113 7239 15147
rect 9413 15113 9447 15147
rect 11345 15113 11379 15147
rect 12541 15113 12575 15147
rect 14013 15113 14047 15147
rect 15485 15113 15519 15147
rect 17325 15113 17359 15147
rect 12081 15045 12115 15079
rect 15025 15045 15059 15079
rect 19073 15045 19107 15079
rect 2237 14977 2271 15011
rect 2881 14977 2915 15011
rect 13369 14977 13403 15011
rect 13553 14977 13587 15011
rect 14473 14977 14507 15011
rect 14657 14977 14691 15011
rect 18521 14977 18555 15011
rect 18705 14977 18739 15011
rect 1501 14909 1535 14943
rect 2053 14909 2087 14943
rect 3148 14909 3182 14943
rect 8033 14909 8067 14943
rect 9689 14909 9723 14943
rect 13277 14909 13311 14943
rect 14381 14909 14415 14943
rect 15945 14909 15979 14943
rect 19993 14909 20027 14943
rect 20260 14909 20294 14943
rect 8300 14841 8334 14875
rect 9956 14841 9990 14875
rect 16212 14841 16246 14875
rect 18429 14841 18463 14875
rect 4261 14773 4295 14807
rect 11069 14773 11103 14807
rect 12909 14773 12943 14807
rect 17601 14773 17635 14807
rect 18061 14773 18095 14807
rect 21373 14773 21407 14807
rect 2421 14569 2455 14603
rect 2973 14569 3007 14603
rect 3341 14569 3375 14603
rect 3433 14569 3467 14603
rect 5457 14569 5491 14603
rect 5733 14569 5767 14603
rect 8953 14569 8987 14603
rect 9689 14569 9723 14603
rect 10517 14569 10551 14603
rect 14289 14569 14323 14603
rect 16681 14569 16715 14603
rect 6101 14501 6135 14535
rect 8493 14501 8527 14535
rect 10885 14501 10919 14535
rect 13154 14501 13188 14535
rect 17960 14501 17994 14535
rect 2329 14433 2363 14467
rect 4333 14433 4367 14467
rect 6193 14433 6227 14467
rect 7104 14433 7138 14467
rect 9137 14433 9171 14467
rect 12909 14433 12943 14467
rect 15301 14433 15335 14467
rect 15568 14433 15602 14467
rect 17693 14433 17727 14467
rect 1685 14365 1719 14399
rect 2513 14365 2547 14399
rect 3617 14365 3651 14399
rect 4077 14365 4111 14399
rect 6377 14365 6411 14399
rect 6837 14365 6871 14399
rect 16957 14365 16991 14399
rect 19349 14365 19383 14399
rect 12173 14297 12207 14331
rect 1961 14229 1995 14263
rect 8217 14229 8251 14263
rect 14565 14229 14599 14263
rect 19073 14229 19107 14263
rect 21373 14229 21407 14263
rect 1685 14025 1719 14059
rect 5917 14025 5951 14059
rect 8217 14025 8251 14059
rect 11345 14025 11379 14059
rect 14197 14025 14231 14059
rect 16221 14025 16255 14059
rect 18061 14025 18095 14059
rect 6377 13957 6411 13991
rect 10149 13957 10183 13991
rect 13829 13957 13863 13991
rect 17325 13957 17359 13991
rect 2237 13889 2271 13923
rect 2973 13889 3007 13923
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 11897 13889 11931 13923
rect 14841 13889 14875 13923
rect 15669 13889 15703 13923
rect 15853 13889 15887 13923
rect 16773 13889 16807 13923
rect 18521 13889 18555 13923
rect 18705 13889 18739 13923
rect 1501 13821 1535 13855
rect 2053 13821 2087 13855
rect 2789 13821 2823 13855
rect 3985 13821 4019 13855
rect 4537 13821 4571 13855
rect 6837 13821 6871 13855
rect 7104 13821 7138 13855
rect 8769 13821 8803 13855
rect 11805 13821 11839 13855
rect 12449 13821 12483 13855
rect 12716 13821 12750 13855
rect 14657 13821 14691 13855
rect 16589 13821 16623 13855
rect 4804 13753 4838 13787
rect 9036 13753 9070 13787
rect 16681 13753 16715 13787
rect 18429 13753 18463 13787
rect 3525 13685 3559 13719
rect 3893 13685 3927 13719
rect 4353 13685 4387 13719
rect 11713 13685 11747 13719
rect 14565 13685 14599 13719
rect 15209 13685 15243 13719
rect 15577 13685 15611 13719
rect 2973 13481 3007 13515
rect 3525 13481 3559 13515
rect 5457 13481 5491 13515
rect 5733 13481 5767 13515
rect 7021 13481 7055 13515
rect 8585 13481 8619 13515
rect 9045 13481 9079 13515
rect 9689 13481 9723 13515
rect 10149 13481 10183 13515
rect 10793 13481 10827 13515
rect 12909 13481 12943 13515
rect 13553 13481 13587 13515
rect 15761 13481 15795 13515
rect 2329 13413 2363 13447
rect 4344 13413 4378 13447
rect 7481 13413 7515 13447
rect 11253 13413 11287 13447
rect 18052 13413 18086 13447
rect 2053 13345 2087 13379
rect 6101 13345 6135 13379
rect 7389 13345 7423 13379
rect 8953 13345 8987 13379
rect 10057 13345 10091 13379
rect 11796 13345 11830 13379
rect 15669 13345 15703 13379
rect 4077 13277 4111 13311
rect 6193 13277 6227 13311
rect 6285 13277 6319 13311
rect 7665 13277 7699 13311
rect 9229 13277 9263 13311
rect 10241 13277 10275 13311
rect 11529 13277 11563 13311
rect 13645 13277 13679 13311
rect 13737 13277 13771 13311
rect 15853 13277 15887 13311
rect 16313 13277 16347 13311
rect 17785 13277 17819 13311
rect 8033 13209 8067 13243
rect 14473 13209 14507 13243
rect 17417 13209 17451 13243
rect 13185 13141 13219 13175
rect 14841 13141 14875 13175
rect 15301 13141 15335 13175
rect 19165 13141 19199 13175
rect 1961 12937 1995 12971
rect 2513 12937 2547 12971
rect 3617 12937 3651 12971
rect 5825 12937 5859 12971
rect 8493 12937 8527 12971
rect 11345 12937 11379 12971
rect 12541 12937 12575 12971
rect 13553 12937 13587 12971
rect 14657 12937 14691 12971
rect 16405 12937 16439 12971
rect 16681 12937 16715 12971
rect 19073 12937 19107 12971
rect 9045 12801 9079 12835
rect 9505 12801 9539 12835
rect 11989 12801 12023 12835
rect 13001 12801 13035 12835
rect 13185 12801 13219 12835
rect 17141 12801 17175 12835
rect 17233 12801 17267 12835
rect 18521 12801 18555 12835
rect 18705 12801 18739 12835
rect 19625 12801 19659 12835
rect 1777 12733 1811 12767
rect 2329 12733 2363 12767
rect 2881 12733 2915 12767
rect 3433 12733 3467 12767
rect 4445 12733 4479 12767
rect 6837 12733 6871 12767
rect 7104 12733 7138 12767
rect 9965 12733 9999 12767
rect 10701 12733 10735 12767
rect 12909 12733 12943 12767
rect 14381 12733 14415 12767
rect 15025 12733 15059 12767
rect 17049 12733 17083 12767
rect 4712 12665 4746 12699
rect 8861 12665 8895 12699
rect 11713 12665 11747 12699
rect 15292 12665 15326 12699
rect 19533 12665 19567 12699
rect 3065 12597 3099 12631
rect 6469 12597 6503 12631
rect 8217 12597 8251 12631
rect 8953 12597 8987 12631
rect 11069 12597 11103 12631
rect 11805 12597 11839 12631
rect 14197 12597 14231 12631
rect 18061 12597 18095 12631
rect 18429 12597 18463 12631
rect 19441 12597 19475 12631
rect 9321 12393 9355 12427
rect 11621 12393 11655 12427
rect 14105 12393 14139 12427
rect 16681 12393 16715 12427
rect 19349 12393 19383 12427
rect 3157 12325 3191 12359
rect 8208 12325 8242 12359
rect 9689 12325 9723 12359
rect 10517 12325 10551 12359
rect 12440 12325 12474 12359
rect 15568 12325 15602 12359
rect 2145 12257 2179 12291
rect 2881 12257 2915 12291
rect 4344 12257 4378 12291
rect 6285 12257 6319 12291
rect 6929 12257 6963 12291
rect 7021 12257 7055 12291
rect 7573 12257 7607 12291
rect 7941 12257 7975 12291
rect 10425 12257 10459 12291
rect 11529 12257 11563 12291
rect 12173 12257 12207 12291
rect 14473 12257 14507 12291
rect 15301 12257 15335 12291
rect 17233 12257 17267 12291
rect 17500 12257 17534 12291
rect 2421 12189 2455 12223
rect 4077 12189 4111 12223
rect 7113 12189 7147 12223
rect 10609 12189 10643 12223
rect 11713 12189 11747 12223
rect 14565 12189 14599 12223
rect 14749 12189 14783 12223
rect 18889 12189 18923 12223
rect 5457 12053 5491 12087
rect 5733 12053 5767 12087
rect 6101 12053 6135 12087
rect 6561 12053 6595 12087
rect 10057 12053 10091 12087
rect 11161 12053 11195 12087
rect 13553 12053 13587 12087
rect 18613 12053 18647 12087
rect 8493 11849 8527 11883
rect 11345 11849 11379 11883
rect 13829 11849 13863 11883
rect 15577 11849 15611 11883
rect 18061 11849 18095 11883
rect 3893 11781 3927 11815
rect 16129 11781 16163 11815
rect 2053 11713 2087 11747
rect 2789 11713 2823 11747
rect 4353 11713 4387 11747
rect 4537 11713 4571 11747
rect 5457 11713 5491 11747
rect 9689 11713 9723 11747
rect 11805 11713 11839 11747
rect 11897 11713 11931 11747
rect 12541 11713 12575 11747
rect 14197 11713 14231 11747
rect 18613 11713 18647 11747
rect 1777 11645 1811 11679
rect 2513 11645 2547 11679
rect 7113 11645 7147 11679
rect 9956 11645 9990 11679
rect 11713 11645 11747 11679
rect 13185 11645 13219 11679
rect 16313 11645 16347 11679
rect 18429 11645 18463 11679
rect 4261 11577 4295 11611
rect 5273 11577 5307 11611
rect 5917 11577 5951 11611
rect 7358 11577 7392 11611
rect 8861 11577 8895 11611
rect 14464 11577 14498 11611
rect 4905 11509 4939 11543
rect 5365 11509 5399 11543
rect 6377 11509 6411 11543
rect 9137 11509 9171 11543
rect 11069 11509 11103 11543
rect 13001 11509 13035 11543
rect 13461 11509 13495 11543
rect 17601 11509 17635 11543
rect 18521 11509 18555 11543
rect 1961 11305 1995 11339
rect 2421 11305 2455 11339
rect 2973 11305 3007 11339
rect 3433 11305 3467 11339
rect 4077 11305 4111 11339
rect 4537 11305 4571 11339
rect 6653 11305 6687 11339
rect 7665 11305 7699 11339
rect 9045 11305 9079 11339
rect 9137 11305 9171 11339
rect 10333 11305 10367 11339
rect 12633 11305 12667 11339
rect 13645 11305 13679 11339
rect 14105 11305 14139 11339
rect 14657 11305 14691 11339
rect 18889 11305 18923 11339
rect 7021 11237 7055 11271
rect 8125 11237 8159 11271
rect 8677 11237 8711 11271
rect 2329 11169 2363 11203
rect 3341 11169 3375 11203
rect 4445 11169 4479 11203
rect 5457 11169 5491 11203
rect 6377 11169 6411 11203
rect 8033 11169 8067 11203
rect 2605 11101 2639 11135
rect 3525 11101 3559 11135
rect 4721 11101 4755 11135
rect 5181 11101 5215 11135
rect 5825 11101 5859 11135
rect 7113 11101 7147 11135
rect 7297 11101 7331 11135
rect 8217 11101 8251 11135
rect 15936 11237 15970 11271
rect 17776 11237 17810 11271
rect 9321 11169 9355 11203
rect 10977 11169 11011 11203
rect 11244 11169 11278 11203
rect 13001 11169 13035 11203
rect 14013 11169 14047 11203
rect 15669 11169 15703 11203
rect 17509 11169 17543 11203
rect 13093 11101 13127 11135
rect 13185 11101 13219 11135
rect 14289 11101 14323 11135
rect 6193 11033 6227 11067
rect 9045 11033 9079 11067
rect 12357 11033 12391 11067
rect 17049 10965 17083 10999
rect 1777 10761 1811 10795
rect 4169 10761 4203 10795
rect 4537 10761 4571 10795
rect 5733 10761 5767 10795
rect 8217 10761 8251 10795
rect 11529 10761 11563 10795
rect 13829 10761 13863 10795
rect 15485 10761 15519 10795
rect 17693 10693 17727 10727
rect 2421 10625 2455 10659
rect 4905 10625 4939 10659
rect 6377 10625 6411 10659
rect 10149 10625 10183 10659
rect 16313 10625 16347 10659
rect 2789 10557 2823 10591
rect 5273 10557 5307 10591
rect 6837 10557 6871 10591
rect 7093 10557 7127 10591
rect 8493 10557 8527 10591
rect 12449 10557 12483 10591
rect 12716 10557 12750 10591
rect 13921 10557 13955 10591
rect 14105 10557 14139 10591
rect 14372 10557 14406 10591
rect 16580 10557 16614 10591
rect 3056 10489 3090 10523
rect 8760 10489 8794 10523
rect 10416 10489 10450 10523
rect 11897 10489 11931 10523
rect 2145 10421 2179 10455
rect 2237 10421 2271 10455
rect 6101 10421 6135 10455
rect 6193 10421 6227 10455
rect 9873 10421 9907 10455
rect 13921 10421 13955 10455
rect 18061 10421 18095 10455
rect 3433 10217 3467 10251
rect 4077 10217 4111 10251
rect 4537 10217 4571 10251
rect 6745 10217 6779 10251
rect 7389 10217 7423 10251
rect 7757 10217 7791 10251
rect 8401 10217 8435 10251
rect 9689 10217 9723 10251
rect 10057 10217 10091 10251
rect 10885 10217 10919 10251
rect 12265 10217 12299 10251
rect 15485 10217 15519 10251
rect 16589 10217 16623 10251
rect 16957 10217 16991 10251
rect 2044 10149 2078 10183
rect 7021 10149 7055 10183
rect 8769 10149 8803 10183
rect 17049 10149 17083 10183
rect 1777 10081 1811 10115
rect 4445 10081 4479 10115
rect 5365 10081 5399 10115
rect 5632 10081 5666 10115
rect 11253 10081 11287 10115
rect 11345 10081 11379 10115
rect 14933 10081 14967 10115
rect 15853 10081 15887 10115
rect 4721 10013 4755 10047
rect 7849 10013 7883 10047
rect 8033 10013 8067 10047
rect 8861 10013 8895 10047
rect 8953 10013 8987 10047
rect 10149 10013 10183 10047
rect 10241 10013 10275 10047
rect 11437 10013 11471 10047
rect 11989 10013 12023 10047
rect 15945 10013 15979 10047
rect 16129 10013 16163 10047
rect 17141 10013 17175 10047
rect 3157 9877 3191 9911
rect 2881 9673 2915 9707
rect 6837 9673 6871 9707
rect 9413 9673 9447 9707
rect 9781 9673 9815 9707
rect 15117 9673 15151 9707
rect 1961 9605 1995 9639
rect 11161 9605 11195 9639
rect 2605 9537 2639 9571
rect 3341 9537 3375 9571
rect 3525 9537 3559 9571
rect 4813 9537 4847 9571
rect 7481 9537 7515 9571
rect 10701 9537 10735 9571
rect 1777 9469 1811 9503
rect 8033 9469 8067 9503
rect 3893 9401 3927 9435
rect 6285 9401 6319 9435
rect 7205 9401 7239 9435
rect 8300 9401 8334 9435
rect 3249 9333 3283 9367
rect 4261 9333 4295 9367
rect 4629 9333 4663 9367
rect 4721 9333 4755 9367
rect 7297 9333 7331 9367
rect 1961 9129 1995 9163
rect 4629 9129 4663 9163
rect 7941 9129 7975 9163
rect 8585 9129 8619 9163
rect 1777 8993 1811 9027
rect 2329 8993 2363 9027
rect 2596 8993 2630 9027
rect 4537 8993 4571 9027
rect 4997 8993 5031 9027
rect 5641 8993 5675 9027
rect 7205 8993 7239 9027
rect 8033 8993 8067 9027
rect 5089 8925 5123 8959
rect 5181 8925 5215 8959
rect 8125 8925 8159 8959
rect 3709 8789 3743 8823
rect 4261 8789 4295 8823
rect 4537 8789 4571 8823
rect 6653 8789 6687 8823
rect 7573 8789 7607 8823
rect 4905 8585 4939 8619
rect 6009 8585 6043 8619
rect 8493 8585 8527 8619
rect 9321 8585 9355 8619
rect 9597 8585 9631 8619
rect 4537 8517 4571 8551
rect 2237 8449 2271 8483
rect 5365 8449 5399 8483
rect 5457 8449 5491 8483
rect 9045 8449 9079 8483
rect 2053 8381 2087 8415
rect 3157 8381 3191 8415
rect 3424 8381 3458 8415
rect 6837 8381 6871 8415
rect 8861 8381 8895 8415
rect 8953 8381 8987 8415
rect 9321 8381 9355 8415
rect 5273 8313 5307 8347
rect 6285 8313 6319 8347
rect 7104 8313 7138 8347
rect 8217 8245 8251 8279
rect 2973 8041 3007 8075
rect 3433 8041 3467 8075
rect 7113 8041 7147 8075
rect 10149 8041 10183 8075
rect 2237 7973 2271 8007
rect 4344 7973 4378 8007
rect 1950 7905 1984 7939
rect 3341 7905 3375 7939
rect 5989 7905 6023 7939
rect 7389 7905 7423 7939
rect 7656 7905 7690 7939
rect 10057 7905 10091 7939
rect 3617 7837 3651 7871
rect 4077 7837 4111 7871
rect 5733 7837 5767 7871
rect 10241 7837 10275 7871
rect 8769 7769 8803 7803
rect 5457 7701 5491 7735
rect 9689 7701 9723 7735
rect 4169 7497 4203 7531
rect 8125 7497 8159 7531
rect 19441 7497 19475 7531
rect 7113 7429 7147 7463
rect 18889 7429 18923 7463
rect 4721 7361 4755 7395
rect 7757 7361 7791 7395
rect 8769 7361 8803 7395
rect 18337 7293 18371 7327
rect 18705 7293 18739 7327
rect 19257 7293 19291 7327
rect 19809 7293 19843 7327
rect 4537 7225 4571 7259
rect 5181 7225 5215 7259
rect 7481 7225 7515 7259
rect 8585 7225 8619 7259
rect 9137 7225 9171 7259
rect 3801 7157 3835 7191
rect 4629 7157 4663 7191
rect 6377 7157 6411 7191
rect 7573 7157 7607 7191
rect 8493 7157 8527 7191
rect 9505 7157 9539 7191
rect 7665 6953 7699 6987
rect 7573 6817 7607 6851
rect 8217 6817 8251 6851
rect 19625 6817 19659 6851
rect 20177 6817 20211 6851
rect 6745 6749 6779 6783
rect 7757 6749 7791 6783
rect 19809 6681 19843 6715
rect 7205 6613 7239 6647
rect 20177 6409 20211 6443
rect 19993 6205 20027 6239
rect 20545 6137 20579 6171
rect 21097 5865 21131 5899
rect 20913 5729 20947 5763
rect 20453 5525 20487 5559
rect 21005 5321 21039 5355
rect 20821 5117 20855 5151
rect 20453 4981 20487 5015
<< metal1 >>
rect 2958 21904 2964 21956
rect 3016 21944 3022 21956
rect 3970 21944 3976 21956
rect 3016 21916 3976 21944
rect 3016 21904 3022 21916
rect 3970 21904 3976 21916
rect 4028 21904 4034 21956
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 1946 20584 1952 20596
rect 1907 20556 1952 20584
rect 1946 20544 1952 20556
rect 2004 20544 2010 20596
rect 2501 20587 2559 20593
rect 2501 20553 2513 20587
rect 2547 20584 2559 20587
rect 2774 20584 2780 20596
rect 2547 20556 2780 20584
rect 2547 20553 2559 20556
rect 2501 20547 2559 20553
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 8938 20584 8944 20596
rect 8588 20556 8944 20584
rect 8588 20457 8616 20556
rect 8938 20544 8944 20556
rect 8996 20584 9002 20596
rect 9125 20587 9183 20593
rect 9125 20584 9137 20587
rect 8996 20556 9137 20584
rect 8996 20544 9002 20556
rect 9125 20553 9137 20556
rect 9171 20553 9183 20587
rect 9125 20547 9183 20553
rect 14277 20587 14335 20593
rect 14277 20553 14289 20587
rect 14323 20584 14335 20587
rect 14918 20584 14924 20596
rect 14323 20556 14924 20584
rect 14323 20553 14335 20556
rect 14277 20547 14335 20553
rect 14918 20544 14924 20556
rect 14976 20544 14982 20596
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20417 8631 20451
rect 8754 20448 8760 20460
rect 8715 20420 8760 20448
rect 8573 20411 8631 20417
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 1762 20380 1768 20392
rect 1723 20352 1768 20380
rect 1762 20340 1768 20352
rect 1820 20340 1826 20392
rect 1854 20340 1860 20392
rect 1912 20380 1918 20392
rect 2317 20383 2375 20389
rect 2317 20380 2329 20383
rect 1912 20352 2329 20380
rect 1912 20340 1918 20352
rect 2317 20349 2329 20352
rect 2363 20349 2375 20383
rect 12802 20380 12808 20392
rect 12763 20352 12808 20380
rect 2317 20343 2375 20349
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 14090 20380 14096 20392
rect 14051 20352 14096 20380
rect 14090 20340 14096 20352
rect 14148 20340 14154 20392
rect 4154 20272 4160 20324
rect 4212 20312 4218 20324
rect 7837 20315 7895 20321
rect 7837 20312 7849 20315
rect 4212 20284 7849 20312
rect 4212 20272 4218 20284
rect 7837 20281 7849 20284
rect 7883 20312 7895 20315
rect 8481 20315 8539 20321
rect 8481 20312 8493 20315
rect 7883 20284 8493 20312
rect 7883 20281 7895 20284
rect 7837 20275 7895 20281
rect 8481 20281 8493 20284
rect 8527 20281 8539 20315
rect 8481 20275 8539 20281
rect 13081 20315 13139 20321
rect 13081 20281 13093 20315
rect 13127 20312 13139 20315
rect 14550 20312 14556 20324
rect 13127 20284 14556 20312
rect 13127 20281 13139 20284
rect 13081 20275 13139 20281
rect 14550 20272 14556 20284
rect 14608 20272 14614 20324
rect 3142 20244 3148 20256
rect 3103 20216 3148 20244
rect 3142 20204 3148 20216
rect 3200 20204 3206 20256
rect 4890 20244 4896 20256
rect 4851 20216 4896 20244
rect 4890 20204 4896 20216
rect 4948 20204 4954 20256
rect 8113 20247 8171 20253
rect 8113 20213 8125 20247
rect 8159 20244 8171 20247
rect 8202 20244 8208 20256
rect 8159 20216 8208 20244
rect 8159 20213 8171 20216
rect 8113 20207 8171 20213
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 11054 20204 11060 20256
rect 11112 20244 11118 20256
rect 12158 20244 12164 20256
rect 11112 20216 12164 20244
rect 11112 20204 11118 20216
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 4154 20040 4160 20052
rect 4115 20012 4160 20040
rect 4154 20000 4160 20012
rect 4212 20000 4218 20052
rect 4890 20040 4896 20052
rect 4851 20012 4896 20040
rect 4890 20000 4896 20012
rect 4948 20000 4954 20052
rect 9033 20043 9091 20049
rect 9033 20009 9045 20043
rect 9079 20040 9091 20043
rect 9398 20040 9404 20052
rect 9079 20012 9404 20040
rect 9079 20009 9091 20012
rect 9033 20003 9091 20009
rect 9398 20000 9404 20012
rect 9456 20040 9462 20052
rect 9677 20043 9735 20049
rect 9677 20040 9689 20043
rect 9456 20012 9689 20040
rect 9456 20000 9462 20012
rect 9677 20009 9689 20012
rect 9723 20009 9735 20043
rect 9677 20003 9735 20009
rect 11517 20043 11575 20049
rect 11517 20009 11529 20043
rect 11563 20009 11575 20043
rect 11517 20003 11575 20009
rect 2866 19972 2872 19984
rect 1596 19944 2872 19972
rect 1596 19913 1624 19944
rect 2866 19932 2872 19944
rect 2924 19932 2930 19984
rect 8754 19932 8760 19984
rect 8812 19972 8818 19984
rect 11532 19972 11560 20003
rect 13538 20000 13544 20052
rect 13596 20040 13602 20052
rect 14185 20043 14243 20049
rect 14185 20040 14197 20043
rect 13596 20012 14197 20040
rect 13596 20000 13602 20012
rect 14185 20009 14197 20012
rect 14231 20009 14243 20043
rect 14185 20003 14243 20009
rect 14458 20000 14464 20052
rect 14516 20040 14522 20052
rect 14737 20043 14795 20049
rect 14737 20040 14749 20043
rect 14516 20012 14749 20040
rect 14516 20000 14522 20012
rect 14737 20009 14749 20012
rect 14783 20009 14795 20043
rect 14737 20003 14795 20009
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 15473 20043 15531 20049
rect 15473 20040 15485 20043
rect 15436 20012 15485 20040
rect 15436 20000 15442 20012
rect 15473 20009 15485 20012
rect 15519 20009 15531 20043
rect 15473 20003 15531 20009
rect 15838 20000 15844 20052
rect 15896 20040 15902 20052
rect 16025 20043 16083 20049
rect 16025 20040 16037 20043
rect 15896 20012 16037 20040
rect 15896 20000 15902 20012
rect 16025 20009 16037 20012
rect 16071 20009 16083 20043
rect 16025 20003 16083 20009
rect 16298 20000 16304 20052
rect 16356 20040 16362 20052
rect 16577 20043 16635 20049
rect 16577 20040 16589 20043
rect 16356 20012 16589 20040
rect 16356 20000 16362 20012
rect 16577 20009 16589 20012
rect 16623 20009 16635 20043
rect 16577 20003 16635 20009
rect 16758 20000 16764 20052
rect 16816 20040 16822 20052
rect 17129 20043 17187 20049
rect 17129 20040 17141 20043
rect 16816 20012 17141 20040
rect 16816 20000 16822 20012
rect 17129 20009 17141 20012
rect 17175 20009 17187 20043
rect 17129 20003 17187 20009
rect 18598 20000 18604 20052
rect 18656 20040 18662 20052
rect 19153 20043 19211 20049
rect 19153 20040 19165 20043
rect 18656 20012 19165 20040
rect 18656 20000 18662 20012
rect 19153 20009 19165 20012
rect 19199 20009 19211 20043
rect 19153 20003 19211 20009
rect 18874 19972 18880 19984
rect 8812 19944 11560 19972
rect 17696 19944 18880 19972
rect 8812 19932 8818 19944
rect 1581 19907 1639 19913
rect 1581 19873 1593 19907
rect 1627 19873 1639 19907
rect 1854 19904 1860 19916
rect 1815 19876 1860 19904
rect 1581 19867 1639 19873
rect 1854 19864 1860 19876
rect 1912 19864 1918 19916
rect 2584 19907 2642 19913
rect 2584 19873 2596 19907
rect 2630 19904 2642 19907
rect 4338 19904 4344 19916
rect 2630 19876 4344 19904
rect 2630 19873 2642 19876
rect 2584 19867 2642 19873
rect 4338 19864 4344 19876
rect 4396 19864 4402 19916
rect 4985 19907 5043 19913
rect 4985 19873 4997 19907
rect 5031 19904 5043 19907
rect 5718 19904 5724 19916
rect 5031 19876 5724 19904
rect 5031 19873 5043 19876
rect 4985 19867 5043 19873
rect 5718 19864 5724 19876
rect 5776 19864 5782 19916
rect 5896 19907 5954 19913
rect 5896 19873 5908 19907
rect 5942 19904 5954 19907
rect 6454 19904 6460 19916
rect 5942 19876 6460 19904
rect 5942 19873 5954 19876
rect 5896 19867 5954 19873
rect 6454 19864 6460 19876
rect 6512 19864 6518 19916
rect 8294 19864 8300 19916
rect 8352 19904 8358 19916
rect 8941 19907 8999 19913
rect 8941 19904 8953 19907
rect 8352 19876 8953 19904
rect 8352 19864 8358 19876
rect 8941 19873 8953 19876
rect 8987 19873 8999 19907
rect 8941 19867 8999 19873
rect 9766 19864 9772 19916
rect 9824 19904 9830 19916
rect 10393 19907 10451 19913
rect 10393 19904 10405 19907
rect 9824 19876 10405 19904
rect 9824 19864 9830 19876
rect 10393 19873 10405 19876
rect 10439 19873 10451 19907
rect 11974 19904 11980 19916
rect 11935 19876 11980 19904
rect 10393 19867 10451 19873
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 12253 19907 12311 19913
rect 12253 19873 12265 19907
rect 12299 19904 12311 19907
rect 12713 19907 12771 19913
rect 12713 19904 12725 19907
rect 12299 19876 12725 19904
rect 12299 19873 12311 19876
rect 12253 19867 12311 19873
rect 12713 19873 12725 19876
rect 12759 19873 12771 19907
rect 12713 19867 12771 19873
rect 13265 19907 13323 19913
rect 13265 19873 13277 19907
rect 13311 19873 13323 19907
rect 13265 19867 13323 19873
rect 13541 19907 13599 19913
rect 13541 19873 13553 19907
rect 13587 19904 13599 19907
rect 14001 19907 14059 19913
rect 14001 19904 14013 19907
rect 13587 19876 14013 19904
rect 13587 19873 13599 19876
rect 13541 19867 13599 19873
rect 14001 19873 14013 19876
rect 14047 19873 14059 19907
rect 14550 19904 14556 19916
rect 14511 19876 14556 19904
rect 14001 19867 14059 19873
rect 2317 19839 2375 19845
rect 2317 19805 2329 19839
rect 2363 19805 2375 19839
rect 2317 19799 2375 19805
rect 5169 19839 5227 19845
rect 5169 19805 5181 19839
rect 5215 19805 5227 19839
rect 5169 19799 5227 19805
rect 2332 19700 2360 19799
rect 2682 19700 2688 19712
rect 2332 19672 2688 19700
rect 2682 19660 2688 19672
rect 2740 19660 2746 19712
rect 3694 19700 3700 19712
rect 3655 19672 3700 19700
rect 3694 19660 3700 19672
rect 3752 19660 3758 19712
rect 4154 19660 4160 19712
rect 4212 19700 4218 19712
rect 4525 19703 4583 19709
rect 4525 19700 4537 19703
rect 4212 19672 4537 19700
rect 4212 19660 4218 19672
rect 4525 19669 4537 19672
rect 4571 19669 4583 19703
rect 4525 19663 4583 19669
rect 4798 19660 4804 19712
rect 4856 19700 4862 19712
rect 5184 19700 5212 19799
rect 5442 19796 5448 19848
rect 5500 19836 5506 19848
rect 5629 19839 5687 19845
rect 5629 19836 5641 19839
rect 5500 19808 5641 19836
rect 5500 19796 5506 19808
rect 5629 19805 5641 19808
rect 5675 19805 5687 19839
rect 5629 19799 5687 19805
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19805 9275 19839
rect 10134 19836 10140 19848
rect 10095 19808 10140 19836
rect 9217 19799 9275 19805
rect 9232 19768 9260 19799
rect 10134 19796 10140 19808
rect 10192 19796 10198 19848
rect 13280 19836 13308 19867
rect 14550 19864 14556 19876
rect 14608 19864 14614 19916
rect 14642 19864 14648 19916
rect 14700 19904 14706 19916
rect 15289 19907 15347 19913
rect 15289 19904 15301 19907
rect 14700 19876 15301 19904
rect 14700 19864 14706 19876
rect 15289 19873 15301 19876
rect 15335 19873 15347 19907
rect 15289 19867 15347 19873
rect 15378 19864 15384 19916
rect 15436 19904 15442 19916
rect 15841 19907 15899 19913
rect 15841 19904 15853 19907
rect 15436 19876 15853 19904
rect 15436 19864 15442 19876
rect 15841 19873 15853 19876
rect 15887 19873 15899 19907
rect 16390 19904 16396 19916
rect 16351 19876 16396 19904
rect 15841 19867 15899 19873
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 16942 19904 16948 19916
rect 16903 19876 16948 19904
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 17696 19913 17724 19944
rect 18874 19932 18880 19944
rect 18932 19932 18938 19984
rect 17681 19907 17739 19913
rect 17681 19873 17693 19907
rect 17727 19873 17739 19907
rect 17681 19867 17739 19873
rect 18138 19864 18144 19916
rect 18196 19904 18202 19916
rect 18417 19907 18475 19913
rect 18417 19904 18429 19907
rect 18196 19876 18429 19904
rect 18196 19864 18202 19876
rect 18417 19873 18429 19876
rect 18463 19873 18475 19907
rect 18417 19867 18475 19873
rect 18969 19907 19027 19913
rect 18969 19873 18981 19907
rect 19015 19873 19027 19907
rect 18969 19867 19027 19873
rect 14182 19836 14188 19848
rect 13280 19808 14188 19836
rect 14182 19796 14188 19808
rect 14240 19796 14246 19848
rect 17957 19839 18015 19845
rect 17957 19805 17969 19839
rect 18003 19836 18015 19839
rect 18984 19836 19012 19867
rect 18003 19808 19012 19836
rect 18003 19805 18015 19808
rect 17957 19799 18015 19805
rect 10042 19768 10048 19780
rect 9232 19740 10048 19768
rect 10042 19728 10048 19740
rect 10100 19728 10106 19780
rect 12897 19771 12955 19777
rect 12897 19737 12909 19771
rect 12943 19768 12955 19771
rect 13998 19768 14004 19780
rect 12943 19740 14004 19768
rect 12943 19737 12955 19740
rect 12897 19731 12955 19737
rect 13998 19728 14004 19740
rect 14056 19728 14062 19780
rect 17678 19728 17684 19780
rect 17736 19768 17742 19780
rect 18601 19771 18659 19777
rect 18601 19768 18613 19771
rect 17736 19740 18613 19768
rect 17736 19728 17742 19740
rect 18601 19737 18613 19740
rect 18647 19737 18659 19771
rect 18601 19731 18659 19737
rect 7009 19703 7067 19709
rect 7009 19700 7021 19703
rect 4856 19672 7021 19700
rect 4856 19660 4862 19672
rect 7009 19669 7021 19672
rect 7055 19669 7067 19703
rect 8294 19700 8300 19712
rect 8255 19672 8300 19700
rect 7009 19663 7067 19669
rect 8294 19660 8300 19672
rect 8352 19660 8358 19712
rect 8573 19703 8631 19709
rect 8573 19669 8585 19703
rect 8619 19700 8631 19703
rect 9030 19700 9036 19712
rect 8619 19672 9036 19700
rect 8619 19669 8631 19672
rect 8573 19663 8631 19669
rect 9030 19660 9036 19672
rect 9088 19660 9094 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 3068 19468 4016 19496
rect 1762 19320 1768 19372
rect 1820 19360 1826 19372
rect 2133 19363 2191 19369
rect 2133 19360 2145 19363
rect 1820 19332 2145 19360
rect 1820 19320 1826 19332
rect 2133 19329 2145 19332
rect 2179 19329 2191 19363
rect 2133 19323 2191 19329
rect 1394 19292 1400 19304
rect 1355 19264 1400 19292
rect 1394 19252 1400 19264
rect 1452 19252 1458 19304
rect 1949 19295 2007 19301
rect 1949 19261 1961 19295
rect 1995 19292 2007 19295
rect 1995 19264 2544 19292
rect 1995 19261 2007 19264
rect 1949 19255 2007 19261
rect 2516 19224 2544 19264
rect 2682 19252 2688 19304
rect 2740 19292 2746 19304
rect 3068 19301 3096 19468
rect 3988 19428 4016 19468
rect 4338 19456 4344 19508
rect 4396 19496 4402 19508
rect 4433 19499 4491 19505
rect 4433 19496 4445 19499
rect 4396 19468 4445 19496
rect 4396 19456 4402 19468
rect 4433 19465 4445 19468
rect 4479 19465 4491 19499
rect 5442 19496 5448 19508
rect 4433 19459 4491 19465
rect 5092 19468 5448 19496
rect 5092 19428 5120 19468
rect 5442 19456 5448 19468
rect 5500 19456 5506 19508
rect 6454 19496 6460 19508
rect 6415 19468 6460 19496
rect 6454 19456 6460 19468
rect 6512 19456 6518 19508
rect 10134 19496 10140 19508
rect 9784 19468 10140 19496
rect 3988 19400 5120 19428
rect 4062 19320 4068 19372
rect 4120 19360 4126 19372
rect 4982 19360 4988 19372
rect 4120 19332 4988 19360
rect 4120 19320 4126 19332
rect 4982 19320 4988 19332
rect 5040 19320 5046 19372
rect 5092 19304 5120 19400
rect 9674 19320 9680 19372
rect 9732 19360 9738 19372
rect 9784 19369 9812 19468
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 14090 19428 14096 19440
rect 11808 19400 14096 19428
rect 11808 19369 11836 19400
rect 14090 19388 14096 19400
rect 14148 19388 14154 19440
rect 9769 19363 9827 19369
rect 9769 19360 9781 19363
rect 9732 19332 9781 19360
rect 9732 19320 9738 19332
rect 9769 19329 9781 19332
rect 9815 19329 9827 19363
rect 9769 19323 9827 19329
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19329 11851 19363
rect 11793 19323 11851 19329
rect 15841 19363 15899 19369
rect 15841 19329 15853 19363
rect 15887 19360 15899 19363
rect 16390 19360 16396 19372
rect 15887 19332 16396 19360
rect 15887 19329 15899 19332
rect 15841 19323 15899 19329
rect 16390 19320 16396 19332
rect 16448 19320 16454 19372
rect 16577 19363 16635 19369
rect 16577 19329 16589 19363
rect 16623 19360 16635 19363
rect 16942 19360 16948 19372
rect 16623 19332 16948 19360
rect 16623 19329 16635 19332
rect 16577 19323 16635 19329
rect 16942 19320 16948 19332
rect 17000 19320 17006 19372
rect 3053 19295 3111 19301
rect 3053 19292 3065 19295
rect 2740 19264 3065 19292
rect 2740 19252 2746 19264
rect 3053 19261 3065 19264
rect 3099 19261 3111 19295
rect 4154 19292 4160 19304
rect 3053 19255 3111 19261
rect 3252 19264 4160 19292
rect 3252 19224 3280 19264
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 4798 19292 4804 19304
rect 4336 19264 4804 19292
rect 2516 19196 3280 19224
rect 3320 19227 3378 19233
rect 3320 19193 3332 19227
rect 3366 19224 3378 19227
rect 4336 19224 4364 19264
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 5074 19292 5080 19304
rect 5035 19264 5080 19292
rect 5074 19252 5080 19264
rect 5132 19252 5138 19304
rect 7374 19292 7380 19304
rect 7335 19264 7380 19292
rect 7374 19252 7380 19264
rect 7432 19252 7438 19304
rect 7644 19295 7702 19301
rect 7644 19261 7656 19295
rect 7690 19292 7702 19295
rect 8754 19292 8760 19304
rect 7690 19264 8760 19292
rect 7690 19261 7702 19264
rect 7644 19255 7702 19261
rect 8754 19252 8760 19264
rect 8812 19252 8818 19304
rect 11238 19252 11244 19304
rect 11296 19292 11302 19304
rect 12618 19301 12624 19304
rect 11517 19295 11575 19301
rect 11517 19292 11529 19295
rect 11296 19264 11529 19292
rect 11296 19252 11302 19264
rect 11517 19261 11529 19264
rect 11563 19261 11575 19295
rect 11517 19255 11575 19261
rect 12560 19295 12624 19301
rect 12560 19261 12572 19295
rect 12606 19261 12624 19295
rect 12560 19255 12624 19261
rect 12618 19252 12624 19255
rect 12676 19252 12682 19304
rect 13354 19292 13360 19304
rect 13315 19264 13360 19292
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19292 13691 19295
rect 14093 19295 14151 19301
rect 14093 19292 14105 19295
rect 13679 19264 14105 19292
rect 13679 19261 13691 19264
rect 13633 19255 13691 19261
rect 14093 19261 14105 19264
rect 14139 19261 14151 19295
rect 14734 19292 14740 19304
rect 14695 19264 14740 19292
rect 14093 19255 14151 19261
rect 14734 19252 14740 19264
rect 14792 19252 14798 19304
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15378 19292 15384 19304
rect 15059 19264 15384 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15378 19252 15384 19264
rect 15436 19252 15442 19304
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19261 15623 19295
rect 16298 19292 16304 19304
rect 16259 19264 16304 19292
rect 15565 19255 15623 19261
rect 3366 19196 4364 19224
rect 5344 19227 5402 19233
rect 3366 19193 3378 19196
rect 3320 19187 3378 19193
rect 5344 19193 5356 19227
rect 5390 19224 5402 19227
rect 6086 19224 6092 19236
rect 5390 19196 6092 19224
rect 5390 19193 5402 19196
rect 5344 19187 5402 19193
rect 6086 19184 6092 19196
rect 6144 19184 6150 19236
rect 10042 19233 10048 19236
rect 10036 19224 10048 19233
rect 10003 19196 10048 19224
rect 10036 19187 10048 19196
rect 10042 19184 10048 19187
rect 10100 19184 10106 19236
rect 12805 19227 12863 19233
rect 12805 19193 12817 19227
rect 12851 19224 12863 19227
rect 14642 19224 14648 19236
rect 12851 19196 14648 19224
rect 12851 19193 12863 19196
rect 12805 19187 12863 19193
rect 14642 19184 14648 19196
rect 14700 19184 14706 19236
rect 15580 19224 15608 19255
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 17034 19292 17040 19304
rect 16995 19264 17040 19292
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 18012 19264 18061 19292
rect 18012 19252 18018 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18325 19295 18383 19301
rect 18325 19261 18337 19295
rect 18371 19292 18383 19295
rect 18785 19295 18843 19301
rect 18785 19292 18797 19295
rect 18371 19264 18797 19292
rect 18371 19261 18383 19264
rect 18325 19255 18383 19261
rect 18785 19261 18797 19264
rect 18831 19261 18843 19295
rect 18785 19255 18843 19261
rect 20533 19295 20591 19301
rect 20533 19261 20545 19295
rect 20579 19292 20591 19295
rect 20714 19292 20720 19304
rect 20579 19264 20720 19292
rect 20579 19261 20591 19264
rect 20533 19255 20591 19261
rect 20714 19252 20720 19264
rect 20772 19252 20778 19304
rect 16574 19224 16580 19236
rect 15580 19196 16580 19224
rect 16574 19184 16580 19196
rect 16632 19184 16638 19236
rect 17313 19227 17371 19233
rect 17313 19193 17325 19227
rect 17359 19224 17371 19227
rect 18230 19224 18236 19236
rect 17359 19196 18236 19224
rect 17359 19193 17371 19196
rect 17313 19187 17371 19193
rect 18230 19184 18236 19196
rect 18288 19184 18294 19236
rect 21174 19224 21180 19236
rect 21135 19196 21180 19224
rect 21174 19184 21180 19196
rect 21232 19184 21238 19236
rect 1670 19116 1676 19168
rect 1728 19156 1734 19168
rect 2590 19156 2596 19168
rect 1728 19128 2596 19156
rect 1728 19116 1734 19128
rect 2590 19116 2596 19128
rect 2648 19116 2654 19168
rect 4522 19116 4528 19168
rect 4580 19156 4586 19168
rect 4801 19159 4859 19165
rect 4801 19156 4813 19159
rect 4580 19128 4813 19156
rect 4580 19116 4586 19128
rect 4801 19125 4813 19128
rect 4847 19156 4859 19159
rect 5258 19156 5264 19168
rect 4847 19128 5264 19156
rect 4847 19125 4859 19128
rect 4801 19119 4859 19125
rect 5258 19116 5264 19128
rect 5316 19116 5322 19168
rect 6730 19116 6736 19168
rect 6788 19156 6794 19168
rect 6825 19159 6883 19165
rect 6825 19156 6837 19159
rect 6788 19128 6837 19156
rect 6788 19116 6794 19128
rect 6825 19125 6837 19128
rect 6871 19125 6883 19159
rect 6825 19119 6883 19125
rect 7742 19116 7748 19168
rect 7800 19156 7806 19168
rect 8757 19159 8815 19165
rect 8757 19156 8769 19159
rect 7800 19128 8769 19156
rect 7800 19116 7806 19128
rect 8757 19125 8769 19128
rect 8803 19125 8815 19159
rect 8757 19119 8815 19125
rect 8938 19116 8944 19168
rect 8996 19156 9002 19168
rect 9309 19159 9367 19165
rect 9309 19156 9321 19159
rect 8996 19128 9321 19156
rect 8996 19116 9002 19128
rect 9309 19125 9321 19128
rect 9355 19125 9367 19159
rect 9309 19119 9367 19125
rect 9766 19116 9772 19168
rect 9824 19156 9830 19168
rect 11149 19159 11207 19165
rect 11149 19156 11161 19159
rect 9824 19128 11161 19156
rect 9824 19116 9830 19128
rect 11149 19125 11161 19128
rect 11195 19125 11207 19159
rect 11149 19119 11207 19125
rect 13078 19116 13084 19168
rect 13136 19156 13142 19168
rect 14277 19159 14335 19165
rect 14277 19156 14289 19159
rect 13136 19128 14289 19156
rect 13136 19116 13142 19128
rect 14277 19125 14289 19128
rect 14323 19125 14335 19159
rect 14277 19119 14335 19125
rect 18046 19116 18052 19168
rect 18104 19156 18110 19168
rect 18969 19159 19027 19165
rect 18969 19156 18981 19159
rect 18104 19128 18981 19156
rect 18104 19116 18110 19128
rect 18969 19125 18981 19128
rect 19015 19125 19027 19159
rect 18969 19119 19027 19125
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 2866 18952 2872 18964
rect 2827 18924 2872 18952
rect 2866 18912 2872 18924
rect 2924 18912 2930 18964
rect 3142 18912 3148 18964
rect 3200 18952 3206 18964
rect 3237 18955 3295 18961
rect 3237 18952 3249 18955
rect 3200 18924 3249 18952
rect 3200 18912 3206 18924
rect 3237 18921 3249 18924
rect 3283 18921 3295 18955
rect 3237 18915 3295 18921
rect 3329 18955 3387 18961
rect 3329 18921 3341 18955
rect 3375 18952 3387 18955
rect 4065 18955 4123 18961
rect 4065 18952 4077 18955
rect 3375 18924 4077 18952
rect 3375 18921 3387 18924
rect 3329 18915 3387 18921
rect 4065 18921 4077 18924
rect 4111 18921 4123 18955
rect 4065 18915 4123 18921
rect 4433 18955 4491 18961
rect 4433 18921 4445 18955
rect 4479 18952 4491 18955
rect 4982 18952 4988 18964
rect 4479 18924 4988 18952
rect 4479 18921 4491 18924
rect 4433 18915 4491 18921
rect 4982 18912 4988 18924
rect 5040 18912 5046 18964
rect 5718 18912 5724 18964
rect 5776 18952 5782 18964
rect 6089 18955 6147 18961
rect 6089 18952 6101 18955
rect 5776 18924 6101 18952
rect 5776 18912 5782 18924
rect 6089 18921 6101 18924
rect 6135 18921 6147 18955
rect 6089 18915 6147 18921
rect 6457 18955 6515 18961
rect 6457 18921 6469 18955
rect 6503 18952 6515 18955
rect 6730 18952 6736 18964
rect 6503 18924 6736 18952
rect 6503 18921 6515 18924
rect 6457 18915 6515 18921
rect 6730 18912 6736 18924
rect 6788 18952 6794 18964
rect 7469 18955 7527 18961
rect 6788 18924 7236 18952
rect 6788 18912 6794 18924
rect 1394 18844 1400 18896
rect 1452 18884 1458 18896
rect 2225 18887 2283 18893
rect 2225 18884 2237 18887
rect 1452 18856 2237 18884
rect 1452 18844 1458 18856
rect 2225 18853 2237 18856
rect 2271 18853 2283 18887
rect 2225 18847 2283 18853
rect 3418 18844 3424 18896
rect 3476 18884 3482 18896
rect 3476 18856 5580 18884
rect 3476 18844 3482 18856
rect 1959 18819 2017 18825
rect 1959 18785 1971 18819
rect 2005 18785 2017 18819
rect 4522 18816 4528 18828
rect 4483 18788 4528 18816
rect 1959 18779 2017 18785
rect 1964 18680 1992 18779
rect 4522 18776 4528 18788
rect 4580 18776 4586 18828
rect 5166 18776 5172 18828
rect 5224 18816 5230 18828
rect 5445 18819 5503 18825
rect 5445 18816 5457 18819
rect 5224 18788 5457 18816
rect 5224 18776 5230 18788
rect 5445 18785 5457 18788
rect 5491 18785 5503 18819
rect 5552 18816 5580 18856
rect 5810 18844 5816 18896
rect 5868 18884 5874 18896
rect 6549 18887 6607 18893
rect 6549 18884 6561 18887
rect 5868 18856 6561 18884
rect 5868 18844 5874 18856
rect 6549 18853 6561 18856
rect 6595 18884 6607 18887
rect 7101 18887 7159 18893
rect 7101 18884 7113 18887
rect 6595 18856 7113 18884
rect 6595 18853 6607 18856
rect 6549 18847 6607 18853
rect 7101 18853 7113 18856
rect 7147 18853 7159 18887
rect 7101 18847 7159 18853
rect 7208 18816 7236 18924
rect 7469 18921 7481 18955
rect 7515 18921 7527 18955
rect 7469 18915 7527 18921
rect 7929 18955 7987 18961
rect 7929 18921 7941 18955
rect 7975 18952 7987 18955
rect 8202 18952 8208 18964
rect 7975 18924 8208 18952
rect 7975 18921 7987 18924
rect 7929 18915 7987 18921
rect 7282 18844 7288 18896
rect 7340 18884 7346 18896
rect 7484 18884 7512 18915
rect 8202 18912 8208 18924
rect 8260 18912 8266 18964
rect 8938 18952 8944 18964
rect 8899 18924 8944 18952
rect 8938 18912 8944 18924
rect 8996 18912 9002 18964
rect 9030 18912 9036 18964
rect 9088 18952 9094 18964
rect 9088 18924 9133 18952
rect 9088 18912 9094 18924
rect 10042 18912 10048 18964
rect 10100 18952 10106 18964
rect 11057 18955 11115 18961
rect 11057 18952 11069 18955
rect 10100 18924 11069 18952
rect 10100 18912 10106 18924
rect 11057 18921 11069 18924
rect 11103 18921 11115 18955
rect 11057 18915 11115 18921
rect 13173 18955 13231 18961
rect 13173 18921 13185 18955
rect 13219 18952 13231 18955
rect 14553 18955 14611 18961
rect 14553 18952 14565 18955
rect 13219 18924 14565 18952
rect 13219 18921 13231 18924
rect 13173 18915 13231 18921
rect 14553 18921 14565 18924
rect 14599 18921 14611 18955
rect 14553 18915 14611 18921
rect 14642 18912 14648 18964
rect 14700 18952 14706 18964
rect 15657 18955 15715 18961
rect 15657 18952 15669 18955
rect 14700 18924 15669 18952
rect 14700 18912 14706 18924
rect 15657 18921 15669 18924
rect 15703 18921 15715 18955
rect 15657 18915 15715 18921
rect 16669 18955 16727 18961
rect 16669 18921 16681 18955
rect 16715 18952 16727 18955
rect 17126 18952 17132 18964
rect 16715 18924 17132 18952
rect 16715 18921 16727 18924
rect 16669 18915 16727 18921
rect 17126 18912 17132 18924
rect 17184 18912 17190 18964
rect 17218 18912 17224 18964
rect 17276 18952 17282 18964
rect 18417 18955 18475 18961
rect 18417 18952 18429 18955
rect 17276 18924 18429 18952
rect 17276 18912 17282 18924
rect 18417 18921 18429 18924
rect 18463 18921 18475 18955
rect 18417 18915 18475 18921
rect 18969 18955 19027 18961
rect 18969 18921 18981 18955
rect 19015 18952 19027 18955
rect 19058 18952 19064 18964
rect 19015 18924 19064 18952
rect 19015 18921 19027 18924
rect 18969 18915 19027 18921
rect 19058 18912 19064 18924
rect 19116 18912 19122 18964
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 21361 18955 21419 18961
rect 21361 18952 21373 18955
rect 20772 18924 21373 18952
rect 20772 18912 20778 18924
rect 21361 18921 21373 18924
rect 21407 18952 21419 18955
rect 22278 18952 22284 18964
rect 21407 18924 22284 18952
rect 21407 18921 21419 18924
rect 21361 18915 21419 18921
rect 22278 18912 22284 18924
rect 22336 18912 22342 18964
rect 8294 18884 8300 18896
rect 7340 18856 7512 18884
rect 7668 18856 8300 18884
rect 7340 18844 7346 18856
rect 7668 18816 7696 18856
rect 8294 18844 8300 18856
rect 8352 18844 8358 18896
rect 10502 18884 10508 18896
rect 9140 18856 10508 18884
rect 7834 18816 7840 18828
rect 5552 18788 6224 18816
rect 5445 18779 5503 18785
rect 3513 18751 3571 18757
rect 3513 18717 3525 18751
rect 3559 18748 3571 18751
rect 3694 18748 3700 18760
rect 3559 18720 3700 18748
rect 3559 18717 3571 18720
rect 3513 18711 3571 18717
rect 3694 18708 3700 18720
rect 3752 18708 3758 18760
rect 4338 18708 4344 18760
rect 4396 18748 4402 18760
rect 4617 18751 4675 18757
rect 4617 18748 4629 18751
rect 4396 18720 4629 18748
rect 4396 18708 4402 18720
rect 4617 18717 4629 18720
rect 4663 18717 4675 18751
rect 5534 18748 5540 18760
rect 5495 18720 5540 18748
rect 4617 18711 4675 18717
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 5721 18751 5779 18757
rect 5721 18717 5733 18751
rect 5767 18748 5779 18751
rect 6086 18748 6092 18760
rect 5767 18720 6092 18748
rect 5767 18717 5779 18720
rect 5721 18711 5779 18717
rect 6086 18708 6092 18720
rect 6144 18708 6150 18760
rect 6196 18748 6224 18788
rect 6564 18788 6776 18816
rect 7208 18788 7696 18816
rect 7795 18788 7840 18816
rect 6564 18748 6592 18788
rect 6196 18720 6592 18748
rect 6641 18751 6699 18757
rect 6641 18717 6653 18751
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 5077 18683 5135 18689
rect 5077 18680 5089 18683
rect 1964 18652 5089 18680
rect 5077 18649 5089 18652
rect 5123 18649 5135 18683
rect 5077 18643 5135 18649
rect 6454 18640 6460 18692
rect 6512 18680 6518 18692
rect 6656 18680 6684 18711
rect 6512 18652 6684 18680
rect 6748 18680 6776 18788
rect 7834 18776 7840 18788
rect 7892 18776 7898 18828
rect 7926 18776 7932 18828
rect 7984 18816 7990 18828
rect 9140 18816 9168 18856
rect 10502 18844 10508 18856
rect 10560 18844 10566 18896
rect 11600 18887 11658 18893
rect 11600 18853 11612 18887
rect 11646 18884 11658 18887
rect 14274 18884 14280 18896
rect 11646 18856 14280 18884
rect 11646 18853 11658 18856
rect 11600 18847 11658 18853
rect 14274 18844 14280 18856
rect 14332 18884 14338 18896
rect 14332 18856 14780 18884
rect 14332 18844 14338 18856
rect 9766 18816 9772 18828
rect 7984 18788 9168 18816
rect 9232 18788 9772 18816
rect 7984 18776 7990 18788
rect 7742 18708 7748 18760
rect 7800 18748 7806 18760
rect 9232 18757 9260 18788
rect 9766 18776 9772 18788
rect 9824 18776 9830 18828
rect 9950 18825 9956 18828
rect 9944 18816 9956 18825
rect 9911 18788 9956 18816
rect 9944 18779 9956 18788
rect 9950 18776 9956 18779
rect 10008 18776 10014 18828
rect 11333 18819 11391 18825
rect 11333 18785 11345 18819
rect 11379 18816 11391 18819
rect 12526 18816 12532 18828
rect 11379 18788 12532 18816
rect 11379 18785 11391 18788
rect 11333 18779 11391 18785
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 13538 18816 13544 18828
rect 13499 18788 13544 18816
rect 13538 18776 13544 18788
rect 13596 18776 13602 18828
rect 8021 18751 8079 18757
rect 8021 18748 8033 18751
rect 7800 18720 8033 18748
rect 7800 18708 7806 18720
rect 8021 18717 8033 18720
rect 8067 18717 8079 18751
rect 8021 18711 8079 18717
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18717 9275 18751
rect 9674 18748 9680 18760
rect 9635 18720 9680 18748
rect 9217 18711 9275 18717
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 12894 18708 12900 18760
rect 12952 18748 12958 18760
rect 13633 18751 13691 18757
rect 13633 18748 13645 18751
rect 12952 18720 13645 18748
rect 12952 18708 12958 18720
rect 13633 18717 13645 18720
rect 13679 18717 13691 18751
rect 13633 18711 13691 18717
rect 13725 18751 13783 18757
rect 13725 18717 13737 18751
rect 13771 18748 13783 18751
rect 14642 18748 14648 18760
rect 13771 18720 14504 18748
rect 14603 18720 14648 18748
rect 13771 18717 13783 18720
rect 13725 18711 13783 18717
rect 14182 18680 14188 18692
rect 6748 18652 8708 18680
rect 6512 18640 6518 18652
rect 2038 18572 2044 18624
rect 2096 18612 2102 18624
rect 7926 18612 7932 18624
rect 2096 18584 7932 18612
rect 2096 18572 2102 18584
rect 7926 18572 7932 18584
rect 7984 18572 7990 18624
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 8573 18615 8631 18621
rect 8573 18612 8585 18615
rect 8352 18584 8585 18612
rect 8352 18572 8358 18584
rect 8573 18581 8585 18584
rect 8619 18581 8631 18615
rect 8680 18612 8708 18652
rect 12544 18652 12848 18680
rect 14143 18652 14188 18680
rect 12544 18612 12572 18652
rect 12710 18612 12716 18624
rect 8680 18584 12572 18612
rect 12671 18584 12716 18612
rect 8573 18575 8631 18581
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 12820 18612 12848 18652
rect 14182 18640 14188 18652
rect 14240 18640 14246 18692
rect 14476 18680 14504 18720
rect 14642 18708 14648 18720
rect 14700 18708 14706 18760
rect 14752 18757 14780 18856
rect 16942 18776 16948 18828
rect 17000 18816 17006 18828
rect 17497 18819 17555 18825
rect 17497 18816 17509 18819
rect 17000 18788 17509 18816
rect 17000 18776 17006 18788
rect 17497 18785 17509 18788
rect 17543 18785 17555 18819
rect 18230 18816 18236 18828
rect 18191 18788 18236 18816
rect 17497 18779 17555 18785
rect 18230 18776 18236 18788
rect 18288 18776 18294 18828
rect 18785 18819 18843 18825
rect 18785 18785 18797 18819
rect 18831 18785 18843 18819
rect 18785 18779 18843 18785
rect 14737 18751 14795 18757
rect 14737 18717 14749 18751
rect 14783 18717 14795 18751
rect 15746 18748 15752 18760
rect 15707 18720 15752 18748
rect 14737 18711 14795 18717
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18717 15991 18751
rect 16758 18748 16764 18760
rect 16719 18720 16764 18748
rect 15933 18711 15991 18717
rect 15378 18680 15384 18692
rect 14476 18652 15384 18680
rect 15378 18640 15384 18652
rect 15436 18640 15442 18692
rect 15948 18680 15976 18711
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18717 16911 18751
rect 16853 18711 16911 18717
rect 17773 18751 17831 18757
rect 17773 18717 17785 18751
rect 17819 18748 17831 18751
rect 18800 18748 18828 18779
rect 17819 18720 18828 18748
rect 17819 18717 17831 18720
rect 17773 18711 17831 18717
rect 16666 18680 16672 18692
rect 15948 18652 16672 18680
rect 16666 18640 16672 18652
rect 16724 18680 16730 18692
rect 16868 18680 16896 18711
rect 16724 18652 16896 18680
rect 16724 18640 16730 18652
rect 14550 18612 14556 18624
rect 12820 18584 14556 18612
rect 14550 18572 14556 18584
rect 14608 18572 14614 18624
rect 15286 18612 15292 18624
rect 15247 18584 15292 18612
rect 15286 18572 15292 18584
rect 15344 18572 15350 18624
rect 15470 18572 15476 18624
rect 15528 18612 15534 18624
rect 16301 18615 16359 18621
rect 16301 18612 16313 18615
rect 15528 18584 16313 18612
rect 15528 18572 15534 18584
rect 16301 18581 16313 18584
rect 16347 18581 16359 18615
rect 16301 18575 16359 18581
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 2332 18380 3924 18408
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18204 1823 18207
rect 1854 18204 1860 18216
rect 1811 18176 1860 18204
rect 1811 18173 1823 18176
rect 1765 18167 1823 18173
rect 1854 18164 1860 18176
rect 1912 18164 1918 18216
rect 2332 18213 2360 18380
rect 3896 18340 3924 18380
rect 4154 18368 4160 18420
rect 4212 18408 4218 18420
rect 4341 18411 4399 18417
rect 4341 18408 4353 18411
rect 4212 18380 4353 18408
rect 4212 18368 4218 18380
rect 4341 18377 4353 18380
rect 4387 18377 4399 18411
rect 4341 18371 4399 18377
rect 4433 18411 4491 18417
rect 4433 18377 4445 18411
rect 4479 18408 4491 18411
rect 12434 18408 12440 18420
rect 4479 18380 12440 18408
rect 4479 18377 4491 18380
rect 4433 18371 4491 18377
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 12805 18411 12863 18417
rect 12805 18377 12817 18411
rect 12851 18408 12863 18411
rect 13630 18408 13636 18420
rect 12851 18380 13636 18408
rect 12851 18377 12863 18380
rect 12805 18371 12863 18377
rect 13630 18368 13636 18380
rect 13688 18368 13694 18420
rect 14274 18408 14280 18420
rect 14235 18380 14280 18408
rect 14274 18368 14280 18380
rect 14332 18368 14338 18420
rect 14642 18368 14648 18420
rect 14700 18408 14706 18420
rect 14829 18411 14887 18417
rect 14829 18408 14841 18411
rect 14700 18380 14841 18408
rect 14700 18368 14706 18380
rect 14829 18377 14841 18380
rect 14875 18377 14887 18411
rect 15378 18408 15384 18420
rect 15291 18380 15384 18408
rect 14829 18371 14887 18377
rect 15378 18368 15384 18380
rect 15436 18408 15442 18420
rect 17221 18411 17279 18417
rect 17221 18408 17233 18411
rect 15436 18380 17233 18408
rect 15436 18368 15442 18380
rect 17221 18377 17233 18380
rect 17267 18377 17279 18411
rect 17221 18371 17279 18377
rect 3896 18312 5028 18340
rect 2682 18232 2688 18284
rect 2740 18272 2746 18284
rect 2961 18275 3019 18281
rect 2961 18272 2973 18275
rect 2740 18244 2973 18272
rect 2740 18232 2746 18244
rect 2961 18241 2973 18244
rect 3007 18241 3019 18275
rect 5000 18272 5028 18312
rect 6086 18300 6092 18352
rect 6144 18340 6150 18352
rect 6457 18343 6515 18349
rect 6457 18340 6469 18343
rect 6144 18312 6469 18340
rect 6144 18300 6150 18312
rect 6457 18309 6469 18312
rect 6503 18309 6515 18343
rect 6457 18303 6515 18309
rect 6546 18300 6552 18352
rect 6604 18340 6610 18352
rect 6604 18312 8616 18340
rect 6604 18300 6610 18312
rect 7193 18275 7251 18281
rect 7193 18272 7205 18275
rect 5000 18244 5212 18272
rect 2961 18235 3019 18241
rect 2317 18207 2375 18213
rect 2317 18173 2329 18207
rect 2363 18173 2375 18207
rect 4433 18207 4491 18213
rect 4433 18204 4445 18207
rect 2317 18167 2375 18173
rect 2424 18176 4445 18204
rect 658 18096 664 18148
rect 716 18136 722 18148
rect 2424 18136 2452 18176
rect 4433 18173 4445 18176
rect 4479 18173 4491 18207
rect 4433 18167 4491 18173
rect 4617 18207 4675 18213
rect 4617 18173 4629 18207
rect 4663 18204 4675 18207
rect 5074 18204 5080 18216
rect 4663 18176 4936 18204
rect 5035 18176 5080 18204
rect 4663 18173 4675 18176
rect 4617 18167 4675 18173
rect 716 18108 2452 18136
rect 3228 18139 3286 18145
rect 716 18096 722 18108
rect 3228 18105 3240 18139
rect 3274 18136 3286 18139
rect 3694 18136 3700 18148
rect 3274 18108 3700 18136
rect 3274 18105 3286 18108
rect 3228 18099 3286 18105
rect 3694 18096 3700 18108
rect 3752 18096 3758 18148
rect 3878 18096 3884 18148
rect 3936 18136 3942 18148
rect 4798 18136 4804 18148
rect 3936 18108 4804 18136
rect 3936 18096 3942 18108
rect 4798 18096 4804 18108
rect 4856 18096 4862 18148
rect 4908 18136 4936 18176
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 5184 18204 5212 18244
rect 6104 18244 7205 18272
rect 6104 18204 6132 18244
rect 7193 18241 7205 18244
rect 7239 18241 7251 18275
rect 7834 18272 7840 18284
rect 7795 18244 7840 18272
rect 7193 18235 7251 18241
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 8588 18281 8616 18312
rect 10410 18300 10416 18352
rect 10468 18340 10474 18352
rect 12529 18343 12587 18349
rect 12529 18340 12541 18343
rect 10468 18312 12541 18340
rect 10468 18300 10474 18312
rect 12529 18309 12541 18312
rect 12575 18340 12587 18343
rect 12894 18340 12900 18352
rect 12575 18312 12900 18340
rect 12575 18309 12587 18312
rect 12529 18303 12587 18309
rect 12894 18300 12900 18312
rect 12952 18300 12958 18352
rect 15396 18340 15424 18368
rect 14844 18312 15424 18340
rect 8573 18275 8631 18281
rect 8573 18241 8585 18275
rect 8619 18241 8631 18275
rect 8573 18235 8631 18241
rect 8662 18232 8668 18284
rect 8720 18272 8726 18284
rect 12342 18272 12348 18284
rect 8720 18244 12348 18272
rect 8720 18232 8726 18244
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 5184 18176 6132 18204
rect 7009 18207 7067 18213
rect 7009 18173 7021 18207
rect 7055 18204 7067 18207
rect 7282 18204 7288 18216
rect 7055 18176 7288 18204
rect 7055 18173 7067 18176
rect 7009 18167 7067 18173
rect 7282 18164 7288 18176
rect 7340 18164 7346 18216
rect 8294 18204 8300 18216
rect 8255 18176 8300 18204
rect 8294 18164 8300 18176
rect 8352 18164 8358 18216
rect 8386 18164 8392 18216
rect 8444 18204 8450 18216
rect 12066 18204 12072 18216
rect 8444 18176 12072 18204
rect 8444 18164 8450 18176
rect 12066 18164 12072 18176
rect 12124 18164 12130 18216
rect 12250 18164 12256 18216
rect 12308 18204 12314 18216
rect 12526 18204 12532 18216
rect 12308 18176 12532 18204
rect 12308 18164 12314 18176
rect 12526 18164 12532 18176
rect 12584 18204 12590 18216
rect 12897 18207 12955 18213
rect 12897 18204 12909 18207
rect 12584 18176 12909 18204
rect 12584 18164 12590 18176
rect 12897 18173 12909 18176
rect 12943 18173 12955 18207
rect 12897 18167 12955 18173
rect 13164 18207 13222 18213
rect 13164 18173 13176 18207
rect 13210 18204 13222 18207
rect 14844 18204 14872 18312
rect 15286 18272 15292 18284
rect 15247 18244 15292 18272
rect 15286 18232 15292 18244
rect 15344 18232 15350 18284
rect 15396 18281 15424 18312
rect 15381 18275 15439 18281
rect 15381 18241 15393 18275
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 18138 18232 18144 18284
rect 18196 18272 18202 18284
rect 18233 18275 18291 18281
rect 18233 18272 18245 18275
rect 18196 18244 18245 18272
rect 18196 18232 18202 18244
rect 18233 18241 18245 18244
rect 18279 18241 18291 18275
rect 18233 18235 18291 18241
rect 13210 18176 14872 18204
rect 15197 18207 15255 18213
rect 13210 18173 13222 18176
rect 13164 18167 13222 18173
rect 15197 18173 15209 18207
rect 15243 18204 15255 18207
rect 15470 18204 15476 18216
rect 15243 18176 15476 18204
rect 15243 18173 15255 18176
rect 15197 18167 15255 18173
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 15841 18207 15899 18213
rect 15841 18173 15853 18207
rect 15887 18173 15899 18207
rect 18046 18204 18052 18216
rect 18007 18176 18052 18204
rect 15841 18167 15899 18173
rect 5166 18136 5172 18148
rect 4908 18108 5172 18136
rect 5166 18096 5172 18108
rect 5224 18096 5230 18148
rect 5344 18139 5402 18145
rect 5344 18105 5356 18139
rect 5390 18136 5402 18139
rect 6178 18136 6184 18148
rect 5390 18108 6184 18136
rect 5390 18105 5402 18108
rect 5344 18099 5402 18105
rect 6178 18096 6184 18108
rect 6236 18096 6242 18148
rect 6288 18108 7687 18136
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 2498 18068 2504 18080
rect 2459 18040 2504 18068
rect 2498 18028 2504 18040
rect 2556 18028 2562 18080
rect 2590 18028 2596 18080
rect 2648 18068 2654 18080
rect 6288 18068 6316 18108
rect 2648 18040 6316 18068
rect 2648 18028 2654 18040
rect 7006 18028 7012 18080
rect 7064 18068 7070 18080
rect 7558 18068 7564 18080
rect 7064 18040 7564 18068
rect 7064 18028 7070 18040
rect 7558 18028 7564 18040
rect 7616 18028 7622 18080
rect 7659 18068 7687 18108
rect 7926 18096 7932 18148
rect 7984 18136 7990 18148
rect 12805 18139 12863 18145
rect 12805 18136 12817 18139
rect 7984 18108 12817 18136
rect 7984 18096 7990 18108
rect 12805 18105 12817 18108
rect 12851 18105 12863 18139
rect 12805 18099 12863 18105
rect 15286 18096 15292 18148
rect 15344 18136 15350 18148
rect 15856 18136 15884 18167
rect 18046 18164 18052 18176
rect 18104 18164 18110 18216
rect 19242 18164 19248 18216
rect 19300 18204 19306 18216
rect 22738 18204 22744 18216
rect 19300 18176 22744 18204
rect 19300 18164 19306 18176
rect 22738 18164 22744 18176
rect 22796 18164 22802 18216
rect 15344 18108 15884 18136
rect 16108 18139 16166 18145
rect 15344 18096 15350 18108
rect 16108 18105 16120 18139
rect 16154 18136 16166 18139
rect 16666 18136 16672 18148
rect 16154 18108 16672 18136
rect 16154 18105 16166 18108
rect 16108 18099 16166 18105
rect 16666 18096 16672 18108
rect 16724 18096 16730 18148
rect 21174 18136 21180 18148
rect 16776 18108 21180 18136
rect 8386 18068 8392 18080
rect 7659 18040 8392 18068
rect 8386 18028 8392 18040
rect 8444 18028 8450 18080
rect 10870 18028 10876 18080
rect 10928 18068 10934 18080
rect 16776 18068 16804 18108
rect 21174 18096 21180 18108
rect 21232 18096 21238 18148
rect 10928 18040 16804 18068
rect 10928 18028 10934 18040
rect 17218 18028 17224 18080
rect 17276 18068 17282 18080
rect 17497 18071 17555 18077
rect 17497 18068 17509 18071
rect 17276 18040 17509 18068
rect 17276 18028 17282 18040
rect 17497 18037 17509 18040
rect 17543 18037 17555 18071
rect 17497 18031 17555 18037
rect 20990 18028 20996 18080
rect 21048 18068 21054 18080
rect 21818 18068 21824 18080
rect 21048 18040 21824 18068
rect 21048 18028 21054 18040
rect 21818 18028 21824 18040
rect 21876 18028 21882 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 1762 17864 1768 17876
rect 1723 17836 1768 17864
rect 1762 17824 1768 17836
rect 1820 17824 1826 17876
rect 2958 17824 2964 17876
rect 3016 17864 3022 17876
rect 3053 17867 3111 17873
rect 3053 17864 3065 17867
rect 3016 17836 3065 17864
rect 3016 17824 3022 17836
rect 3053 17833 3065 17836
rect 3099 17833 3111 17867
rect 3053 17827 3111 17833
rect 4525 17867 4583 17873
rect 4525 17833 4537 17867
rect 4571 17864 4583 17867
rect 4890 17864 4896 17876
rect 4571 17836 4896 17864
rect 4571 17833 4583 17836
rect 4525 17827 4583 17833
rect 4890 17824 4896 17836
rect 4948 17864 4954 17876
rect 5077 17867 5135 17873
rect 5077 17864 5089 17867
rect 4948 17836 5089 17864
rect 4948 17824 4954 17836
rect 5077 17833 5089 17836
rect 5123 17833 5135 17867
rect 5077 17827 5135 17833
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 5629 17867 5687 17873
rect 5629 17864 5641 17867
rect 5592 17836 5641 17864
rect 5592 17824 5598 17836
rect 5629 17833 5641 17836
rect 5675 17833 5687 17867
rect 5629 17827 5687 17833
rect 6089 17867 6147 17873
rect 6089 17833 6101 17867
rect 6135 17864 6147 17867
rect 6270 17864 6276 17876
rect 6135 17836 6276 17864
rect 6135 17833 6147 17836
rect 6089 17827 6147 17833
rect 6270 17824 6276 17836
rect 6328 17864 6334 17876
rect 6641 17867 6699 17873
rect 6641 17864 6653 17867
rect 6328 17836 6653 17864
rect 6328 17824 6334 17836
rect 6641 17833 6653 17836
rect 6687 17833 6699 17867
rect 6641 17827 6699 17833
rect 8573 17867 8631 17873
rect 8573 17833 8585 17867
rect 8619 17833 8631 17867
rect 8573 17827 8631 17833
rect 11333 17867 11391 17873
rect 11333 17833 11345 17867
rect 11379 17864 11391 17867
rect 11974 17864 11980 17876
rect 11379 17836 11980 17864
rect 11379 17833 11391 17836
rect 11333 17827 11391 17833
rect 2038 17756 2044 17808
rect 2096 17796 2102 17808
rect 8588 17796 8616 17827
rect 11974 17824 11980 17836
rect 12032 17824 12038 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 12894 17864 12900 17876
rect 12492 17836 12900 17864
rect 12492 17824 12498 17836
rect 12894 17824 12900 17836
rect 12952 17864 12958 17876
rect 13538 17864 13544 17876
rect 12952 17836 13400 17864
rect 13499 17836 13544 17864
rect 12952 17824 12958 17836
rect 2096 17768 8616 17796
rect 9944 17799 10002 17805
rect 2096 17756 2102 17768
rect 9944 17765 9956 17799
rect 9990 17796 10002 17799
rect 10042 17796 10048 17808
rect 9990 17768 10048 17796
rect 9990 17765 10002 17768
rect 9944 17759 10002 17765
rect 10042 17756 10048 17768
rect 10100 17756 10106 17808
rect 10134 17756 10140 17808
rect 10192 17796 10198 17808
rect 11882 17796 11888 17808
rect 10192 17768 11888 17796
rect 10192 17756 10198 17768
rect 11882 17756 11888 17768
rect 11940 17756 11946 17808
rect 12342 17796 12348 17808
rect 12255 17768 12348 17796
rect 12342 17756 12348 17768
rect 12400 17796 12406 17808
rect 12526 17796 12532 17808
rect 12400 17768 12532 17796
rect 12400 17756 12406 17768
rect 12526 17756 12532 17768
rect 12584 17756 12590 17808
rect 13372 17796 13400 17836
rect 13538 17824 13544 17836
rect 13596 17824 13602 17876
rect 14550 17864 14556 17876
rect 14511 17836 14556 17864
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 16666 17864 16672 17876
rect 16627 17836 16672 17864
rect 16666 17824 16672 17836
rect 16724 17824 16730 17876
rect 18046 17824 18052 17876
rect 18104 17864 18110 17876
rect 18141 17867 18199 17873
rect 18141 17864 18153 17867
rect 18104 17836 18153 17864
rect 18104 17824 18110 17836
rect 18141 17833 18153 17836
rect 18187 17833 18199 17867
rect 18141 17827 18199 17833
rect 14829 17799 14887 17805
rect 14829 17796 14841 17799
rect 13372 17768 14841 17796
rect 14829 17765 14841 17768
rect 14875 17796 14887 17799
rect 15746 17796 15752 17808
rect 14875 17768 15752 17796
rect 14875 17765 14887 17768
rect 14829 17759 14887 17765
rect 15746 17756 15752 17768
rect 15804 17756 15810 17808
rect 1578 17728 1584 17740
rect 1539 17700 1584 17728
rect 1578 17688 1584 17700
rect 1636 17688 1642 17740
rect 2130 17728 2136 17740
rect 2091 17700 2136 17728
rect 2130 17688 2136 17700
rect 2188 17688 2194 17740
rect 2409 17731 2467 17737
rect 2409 17697 2421 17731
rect 2455 17728 2467 17731
rect 2869 17731 2927 17737
rect 2869 17728 2881 17731
rect 2455 17700 2881 17728
rect 2455 17697 2467 17700
rect 2409 17691 2467 17697
rect 2869 17697 2881 17700
rect 2915 17697 2927 17731
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 2869 17691 2927 17697
rect 3620 17700 4445 17728
rect 3418 17484 3424 17536
rect 3476 17524 3482 17536
rect 3620 17533 3648 17700
rect 4433 17697 4445 17700
rect 4479 17697 4491 17731
rect 5994 17728 6000 17740
rect 5955 17700 6000 17728
rect 4433 17691 4491 17697
rect 5994 17688 6000 17700
rect 6052 17688 6058 17740
rect 8294 17728 8300 17740
rect 8255 17700 8300 17728
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 8938 17728 8944 17740
rect 8899 17700 8944 17728
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 9674 17728 9680 17740
rect 9140 17700 9680 17728
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4617 17663 4675 17669
rect 4617 17660 4629 17663
rect 4212 17632 4629 17660
rect 4212 17620 4218 17632
rect 4617 17629 4629 17632
rect 4663 17629 4675 17663
rect 4617 17623 4675 17629
rect 6178 17620 6184 17672
rect 6236 17660 6242 17672
rect 7190 17660 7196 17672
rect 6236 17632 6281 17660
rect 7151 17632 7196 17660
rect 6236 17620 6242 17632
rect 7190 17620 7196 17632
rect 7248 17620 7254 17672
rect 9030 17660 9036 17672
rect 8991 17632 9036 17660
rect 9030 17620 9036 17632
rect 9088 17620 9094 17672
rect 3970 17552 3976 17604
rect 4028 17592 4034 17604
rect 4028 17564 7236 17592
rect 4028 17552 4034 17564
rect 3605 17527 3663 17533
rect 3605 17524 3617 17527
rect 3476 17496 3617 17524
rect 3476 17484 3482 17496
rect 3605 17493 3617 17496
rect 3651 17493 3663 17527
rect 4062 17524 4068 17536
rect 4023 17496 4068 17524
rect 3605 17487 3663 17493
rect 4062 17484 4068 17496
rect 4120 17484 4126 17536
rect 7208 17524 7236 17564
rect 7374 17552 7380 17604
rect 7432 17592 7438 17604
rect 8113 17595 8171 17601
rect 8113 17592 8125 17595
rect 7432 17564 8125 17592
rect 7432 17552 7438 17564
rect 8113 17561 8125 17564
rect 8159 17592 8171 17595
rect 8662 17592 8668 17604
rect 8159 17564 8668 17592
rect 8159 17561 8171 17564
rect 8113 17555 8171 17561
rect 8662 17552 8668 17564
rect 8720 17592 8726 17604
rect 9140 17592 9168 17700
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 11698 17728 11704 17740
rect 11659 17700 11704 17728
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 15102 17688 15108 17740
rect 15160 17728 15166 17740
rect 15545 17731 15603 17737
rect 15545 17728 15557 17731
rect 15160 17700 15557 17728
rect 15160 17688 15166 17700
rect 15545 17697 15557 17700
rect 15591 17697 15603 17731
rect 15545 17691 15603 17697
rect 18509 17731 18567 17737
rect 18509 17697 18521 17731
rect 18555 17728 18567 17731
rect 19153 17731 19211 17737
rect 19153 17728 19165 17731
rect 18555 17700 19165 17728
rect 18555 17697 18567 17700
rect 18509 17691 18567 17697
rect 19153 17697 19165 17700
rect 19199 17697 19211 17731
rect 19153 17691 19211 17697
rect 9217 17663 9275 17669
rect 9217 17629 9229 17663
rect 9263 17660 9275 17663
rect 11790 17660 11796 17672
rect 9263 17632 9444 17660
rect 11751 17632 11796 17660
rect 9263 17629 9275 17632
rect 9217 17623 9275 17629
rect 8720 17564 9168 17592
rect 8720 17552 8726 17564
rect 9306 17524 9312 17536
rect 7208 17496 9312 17524
rect 9306 17484 9312 17496
rect 9364 17484 9370 17536
rect 9416 17524 9444 17632
rect 11790 17620 11796 17632
rect 11848 17620 11854 17672
rect 11977 17663 12035 17669
rect 11977 17629 11989 17663
rect 12023 17660 12035 17663
rect 12434 17660 12440 17672
rect 12023 17632 12440 17660
rect 12023 17629 12035 17632
rect 11977 17623 12035 17629
rect 12434 17620 12440 17632
rect 12492 17620 12498 17672
rect 15286 17660 15292 17672
rect 15247 17632 15292 17660
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 18046 17620 18052 17672
rect 18104 17660 18110 17672
rect 18601 17663 18659 17669
rect 18601 17660 18613 17663
rect 18104 17632 18613 17660
rect 18104 17620 18110 17632
rect 18601 17629 18613 17632
rect 18647 17629 18659 17663
rect 18782 17660 18788 17672
rect 18743 17632 18788 17660
rect 18601 17623 18659 17629
rect 18782 17620 18788 17632
rect 18840 17620 18846 17672
rect 9950 17524 9956 17536
rect 9416 17496 9956 17524
rect 9950 17484 9956 17496
rect 10008 17524 10014 17536
rect 11057 17527 11115 17533
rect 11057 17524 11069 17527
rect 10008 17496 11069 17524
rect 10008 17484 10014 17496
rect 11057 17493 11069 17496
rect 11103 17493 11115 17527
rect 11057 17487 11115 17493
rect 12805 17527 12863 17533
rect 12805 17493 12817 17527
rect 12851 17524 12863 17527
rect 13170 17524 13176 17536
rect 12851 17496 13176 17524
rect 12851 17493 12863 17496
rect 12805 17487 12863 17493
rect 13170 17484 13176 17496
rect 13228 17524 13234 17536
rect 14093 17527 14151 17533
rect 14093 17524 14105 17527
rect 13228 17496 14105 17524
rect 13228 17484 13234 17496
rect 14093 17493 14105 17496
rect 14139 17524 14151 17527
rect 14274 17524 14280 17536
rect 14139 17496 14280 17524
rect 14139 17493 14151 17496
rect 14093 17487 14151 17493
rect 14274 17484 14280 17496
rect 14332 17484 14338 17536
rect 16666 17484 16672 17536
rect 16724 17524 16730 17536
rect 16945 17527 17003 17533
rect 16945 17524 16957 17527
rect 16724 17496 16957 17524
rect 16724 17484 16730 17496
rect 16945 17493 16957 17496
rect 16991 17493 17003 17527
rect 16945 17487 17003 17493
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 5074 17320 5080 17332
rect 3528 17292 5080 17320
rect 1578 17212 1584 17264
rect 1636 17252 1642 17264
rect 1636 17224 2360 17252
rect 1636 17212 1642 17224
rect 2225 17187 2283 17193
rect 2225 17184 2237 17187
rect 1504 17156 2237 17184
rect 1504 17125 1532 17156
rect 2225 17153 2237 17156
rect 2271 17153 2283 17187
rect 2332 17184 2360 17224
rect 3528 17193 3556 17292
rect 4816 17264 4844 17292
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 7374 17320 7380 17332
rect 7116 17292 7380 17320
rect 4798 17212 4804 17264
rect 4856 17212 4862 17264
rect 2961 17187 3019 17193
rect 2961 17184 2973 17187
rect 2332 17156 2973 17184
rect 2225 17147 2283 17153
rect 2961 17153 2973 17156
rect 3007 17153 3019 17187
rect 2961 17147 3019 17153
rect 3513 17187 3571 17193
rect 3513 17153 3525 17187
rect 3559 17153 3571 17187
rect 3513 17147 3571 17153
rect 6914 17144 6920 17196
rect 6972 17184 6978 17196
rect 7116 17193 7144 17292
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 8478 17280 8484 17332
rect 8536 17320 8542 17332
rect 8757 17323 8815 17329
rect 8757 17320 8769 17323
rect 8536 17292 8769 17320
rect 8536 17280 8542 17292
rect 8757 17289 8769 17292
rect 8803 17289 8815 17323
rect 8757 17283 8815 17289
rect 9030 17280 9036 17332
rect 9088 17320 9094 17332
rect 9125 17323 9183 17329
rect 9125 17320 9137 17323
rect 9088 17292 9137 17320
rect 9088 17280 9094 17292
rect 9125 17289 9137 17292
rect 9171 17289 9183 17323
rect 9125 17283 9183 17289
rect 11333 17323 11391 17329
rect 11333 17289 11345 17323
rect 11379 17320 11391 17323
rect 11790 17320 11796 17332
rect 11379 17292 11796 17320
rect 11379 17289 11391 17292
rect 11333 17283 11391 17289
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 11974 17280 11980 17332
rect 12032 17320 12038 17332
rect 12250 17320 12256 17332
rect 12032 17292 12256 17320
rect 12032 17280 12038 17292
rect 12250 17280 12256 17292
rect 12308 17320 12314 17332
rect 13449 17323 13507 17329
rect 13449 17320 13461 17323
rect 12308 17292 13461 17320
rect 12308 17280 12314 17292
rect 13449 17289 13461 17292
rect 13495 17289 13507 17323
rect 13449 17283 13507 17289
rect 16945 17323 17003 17329
rect 16945 17289 16957 17323
rect 16991 17320 17003 17323
rect 17034 17320 17040 17332
rect 16991 17292 17040 17320
rect 16991 17289 17003 17292
rect 16945 17283 17003 17289
rect 8938 17212 8944 17264
rect 8996 17252 9002 17264
rect 8996 17224 10180 17252
rect 8996 17212 9002 17224
rect 7101 17187 7159 17193
rect 7101 17184 7113 17187
rect 6972 17156 7113 17184
rect 6972 17144 6978 17156
rect 7101 17153 7113 17156
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 9769 17187 9827 17193
rect 9769 17153 9781 17187
rect 9815 17184 9827 17187
rect 10042 17184 10048 17196
rect 9815 17156 10048 17184
rect 9815 17153 9827 17156
rect 9769 17147 9827 17153
rect 10042 17144 10048 17156
rect 10100 17144 10106 17196
rect 10152 17193 10180 17224
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17153 10195 17187
rect 10137 17147 10195 17153
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 1489 17119 1547 17125
rect 1489 17085 1501 17119
rect 1535 17085 1547 17119
rect 2038 17116 2044 17128
rect 1999 17088 2044 17116
rect 1489 17079 1547 17085
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17116 2835 17119
rect 3142 17116 3148 17128
rect 2823 17088 3148 17116
rect 2823 17085 2835 17088
rect 2777 17079 2835 17085
rect 3142 17076 3148 17088
rect 3200 17076 3206 17128
rect 3780 17119 3838 17125
rect 3780 17085 3792 17119
rect 3826 17116 3838 17119
rect 4154 17116 4160 17128
rect 3826 17088 4160 17116
rect 3826 17085 3838 17088
rect 3780 17079 3838 17085
rect 4154 17076 4160 17088
rect 4212 17076 4218 17128
rect 7368 17119 7426 17125
rect 7368 17085 7380 17119
rect 7414 17116 7426 17119
rect 7742 17116 7748 17128
rect 7414 17088 7748 17116
rect 7414 17085 7426 17088
rect 7368 17079 7426 17085
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 8846 17116 8852 17128
rect 7944 17088 8852 17116
rect 1670 16980 1676 16992
rect 1631 16952 1676 16980
rect 1670 16940 1676 16952
rect 1728 16940 1734 16992
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 4893 16983 4951 16989
rect 4893 16980 4905 16983
rect 4212 16952 4905 16980
rect 4212 16940 4218 16952
rect 4893 16949 4905 16952
rect 4939 16949 4951 16983
rect 4893 16943 4951 16949
rect 5537 16983 5595 16989
rect 5537 16949 5549 16983
rect 5583 16980 5595 16983
rect 5994 16980 6000 16992
rect 5583 16952 6000 16980
rect 5583 16949 5595 16952
rect 5537 16943 5595 16949
rect 5994 16940 6000 16952
rect 6052 16980 6058 16992
rect 7944 16980 7972 17088
rect 8846 17076 8852 17088
rect 8904 17076 8910 17128
rect 9585 17119 9643 17125
rect 9585 17085 9597 17119
rect 9631 17116 9643 17119
rect 9858 17116 9864 17128
rect 9631 17088 9864 17116
rect 9631 17085 9643 17088
rect 9585 17079 9643 17085
rect 9858 17076 9864 17088
rect 9916 17116 9922 17128
rect 10597 17119 10655 17125
rect 10597 17116 10609 17119
rect 9916 17088 10609 17116
rect 9916 17076 9922 17088
rect 10597 17085 10609 17088
rect 10643 17085 10655 17119
rect 10597 17079 10655 17085
rect 11057 17119 11115 17125
rect 11057 17085 11069 17119
rect 11103 17116 11115 17119
rect 11882 17116 11888 17128
rect 11103 17088 11888 17116
rect 11103 17085 11115 17088
rect 11057 17079 11115 17085
rect 11882 17076 11888 17088
rect 11940 17076 11946 17128
rect 11992 17116 12020 17147
rect 12250 17144 12256 17196
rect 12308 17184 12314 17196
rect 12526 17184 12532 17196
rect 12308 17156 12532 17184
rect 12308 17144 12314 17156
rect 12342 17116 12348 17128
rect 11992 17088 12348 17116
rect 12342 17076 12348 17088
rect 12400 17076 12406 17128
rect 12443 17116 12471 17156
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 12710 17144 12716 17196
rect 12768 17184 12774 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 12768 17156 13001 17184
rect 12768 17144 12774 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 13464 17184 13492 17283
rect 17034 17280 17040 17292
rect 17092 17280 17098 17332
rect 13722 17184 13728 17196
rect 13464 17156 13728 17184
rect 12989 17147 13047 17153
rect 13722 17144 13728 17156
rect 13780 17184 13786 17196
rect 14185 17187 14243 17193
rect 14185 17184 14197 17187
rect 13780 17156 14197 17184
rect 13780 17144 13786 17156
rect 14185 17153 14197 17156
rect 14231 17153 14243 17187
rect 14185 17147 14243 17153
rect 17589 17187 17647 17193
rect 17589 17153 17601 17187
rect 17635 17184 17647 17187
rect 17770 17184 17776 17196
rect 17635 17156 17776 17184
rect 17635 17153 17647 17156
rect 17589 17147 17647 17153
rect 17770 17144 17776 17156
rect 17828 17144 17834 17196
rect 13633 17119 13691 17125
rect 12443 17088 12940 17116
rect 11701 17051 11759 17057
rect 11701 17017 11713 17051
rect 11747 17048 11759 17051
rect 12526 17048 12532 17060
rect 11747 17020 12532 17048
rect 11747 17017 11759 17020
rect 11701 17011 11759 17017
rect 12526 17008 12532 17020
rect 12584 17008 12590 17060
rect 12912 17057 12940 17088
rect 13633 17085 13645 17119
rect 13679 17116 13691 17119
rect 14090 17116 14096 17128
rect 13679 17088 14096 17116
rect 13679 17085 13691 17088
rect 13633 17079 13691 17085
rect 14090 17076 14096 17088
rect 14148 17076 14154 17128
rect 18138 17116 18144 17128
rect 18099 17088 18144 17116
rect 18138 17076 18144 17088
rect 18196 17076 18202 17128
rect 12897 17051 12955 17057
rect 12897 17017 12909 17051
rect 12943 17048 12955 17051
rect 13998 17048 14004 17060
rect 12943 17020 14004 17048
rect 12943 17017 12955 17020
rect 12897 17011 12955 17017
rect 13998 17008 14004 17020
rect 14056 17008 14062 17060
rect 14452 17051 14510 17057
rect 14452 17017 14464 17051
rect 14498 17048 14510 17051
rect 14642 17048 14648 17060
rect 14498 17020 14648 17048
rect 14498 17017 14510 17020
rect 14452 17011 14510 17017
rect 14642 17008 14648 17020
rect 14700 17008 14706 17060
rect 15102 17008 15108 17060
rect 15160 17008 15166 17060
rect 18408 17051 18466 17057
rect 18408 17017 18420 17051
rect 18454 17048 18466 17051
rect 18598 17048 18604 17060
rect 18454 17020 18604 17048
rect 18454 17017 18466 17020
rect 18408 17011 18466 17017
rect 18598 17008 18604 17020
rect 18656 17008 18662 17060
rect 6052 16952 7972 16980
rect 6052 16940 6058 16952
rect 8202 16940 8208 16992
rect 8260 16980 8266 16992
rect 8481 16983 8539 16989
rect 8481 16980 8493 16983
rect 8260 16952 8493 16980
rect 8260 16940 8266 16952
rect 8481 16949 8493 16952
rect 8527 16949 8539 16983
rect 9490 16980 9496 16992
rect 9451 16952 9496 16980
rect 8481 16943 8539 16949
rect 9490 16940 9496 16952
rect 9548 16940 9554 16992
rect 11793 16983 11851 16989
rect 11793 16949 11805 16983
rect 11839 16980 11851 16983
rect 12437 16983 12495 16989
rect 12437 16980 12449 16983
rect 11839 16952 12449 16980
rect 11839 16949 11851 16952
rect 11793 16943 11851 16949
rect 12437 16949 12449 16952
rect 12483 16949 12495 16983
rect 12437 16943 12495 16949
rect 12805 16983 12863 16989
rect 12805 16949 12817 16983
rect 12851 16980 12863 16983
rect 13170 16980 13176 16992
rect 12851 16952 13176 16980
rect 12851 16949 12863 16952
rect 12805 16943 12863 16949
rect 13170 16940 13176 16952
rect 13228 16940 13234 16992
rect 14182 16940 14188 16992
rect 14240 16980 14246 16992
rect 15120 16980 15148 17008
rect 15565 16983 15623 16989
rect 15565 16980 15577 16983
rect 14240 16952 15577 16980
rect 14240 16940 14246 16952
rect 15565 16949 15577 16952
rect 15611 16949 15623 16983
rect 17310 16980 17316 16992
rect 17271 16952 17316 16980
rect 15565 16943 15623 16949
rect 17310 16940 17316 16952
rect 17368 16940 17374 16992
rect 17402 16940 17408 16992
rect 17460 16980 17466 16992
rect 17460 16952 17505 16980
rect 17460 16940 17466 16952
rect 18782 16940 18788 16992
rect 18840 16980 18846 16992
rect 19521 16983 19579 16989
rect 19521 16980 19533 16983
rect 18840 16952 19533 16980
rect 18840 16940 18846 16952
rect 19521 16949 19533 16952
rect 19567 16949 19579 16983
rect 19521 16943 19579 16949
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 1949 16779 2007 16785
rect 1949 16745 1961 16779
rect 1995 16745 2007 16779
rect 1949 16739 2007 16745
rect 1964 16708 1992 16739
rect 2130 16736 2136 16788
rect 2188 16776 2194 16788
rect 2961 16779 3019 16785
rect 2961 16776 2973 16779
rect 2188 16748 2973 16776
rect 2188 16736 2194 16748
rect 2961 16745 2973 16748
rect 3007 16745 3019 16779
rect 2961 16739 3019 16745
rect 3421 16779 3479 16785
rect 3421 16745 3433 16779
rect 3467 16776 3479 16779
rect 4062 16776 4068 16788
rect 3467 16748 4068 16776
rect 3467 16745 3479 16748
rect 3421 16739 3479 16745
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 6178 16736 6184 16788
rect 6236 16776 6242 16788
rect 6273 16779 6331 16785
rect 6273 16776 6285 16779
rect 6236 16748 6285 16776
rect 6236 16736 6242 16748
rect 6273 16745 6285 16748
rect 6319 16745 6331 16779
rect 6273 16739 6331 16745
rect 7190 16736 7196 16788
rect 7248 16776 7254 16788
rect 8941 16779 8999 16785
rect 8941 16776 8953 16779
rect 7248 16748 8953 16776
rect 7248 16736 7254 16748
rect 8941 16745 8953 16748
rect 8987 16745 8999 16779
rect 8941 16739 8999 16745
rect 9306 16736 9312 16788
rect 9364 16776 9370 16788
rect 10226 16776 10232 16788
rect 9364 16748 10232 16776
rect 9364 16736 9370 16748
rect 10226 16736 10232 16748
rect 10284 16736 10290 16788
rect 11146 16736 11152 16788
rect 11204 16776 11210 16788
rect 12342 16776 12348 16788
rect 11204 16748 12348 16776
rect 11204 16736 11210 16748
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 12897 16779 12955 16785
rect 12897 16745 12909 16779
rect 12943 16776 12955 16779
rect 13354 16776 13360 16788
rect 12943 16748 13360 16776
rect 12943 16745 12955 16748
rect 12897 16739 12955 16745
rect 13354 16736 13360 16748
rect 13412 16736 13418 16788
rect 13998 16736 14004 16788
rect 14056 16776 14062 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 14056 16748 14381 16776
rect 14056 16736 14062 16748
rect 14369 16745 14381 16748
rect 14415 16776 14427 16779
rect 15289 16779 15347 16785
rect 15289 16776 15301 16779
rect 14415 16748 15301 16776
rect 14415 16745 14427 16748
rect 14369 16739 14427 16745
rect 15289 16745 15301 16748
rect 15335 16745 15347 16779
rect 17770 16776 17776 16788
rect 17731 16748 17776 16776
rect 15289 16739 15347 16745
rect 17770 16736 17776 16748
rect 17828 16736 17834 16788
rect 18598 16736 18604 16788
rect 18656 16776 18662 16788
rect 19429 16779 19487 16785
rect 19429 16776 19441 16779
rect 18656 16748 19441 16776
rect 18656 16736 18662 16748
rect 19429 16745 19441 16748
rect 19475 16745 19487 16779
rect 19429 16739 19487 16745
rect 3050 16708 3056 16720
rect 1964 16680 3056 16708
rect 3050 16668 3056 16680
rect 3108 16668 3114 16720
rect 3142 16668 3148 16720
rect 3200 16708 3206 16720
rect 11232 16711 11290 16717
rect 3200 16680 8340 16708
rect 3200 16668 3206 16680
rect 1765 16643 1823 16649
rect 1765 16609 1777 16643
rect 1811 16640 1823 16643
rect 2222 16640 2228 16652
rect 1811 16612 2228 16640
rect 1811 16609 1823 16612
rect 1765 16603 1823 16609
rect 2222 16600 2228 16612
rect 2280 16600 2286 16652
rect 3329 16643 3387 16649
rect 3329 16609 3341 16643
rect 3375 16640 3387 16643
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 3375 16612 4077 16640
rect 3375 16609 3387 16612
rect 3329 16603 3387 16609
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 5160 16643 5218 16649
rect 5160 16609 5172 16643
rect 5206 16640 5218 16643
rect 5442 16640 5448 16652
rect 5206 16612 5448 16640
rect 5206 16609 5218 16612
rect 5160 16603 5218 16609
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 6914 16640 6920 16652
rect 6875 16612 6920 16640
rect 6914 16600 6920 16612
rect 6972 16600 6978 16652
rect 7184 16643 7242 16649
rect 7184 16609 7196 16643
rect 7230 16640 7242 16643
rect 8202 16640 8208 16652
rect 7230 16612 8208 16640
rect 7230 16609 7242 16612
rect 7184 16603 7242 16609
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 8312 16640 8340 16680
rect 11232 16677 11244 16711
rect 11278 16708 11290 16711
rect 12710 16708 12716 16720
rect 11278 16680 12716 16708
rect 11278 16677 11290 16680
rect 11232 16671 11290 16677
rect 12710 16668 12716 16680
rect 12768 16668 12774 16720
rect 13265 16711 13323 16717
rect 13265 16677 13277 16711
rect 13311 16708 13323 16711
rect 13906 16708 13912 16720
rect 13311 16680 13912 16708
rect 13311 16677 13323 16680
rect 13265 16671 13323 16677
rect 13906 16668 13912 16680
rect 13964 16668 13970 16720
rect 16660 16711 16718 16717
rect 16660 16677 16672 16711
rect 16706 16708 16718 16711
rect 16758 16708 16764 16720
rect 16706 16680 16764 16708
rect 16706 16677 16718 16680
rect 16660 16671 16718 16677
rect 16758 16668 16764 16680
rect 16816 16668 16822 16720
rect 17788 16708 17816 16736
rect 18294 16711 18352 16717
rect 18294 16708 18306 16711
rect 17788 16680 18306 16708
rect 18294 16677 18306 16680
rect 18340 16677 18352 16711
rect 18294 16671 18352 16677
rect 8312 16612 8616 16640
rect 3605 16575 3663 16581
rect 3605 16541 3617 16575
rect 3651 16572 3663 16575
rect 4154 16572 4160 16584
rect 3651 16544 4160 16572
rect 3651 16541 3663 16544
rect 3605 16535 3663 16541
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 4798 16532 4804 16584
rect 4856 16572 4862 16584
rect 4893 16575 4951 16581
rect 4893 16572 4905 16575
rect 4856 16544 4905 16572
rect 4856 16532 4862 16544
rect 4893 16541 4905 16544
rect 4939 16541 4951 16575
rect 4893 16535 4951 16541
rect 8588 16513 8616 16612
rect 8846 16600 8852 16652
rect 8904 16640 8910 16652
rect 9490 16640 9496 16652
rect 8904 16612 9496 16640
rect 8904 16600 8910 16612
rect 9490 16600 9496 16612
rect 9548 16640 9554 16652
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 9548 16612 9689 16640
rect 9548 16600 9554 16612
rect 9677 16609 9689 16612
rect 9723 16609 9735 16643
rect 10594 16640 10600 16652
rect 10555 16612 10600 16640
rect 9677 16603 9735 16609
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 10962 16640 10968 16652
rect 10875 16612 10968 16640
rect 10962 16600 10968 16612
rect 11020 16640 11026 16652
rect 11974 16640 11980 16652
rect 11020 16612 11980 16640
rect 11020 16600 11026 16612
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 13357 16643 13415 16649
rect 13357 16609 13369 16643
rect 13403 16640 13415 16643
rect 13998 16640 14004 16652
rect 13403 16612 14004 16640
rect 13403 16609 13415 16612
rect 13357 16603 13415 16609
rect 13998 16600 14004 16612
rect 14056 16600 14062 16652
rect 14274 16640 14280 16652
rect 14235 16612 14280 16640
rect 14274 16600 14280 16612
rect 14332 16600 14338 16652
rect 15286 16600 15292 16652
rect 15344 16640 15350 16652
rect 16393 16643 16451 16649
rect 16393 16640 16405 16643
rect 15344 16612 16405 16640
rect 15344 16600 15350 16612
rect 16393 16609 16405 16612
rect 16439 16640 16451 16643
rect 18049 16643 18107 16649
rect 18049 16640 18061 16643
rect 16439 16612 18061 16640
rect 16439 16609 16451 16612
rect 16393 16603 16451 16609
rect 18049 16609 18061 16612
rect 18095 16640 18107 16643
rect 18138 16640 18144 16652
rect 18095 16612 18144 16640
rect 18095 16609 18107 16612
rect 18049 16603 18107 16609
rect 18138 16600 18144 16612
rect 18196 16600 18202 16652
rect 9030 16572 9036 16584
rect 8991 16544 9036 16572
rect 9030 16532 9036 16544
rect 9088 16532 9094 16584
rect 9125 16575 9183 16581
rect 9125 16541 9137 16575
rect 9171 16541 9183 16575
rect 9125 16535 9183 16541
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16572 13599 16575
rect 14182 16572 14188 16584
rect 13587 16544 14188 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 8573 16507 8631 16513
rect 8573 16473 8585 16507
rect 8619 16473 8631 16507
rect 9140 16504 9168 16535
rect 14182 16532 14188 16544
rect 14240 16532 14246 16584
rect 14553 16575 14611 16581
rect 14553 16541 14565 16575
rect 14599 16572 14611 16575
rect 15194 16572 15200 16584
rect 14599 16544 15200 16572
rect 14599 16541 14611 16544
rect 14553 16535 14611 16541
rect 15194 16532 15200 16544
rect 15252 16572 15258 16584
rect 16022 16572 16028 16584
rect 15252 16544 16028 16572
rect 15252 16532 15258 16544
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 8573 16467 8631 16473
rect 9048 16476 9168 16504
rect 8297 16439 8355 16445
rect 8297 16405 8309 16439
rect 8343 16436 8355 16439
rect 8386 16436 8392 16448
rect 8343 16408 8392 16436
rect 8343 16405 8355 16408
rect 8297 16399 8355 16405
rect 8386 16396 8392 16408
rect 8444 16436 8450 16448
rect 9048 16436 9076 16476
rect 8444 16408 9076 16436
rect 13909 16439 13967 16445
rect 8444 16396 8450 16408
rect 13909 16405 13921 16439
rect 13955 16436 13967 16439
rect 14550 16436 14556 16448
rect 13955 16408 14556 16436
rect 13955 16405 13967 16408
rect 13909 16399 13967 16405
rect 14550 16396 14556 16408
rect 14608 16396 14614 16448
rect 15654 16436 15660 16448
rect 15615 16408 15660 16436
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 1670 16232 1676 16244
rect 1631 16204 1676 16232
rect 1670 16192 1676 16204
rect 1728 16192 1734 16244
rect 7377 16235 7435 16241
rect 7377 16201 7389 16235
rect 7423 16232 7435 16235
rect 9030 16232 9036 16244
rect 7423 16204 9036 16232
rect 7423 16201 7435 16204
rect 7377 16195 7435 16201
rect 9030 16192 9036 16204
rect 9088 16192 9094 16244
rect 10042 16232 10048 16244
rect 10003 16204 10048 16232
rect 10042 16192 10048 16204
rect 10100 16192 10106 16244
rect 10321 16235 10379 16241
rect 10321 16201 10333 16235
rect 10367 16232 10379 16235
rect 11698 16232 11704 16244
rect 10367 16204 11704 16232
rect 10367 16201 10379 16204
rect 10321 16195 10379 16201
rect 11698 16192 11704 16204
rect 11756 16192 11762 16244
rect 12437 16235 12495 16241
rect 12437 16201 12449 16235
rect 12483 16232 12495 16235
rect 12526 16232 12532 16244
rect 12483 16204 12532 16232
rect 12483 16201 12495 16204
rect 12437 16195 12495 16201
rect 12526 16192 12532 16204
rect 12584 16192 12590 16244
rect 14642 16192 14648 16244
rect 14700 16232 14706 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 14700 16204 15025 16232
rect 14700 16192 14706 16204
rect 15013 16201 15025 16204
rect 15059 16201 15071 16235
rect 18046 16232 18052 16244
rect 18007 16204 18052 16232
rect 15013 16195 15071 16201
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 4893 16167 4951 16173
rect 4893 16164 4905 16167
rect 2056 16136 4905 16164
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 16028 1547 16031
rect 1578 16028 1584 16040
rect 1535 16000 1584 16028
rect 1535 15997 1547 16000
rect 1489 15991 1547 15997
rect 1578 15988 1584 16000
rect 1636 15988 1642 16040
rect 2056 16037 2084 16136
rect 4893 16133 4905 16136
rect 4939 16133 4951 16167
rect 4893 16127 4951 16133
rect 10226 16124 10232 16176
rect 10284 16164 10290 16176
rect 16577 16167 16635 16173
rect 10284 16136 11928 16164
rect 10284 16124 10290 16136
rect 2222 16096 2228 16108
rect 2183 16068 2228 16096
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 5442 16096 5448 16108
rect 5403 16068 5448 16096
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 8021 16099 8079 16105
rect 8021 16065 8033 16099
rect 8067 16096 8079 16099
rect 8202 16096 8208 16108
rect 8067 16068 8208 16096
rect 8067 16065 8079 16068
rect 8021 16059 8079 16065
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 8662 16096 8668 16108
rect 8623 16068 8668 16096
rect 8662 16056 8668 16068
rect 8720 16056 8726 16108
rect 10965 16099 11023 16105
rect 10965 16065 10977 16099
rect 11011 16096 11023 16099
rect 11146 16096 11152 16108
rect 11011 16068 11152 16096
rect 11011 16065 11023 16068
rect 10965 16059 11023 16065
rect 11146 16056 11152 16068
rect 11204 16056 11210 16108
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 3418 15988 3424 16040
rect 3476 16028 3482 16040
rect 6365 16031 6423 16037
rect 6365 16028 6377 16031
rect 3476 16000 6377 16028
rect 3476 15988 3482 16000
rect 6365 15997 6377 16000
rect 6411 15997 6423 16031
rect 6365 15991 6423 15997
rect 7009 16031 7067 16037
rect 7009 15997 7021 16031
rect 7055 16028 7067 16031
rect 8294 16028 8300 16040
rect 7055 16000 8300 16028
rect 7055 15997 7067 16000
rect 7009 15991 7067 15997
rect 5261 15963 5319 15969
rect 5261 15929 5273 15963
rect 5307 15960 5319 15963
rect 5905 15963 5963 15969
rect 5905 15960 5917 15963
rect 5307 15932 5917 15960
rect 5307 15929 5319 15932
rect 5261 15923 5319 15929
rect 5905 15929 5917 15932
rect 5951 15929 5963 15963
rect 6380 15960 6408 15991
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 9214 15988 9220 16040
rect 9272 16028 9278 16040
rect 11900 16028 11928 16136
rect 13464 16136 13676 16164
rect 11977 16099 12035 16105
rect 11977 16065 11989 16099
rect 12023 16096 12035 16099
rect 12710 16096 12716 16108
rect 12023 16068 12716 16096
rect 12023 16065 12035 16068
rect 11977 16059 12035 16065
rect 12710 16056 12716 16068
rect 12768 16096 12774 16108
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 12768 16068 13001 16096
rect 12768 16056 12774 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 12805 16031 12863 16037
rect 12805 16028 12817 16031
rect 9272 16000 11836 16028
rect 11900 16000 12817 16028
rect 9272 15988 9278 16000
rect 7745 15963 7803 15969
rect 7745 15960 7757 15963
rect 6380 15932 7757 15960
rect 5905 15923 5963 15929
rect 7745 15929 7757 15932
rect 7791 15929 7803 15963
rect 7745 15923 7803 15929
rect 7837 15963 7895 15969
rect 7837 15929 7849 15963
rect 7883 15960 7895 15963
rect 8478 15960 8484 15972
rect 7883 15932 8484 15960
rect 7883 15929 7895 15932
rect 7837 15923 7895 15929
rect 8478 15920 8484 15932
rect 8536 15920 8542 15972
rect 8932 15963 8990 15969
rect 8932 15929 8944 15963
rect 8978 15960 8990 15963
rect 9398 15960 9404 15972
rect 8978 15932 9404 15960
rect 8978 15929 8990 15932
rect 8932 15923 8990 15929
rect 9398 15920 9404 15932
rect 9456 15920 9462 15972
rect 10594 15920 10600 15972
rect 10652 15960 10658 15972
rect 11701 15963 11759 15969
rect 11701 15960 11713 15963
rect 10652 15932 11713 15960
rect 10652 15920 10658 15932
rect 11701 15929 11713 15932
rect 11747 15929 11759 15963
rect 11808 15960 11836 16000
rect 12805 15997 12817 16000
rect 12851 16028 12863 16031
rect 13464 16028 13492 16136
rect 13648 16096 13676 16136
rect 16577 16133 16589 16167
rect 16623 16164 16635 16167
rect 18138 16164 18144 16176
rect 16623 16136 18144 16164
rect 16623 16133 16635 16136
rect 16577 16127 16635 16133
rect 18138 16124 18144 16136
rect 18196 16124 18202 16176
rect 13648 16068 13768 16096
rect 13630 16028 13636 16040
rect 12851 16000 13492 16028
rect 13591 16000 13636 16028
rect 12851 15997 12863 16000
rect 12805 15991 12863 15997
rect 13630 15988 13636 16000
rect 13688 15988 13694 16040
rect 13740 16028 13768 16068
rect 15654 16056 15660 16108
rect 15712 16096 15718 16108
rect 15749 16099 15807 16105
rect 15749 16096 15761 16099
rect 15712 16068 15761 16096
rect 15712 16056 15718 16068
rect 15749 16065 15761 16068
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 16022 16096 16028 16108
rect 15979 16068 16028 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16096 17095 16099
rect 17310 16096 17316 16108
rect 17083 16068 17316 16096
rect 17083 16065 17095 16068
rect 17037 16059 17095 16065
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 18598 16096 18604 16108
rect 18559 16068 18604 16096
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 13740 16000 15332 16028
rect 13446 15960 13452 15972
rect 11808 15932 13452 15960
rect 11701 15923 11759 15929
rect 13446 15920 13452 15932
rect 13504 15920 13510 15972
rect 13900 15963 13958 15969
rect 13900 15929 13912 15963
rect 13946 15960 13958 15963
rect 15194 15960 15200 15972
rect 13946 15932 15200 15960
rect 13946 15929 13958 15932
rect 13900 15923 13958 15929
rect 15194 15920 15200 15932
rect 15252 15920 15258 15972
rect 15304 15960 15332 16000
rect 15378 15988 15384 16040
rect 15436 16028 15442 16040
rect 16761 16031 16819 16037
rect 16761 16028 16773 16031
rect 15436 16000 16773 16028
rect 15436 15988 15442 16000
rect 16761 15997 16773 16000
rect 16807 15997 16819 16031
rect 16761 15991 16819 15997
rect 15470 15960 15476 15972
rect 15304 15932 15476 15960
rect 15470 15920 15476 15932
rect 15528 15960 15534 15972
rect 15657 15963 15715 15969
rect 15657 15960 15669 15963
rect 15528 15932 15669 15960
rect 15528 15920 15534 15932
rect 15657 15929 15669 15932
rect 15703 15929 15715 15963
rect 15657 15923 15715 15929
rect 5350 15892 5356 15904
rect 5311 15864 5356 15892
rect 5350 15852 5356 15864
rect 5408 15852 5414 15904
rect 6822 15892 6828 15904
rect 6783 15864 6828 15892
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 10686 15892 10692 15904
rect 10647 15864 10692 15892
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 10781 15895 10839 15901
rect 10781 15861 10793 15895
rect 10827 15892 10839 15895
rect 11333 15895 11391 15901
rect 11333 15892 11345 15895
rect 10827 15864 11345 15892
rect 10827 15861 10839 15864
rect 10781 15855 10839 15861
rect 11333 15861 11345 15864
rect 11379 15861 11391 15895
rect 11333 15855 11391 15861
rect 11793 15895 11851 15901
rect 11793 15861 11805 15895
rect 11839 15892 11851 15895
rect 11882 15892 11888 15904
rect 11839 15864 11888 15892
rect 11839 15861 11851 15864
rect 11793 15855 11851 15861
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 12526 15852 12532 15904
rect 12584 15892 12590 15904
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 12584 15864 12909 15892
rect 12584 15852 12590 15864
rect 12897 15861 12909 15864
rect 12943 15892 12955 15895
rect 13538 15892 13544 15904
rect 12943 15864 13544 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 15286 15892 15292 15904
rect 15247 15864 15292 15892
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 17589 15895 17647 15901
rect 17589 15892 17601 15895
rect 17368 15864 17601 15892
rect 17368 15852 17374 15864
rect 17589 15861 17601 15864
rect 17635 15892 17647 15895
rect 18417 15895 18475 15901
rect 18417 15892 18429 15895
rect 17635 15864 18429 15892
rect 17635 15861 17647 15864
rect 17589 15855 17647 15861
rect 18417 15861 18429 15864
rect 18463 15861 18475 15895
rect 18417 15855 18475 15861
rect 18506 15852 18512 15904
rect 18564 15892 18570 15904
rect 18564 15864 18609 15892
rect 18564 15852 18570 15864
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 1673 15691 1731 15697
rect 1673 15657 1685 15691
rect 1719 15688 1731 15691
rect 2774 15688 2780 15700
rect 1719 15660 2780 15688
rect 1719 15657 1731 15660
rect 1673 15651 1731 15657
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 2961 15691 3019 15697
rect 2961 15657 2973 15691
rect 3007 15688 3019 15691
rect 3234 15688 3240 15700
rect 3007 15660 3240 15688
rect 3007 15657 3019 15660
rect 2961 15651 3019 15657
rect 3234 15648 3240 15660
rect 3292 15648 3298 15700
rect 5350 15648 5356 15700
rect 5408 15688 5414 15700
rect 6365 15691 6423 15697
rect 6365 15688 6377 15691
rect 5408 15660 6377 15688
rect 5408 15648 5414 15660
rect 6365 15657 6377 15660
rect 6411 15657 6423 15691
rect 6365 15651 6423 15657
rect 6638 15648 6644 15700
rect 6696 15688 6702 15700
rect 6825 15691 6883 15697
rect 6825 15688 6837 15691
rect 6696 15660 6837 15688
rect 6696 15648 6702 15660
rect 6825 15657 6837 15660
rect 6871 15657 6883 15691
rect 6825 15651 6883 15657
rect 7377 15691 7435 15697
rect 7377 15657 7389 15691
rect 7423 15688 7435 15691
rect 8294 15688 8300 15700
rect 7423 15660 8300 15688
rect 7423 15657 7435 15660
rect 7377 15651 7435 15657
rect 8294 15648 8300 15660
rect 8352 15648 8358 15700
rect 8573 15691 8631 15697
rect 8573 15657 8585 15691
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 9033 15691 9091 15697
rect 9033 15657 9045 15691
rect 9079 15688 9091 15691
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 9079 15660 9689 15688
rect 9079 15657 9091 15660
rect 9033 15651 9091 15657
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 9677 15651 9735 15657
rect 10137 15691 10195 15697
rect 10137 15657 10149 15691
rect 10183 15688 10195 15691
rect 10318 15688 10324 15700
rect 10183 15660 10324 15688
rect 10183 15657 10195 15660
rect 10137 15651 10195 15657
rect 8588 15620 8616 15651
rect 10318 15648 10324 15660
rect 10376 15648 10382 15700
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 12529 15691 12587 15697
rect 12529 15688 12541 15691
rect 10744 15660 12541 15688
rect 10744 15648 10750 15660
rect 12529 15657 12541 15660
rect 12575 15657 12587 15691
rect 13998 15688 14004 15700
rect 13959 15660 14004 15688
rect 12529 15651 12587 15657
rect 13998 15648 14004 15660
rect 14056 15648 14062 15700
rect 14369 15691 14427 15697
rect 14369 15657 14381 15691
rect 14415 15688 14427 15691
rect 15286 15688 15292 15700
rect 14415 15660 15292 15688
rect 14415 15657 14427 15660
rect 14369 15651 14427 15657
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 16209 15691 16267 15697
rect 16209 15657 16221 15691
rect 16255 15688 16267 15691
rect 17402 15688 17408 15700
rect 16255 15660 17408 15688
rect 16255 15657 16267 15660
rect 16209 15651 16267 15657
rect 17402 15648 17408 15660
rect 17460 15648 17466 15700
rect 11146 15629 11152 15632
rect 11140 15620 11152 15629
rect 2056 15592 8616 15620
rect 11107 15592 11152 15620
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15552 1547 15555
rect 1946 15552 1952 15564
rect 1535 15524 1952 15552
rect 1535 15521 1547 15524
rect 1489 15515 1547 15521
rect 1946 15512 1952 15524
rect 2004 15512 2010 15564
rect 2056 15561 2084 15592
rect 11140 15583 11152 15592
rect 11146 15580 11152 15583
rect 11204 15580 11210 15632
rect 14461 15623 14519 15629
rect 14461 15589 14473 15623
rect 14507 15620 14519 15623
rect 14550 15620 14556 15632
rect 14507 15592 14556 15620
rect 14507 15589 14519 15592
rect 14461 15583 14519 15589
rect 14550 15580 14556 15592
rect 14608 15580 14614 15632
rect 18782 15629 18788 15632
rect 17221 15623 17279 15629
rect 17221 15620 17233 15623
rect 16592 15592 17233 15620
rect 2041 15555 2099 15561
rect 2041 15521 2053 15555
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15552 2835 15555
rect 2958 15552 2964 15564
rect 2823 15524 2964 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 4709 15555 4767 15561
rect 4709 15521 4721 15555
rect 4755 15552 4767 15555
rect 4798 15552 4804 15564
rect 4755 15524 4804 15552
rect 4755 15521 4767 15524
rect 4709 15515 4767 15521
rect 4798 15512 4804 15524
rect 4856 15512 4862 15564
rect 4976 15555 5034 15561
rect 4976 15521 4988 15555
rect 5022 15552 5034 15555
rect 5022 15524 5948 15552
rect 5022 15521 5034 15524
rect 4976 15515 5034 15521
rect 1578 15444 1584 15496
rect 1636 15484 1642 15496
rect 2225 15487 2283 15493
rect 2225 15484 2237 15487
rect 1636 15456 2237 15484
rect 1636 15444 1642 15456
rect 2225 15453 2237 15456
rect 2271 15453 2283 15487
rect 2225 15447 2283 15453
rect 5920 15428 5948 15524
rect 6270 15512 6276 15564
rect 6328 15552 6334 15564
rect 6733 15555 6791 15561
rect 6733 15552 6745 15555
rect 6328 15524 6745 15552
rect 6328 15512 6334 15524
rect 6733 15521 6745 15524
rect 6779 15552 6791 15555
rect 7561 15555 7619 15561
rect 6779 15524 7052 15552
rect 6779 15521 6791 15524
rect 6733 15515 6791 15521
rect 6917 15487 6975 15493
rect 6917 15453 6929 15487
rect 6963 15453 6975 15487
rect 6917 15447 6975 15453
rect 5902 15416 5908 15428
rect 5815 15388 5908 15416
rect 5902 15376 5908 15388
rect 5960 15416 5966 15428
rect 6932 15416 6960 15447
rect 5960 15388 6960 15416
rect 7024 15416 7052 15524
rect 7561 15521 7573 15555
rect 7607 15552 7619 15555
rect 7650 15552 7656 15564
rect 7607 15524 7656 15552
rect 7607 15521 7619 15524
rect 7561 15515 7619 15521
rect 7650 15512 7656 15524
rect 7708 15512 7714 15564
rect 8113 15555 8171 15561
rect 8113 15521 8125 15555
rect 8159 15552 8171 15555
rect 8941 15555 8999 15561
rect 8941 15552 8953 15555
rect 8159 15524 8953 15552
rect 8159 15521 8171 15524
rect 8113 15515 8171 15521
rect 8941 15521 8953 15524
rect 8987 15521 8999 15555
rect 8941 15515 8999 15521
rect 10045 15555 10103 15561
rect 10045 15521 10057 15555
rect 10091 15521 10103 15555
rect 10045 15515 10103 15521
rect 10873 15555 10931 15561
rect 10873 15521 10885 15555
rect 10919 15552 10931 15555
rect 10962 15552 10968 15564
rect 10919 15524 10968 15552
rect 10919 15521 10931 15524
rect 10873 15515 10931 15521
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15484 9275 15487
rect 9398 15484 9404 15496
rect 9263 15456 9404 15484
rect 9263 15453 9275 15456
rect 9217 15447 9275 15453
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 9674 15416 9680 15428
rect 7024 15388 9680 15416
rect 5960 15376 5966 15388
rect 9674 15376 9680 15388
rect 9732 15416 9738 15428
rect 10060 15416 10088 15515
rect 10962 15512 10968 15524
rect 11020 15512 11026 15564
rect 13262 15552 13268 15564
rect 13223 15524 13268 15552
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 14274 15552 14280 15564
rect 13464 15524 14280 15552
rect 10226 15484 10232 15496
rect 10187 15456 10232 15484
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 9732 15388 10088 15416
rect 13081 15419 13139 15425
rect 9732 15376 9738 15388
rect 13081 15385 13093 15419
rect 13127 15416 13139 15419
rect 13464 15416 13492 15524
rect 14274 15512 14280 15524
rect 14332 15552 14338 15564
rect 16592 15561 16620 15592
rect 17221 15589 17233 15592
rect 17267 15589 17279 15623
rect 17221 15583 17279 15589
rect 18776 15583 18788 15629
rect 18840 15620 18846 15632
rect 18840 15592 18876 15620
rect 18782 15580 18788 15583
rect 18840 15580 18846 15592
rect 15657 15555 15715 15561
rect 15657 15552 15669 15555
rect 14332 15524 15669 15552
rect 14332 15512 14338 15524
rect 15657 15521 15669 15524
rect 15703 15521 15715 15555
rect 15657 15515 15715 15521
rect 16117 15555 16175 15561
rect 16117 15521 16129 15555
rect 16163 15552 16175 15555
rect 16577 15555 16635 15561
rect 16577 15552 16589 15555
rect 16163 15524 16589 15552
rect 16163 15521 16175 15524
rect 16117 15515 16175 15521
rect 16577 15521 16589 15524
rect 16623 15521 16635 15555
rect 17589 15555 17647 15561
rect 17589 15552 17601 15555
rect 16577 15515 16635 15521
rect 16684 15524 17601 15552
rect 16684 15496 16712 15524
rect 17589 15521 17601 15524
rect 17635 15521 17647 15555
rect 17589 15515 17647 15521
rect 18138 15512 18144 15564
rect 18196 15552 18202 15564
rect 18509 15555 18567 15561
rect 18509 15552 18521 15555
rect 18196 15524 18521 15552
rect 18196 15512 18202 15524
rect 18509 15521 18521 15524
rect 18555 15552 18567 15555
rect 18598 15552 18604 15564
rect 18555 15524 18604 15552
rect 18555 15521 18567 15524
rect 18509 15515 18567 15521
rect 18598 15512 18604 15524
rect 18656 15512 18662 15564
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15484 13599 15487
rect 14366 15484 14372 15496
rect 13587 15456 14372 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 14642 15484 14648 15496
rect 14603 15456 14648 15484
rect 14642 15444 14648 15456
rect 14700 15444 14706 15496
rect 15838 15444 15844 15496
rect 15896 15484 15902 15496
rect 16666 15484 16672 15496
rect 15896 15456 16672 15484
rect 15896 15444 15902 15456
rect 16666 15444 16672 15456
rect 16724 15444 16730 15496
rect 16758 15444 16764 15496
rect 16816 15484 16822 15496
rect 16816 15456 16861 15484
rect 16816 15444 16822 15456
rect 13127 15388 13492 15416
rect 13127 15385 13139 15388
rect 13081 15379 13139 15385
rect 14090 15376 14096 15428
rect 14148 15416 14154 15428
rect 15378 15416 15384 15428
rect 14148 15388 15384 15416
rect 14148 15376 14154 15388
rect 15378 15376 15384 15388
rect 15436 15416 15442 15428
rect 15473 15419 15531 15425
rect 15473 15416 15485 15419
rect 15436 15388 15485 15416
rect 15436 15376 15442 15388
rect 15473 15385 15485 15388
rect 15519 15385 15531 15419
rect 15473 15379 15531 15385
rect 15562 15376 15568 15428
rect 15620 15416 15626 15428
rect 17957 15419 18015 15425
rect 17957 15416 17969 15419
rect 15620 15388 17969 15416
rect 15620 15376 15626 15388
rect 17957 15385 17969 15388
rect 18003 15416 18015 15419
rect 18506 15416 18512 15428
rect 18003 15388 18512 15416
rect 18003 15385 18015 15388
rect 17957 15379 18015 15385
rect 18506 15376 18512 15388
rect 18564 15376 18570 15428
rect 3326 15348 3332 15360
rect 3287 15320 3332 15348
rect 3326 15308 3332 15320
rect 3384 15308 3390 15360
rect 5442 15308 5448 15360
rect 5500 15348 5506 15360
rect 6089 15351 6147 15357
rect 6089 15348 6101 15351
rect 5500 15320 6101 15348
rect 5500 15308 5506 15320
rect 6089 15317 6101 15320
rect 6135 15317 6147 15351
rect 6089 15311 6147 15317
rect 12253 15351 12311 15357
rect 12253 15317 12265 15351
rect 12299 15348 12311 15351
rect 12434 15348 12440 15360
rect 12299 15320 12440 15348
rect 12299 15317 12311 15320
rect 12253 15311 12311 15317
rect 12434 15308 12440 15320
rect 12492 15308 12498 15360
rect 13446 15308 13452 15360
rect 13504 15348 13510 15360
rect 16117 15351 16175 15357
rect 16117 15348 16129 15351
rect 13504 15320 16129 15348
rect 13504 15308 13510 15320
rect 16117 15317 16129 15320
rect 16163 15317 16175 15351
rect 19886 15348 19892 15360
rect 19847 15320 19892 15348
rect 16117 15311 16175 15317
rect 19886 15308 19892 15320
rect 19944 15308 19950 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 1670 15144 1676 15156
rect 1631 15116 1676 15144
rect 1670 15104 1676 15116
rect 1728 15104 1734 15156
rect 2884 15116 3832 15144
rect 1946 14968 1952 15020
rect 2004 15008 2010 15020
rect 2884 15017 2912 15116
rect 3804 15076 3832 15116
rect 4246 15104 4252 15156
rect 4304 15144 4310 15156
rect 4525 15147 4583 15153
rect 4525 15144 4537 15147
rect 4304 15116 4537 15144
rect 4304 15104 4310 15116
rect 4525 15113 4537 15116
rect 4571 15113 4583 15147
rect 6270 15144 6276 15156
rect 6231 15116 6276 15144
rect 4525 15107 4583 15113
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 6638 15104 6644 15156
rect 6696 15144 6702 15156
rect 7193 15147 7251 15153
rect 7193 15144 7205 15147
rect 6696 15116 7205 15144
rect 6696 15104 6702 15116
rect 7193 15113 7205 15116
rect 7239 15113 7251 15147
rect 9398 15144 9404 15156
rect 9359 15116 9404 15144
rect 7193 15107 7251 15113
rect 9398 15104 9404 15116
rect 9456 15104 9462 15156
rect 10318 15104 10324 15156
rect 10376 15144 10382 15156
rect 11333 15147 11391 15153
rect 11333 15144 11345 15147
rect 10376 15116 11345 15144
rect 10376 15104 10382 15116
rect 11333 15113 11345 15116
rect 11379 15113 11391 15147
rect 12526 15144 12532 15156
rect 12487 15116 12532 15144
rect 11333 15107 11391 15113
rect 12526 15104 12532 15116
rect 12584 15104 12590 15156
rect 13906 15104 13912 15156
rect 13964 15144 13970 15156
rect 14001 15147 14059 15153
rect 14001 15144 14013 15147
rect 13964 15116 14013 15144
rect 13964 15104 13970 15116
rect 14001 15113 14013 15116
rect 14047 15113 14059 15147
rect 15470 15144 15476 15156
rect 15431 15116 15476 15144
rect 14001 15107 14059 15113
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 16850 15104 16856 15156
rect 16908 15144 16914 15156
rect 17313 15147 17371 15153
rect 17313 15144 17325 15147
rect 16908 15116 17325 15144
rect 16908 15104 16914 15116
rect 17313 15113 17325 15116
rect 17359 15113 17371 15147
rect 17313 15107 17371 15113
rect 3804 15048 4384 15076
rect 4356 15020 4384 15048
rect 4798 15036 4804 15088
rect 4856 15076 4862 15088
rect 6822 15076 6828 15088
rect 4856 15048 6828 15076
rect 4856 15036 4862 15048
rect 6822 15036 6828 15048
rect 6880 15036 6886 15088
rect 12066 15076 12072 15088
rect 12027 15048 12072 15076
rect 12066 15036 12072 15048
rect 12124 15036 12130 15088
rect 12544 15076 12572 15104
rect 15013 15079 15071 15085
rect 15013 15076 15025 15079
rect 12544 15048 15025 15076
rect 15013 15045 15025 15048
rect 15059 15076 15071 15079
rect 15654 15076 15660 15088
rect 15059 15048 15660 15076
rect 15059 15045 15071 15048
rect 15013 15039 15071 15045
rect 15654 15036 15660 15048
rect 15712 15036 15718 15088
rect 19061 15079 19119 15085
rect 19061 15076 19073 15079
rect 18524 15048 19073 15076
rect 2225 15011 2283 15017
rect 2225 15008 2237 15011
rect 2004 14980 2237 15008
rect 2004 14968 2010 14980
rect 2225 14977 2237 14980
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 14977 2927 15011
rect 2869 14971 2927 14977
rect 4338 14968 4344 15020
rect 4396 15008 4402 15020
rect 4816 15008 4844 15036
rect 4396 14980 4844 15008
rect 12084 15008 12112 15036
rect 13357 15011 13415 15017
rect 13357 15008 13369 15011
rect 12084 14980 13369 15008
rect 4396 14968 4402 14980
rect 13357 14977 13369 14980
rect 13403 14977 13415 15011
rect 13538 15008 13544 15020
rect 13499 14980 13544 15008
rect 13357 14971 13415 14977
rect 1489 14943 1547 14949
rect 1489 14909 1501 14943
rect 1535 14909 1547 14943
rect 1489 14903 1547 14909
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14940 2099 14943
rect 3136 14943 3194 14949
rect 2087 14912 3096 14940
rect 2087 14909 2099 14912
rect 2041 14903 2099 14909
rect 1504 14872 1532 14903
rect 2222 14872 2228 14884
rect 1504 14844 2228 14872
rect 2222 14832 2228 14844
rect 2280 14832 2286 14884
rect 3068 14872 3096 14912
rect 3136 14909 3148 14943
rect 3182 14940 3194 14943
rect 4154 14940 4160 14952
rect 3182 14912 4160 14940
rect 3182 14909 3194 14912
rect 3136 14903 3194 14909
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14940 8079 14943
rect 8662 14940 8668 14952
rect 8067 14912 8668 14940
rect 8067 14909 8079 14912
rect 8021 14903 8079 14909
rect 8662 14900 8668 14912
rect 8720 14940 8726 14952
rect 9677 14943 9735 14949
rect 9677 14940 9689 14943
rect 8720 14912 9689 14940
rect 8720 14900 8726 14912
rect 9677 14909 9689 14912
rect 9723 14909 9735 14943
rect 10226 14940 10232 14952
rect 9677 14903 9735 14909
rect 9784 14912 10232 14940
rect 5718 14872 5724 14884
rect 3068 14844 5724 14872
rect 5718 14832 5724 14844
rect 5776 14832 5782 14884
rect 8288 14875 8346 14881
rect 5828 14844 6316 14872
rect 3786 14764 3792 14816
rect 3844 14804 3850 14816
rect 4249 14807 4307 14813
rect 4249 14804 4261 14807
rect 3844 14776 4261 14804
rect 3844 14764 3850 14776
rect 4249 14773 4261 14776
rect 4295 14773 4307 14807
rect 4249 14767 4307 14773
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 5828 14804 5856 14844
rect 5500 14776 5856 14804
rect 6288 14804 6316 14844
rect 8288 14841 8300 14875
rect 8334 14872 8346 14875
rect 9784 14872 9812 14912
rect 10226 14900 10232 14912
rect 10284 14900 10290 14952
rect 10502 14900 10508 14952
rect 10560 14940 10566 14952
rect 13265 14943 13323 14949
rect 13265 14940 13277 14943
rect 10560 14912 13277 14940
rect 10560 14900 10566 14912
rect 13265 14909 13277 14912
rect 13311 14909 13323 14943
rect 13265 14903 13323 14909
rect 9950 14881 9956 14884
rect 9944 14872 9956 14881
rect 8334 14844 9812 14872
rect 9911 14844 9956 14872
rect 8334 14841 8346 14844
rect 8288 14835 8346 14841
rect 9944 14835 9956 14844
rect 9950 14832 9956 14835
rect 10008 14832 10014 14884
rect 12066 14872 12072 14884
rect 10060 14844 12072 14872
rect 10060 14804 10088 14844
rect 12066 14832 12072 14844
rect 12124 14832 12130 14884
rect 6288 14776 10088 14804
rect 5500 14764 5506 14776
rect 10226 14764 10232 14816
rect 10284 14804 10290 14816
rect 11057 14807 11115 14813
rect 11057 14804 11069 14807
rect 10284 14776 11069 14804
rect 10284 14764 10290 14776
rect 11057 14773 11069 14776
rect 11103 14773 11115 14807
rect 12894 14804 12900 14816
rect 12855 14776 12900 14804
rect 11057 14767 11115 14773
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 13280 14804 13308 14903
rect 13372 14872 13400 14971
rect 13538 14968 13544 14980
rect 13596 14968 13602 15020
rect 14461 15011 14519 15017
rect 14461 15008 14473 15011
rect 14200 14980 14473 15008
rect 14200 14952 14228 14980
rect 14461 14977 14473 14980
rect 14507 14977 14519 15011
rect 14642 15008 14648 15020
rect 14603 14980 14648 15008
rect 14461 14971 14519 14977
rect 14642 14968 14648 14980
rect 14700 14968 14706 15020
rect 17218 14968 17224 15020
rect 17276 15008 17282 15020
rect 18524 15017 18552 15048
rect 19061 15045 19073 15048
rect 19107 15045 19119 15079
rect 19061 15039 19119 15045
rect 18509 15011 18567 15017
rect 18509 15008 18521 15011
rect 17276 14980 18521 15008
rect 17276 14968 17282 14980
rect 18509 14977 18521 14980
rect 18555 14977 18567 15011
rect 18509 14971 18567 14977
rect 18693 15011 18751 15017
rect 18693 14977 18705 15011
rect 18739 15008 18751 15011
rect 19334 15008 19340 15020
rect 18739 14980 19340 15008
rect 18739 14977 18751 14980
rect 18693 14971 18751 14977
rect 19334 14968 19340 14980
rect 19392 15008 19398 15020
rect 19886 15008 19892 15020
rect 19392 14980 19892 15008
rect 19392 14968 19398 14980
rect 19886 14968 19892 14980
rect 19944 14968 19950 15020
rect 14182 14900 14188 14952
rect 14240 14900 14246 14952
rect 14366 14940 14372 14952
rect 14327 14912 14372 14940
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 15930 14940 15936 14952
rect 15891 14912 15936 14940
rect 15930 14900 15936 14912
rect 15988 14900 15994 14952
rect 16022 14900 16028 14952
rect 16080 14940 16086 14952
rect 16080 14912 18552 14940
rect 16080 14900 16086 14912
rect 15838 14872 15844 14884
rect 13372 14844 15844 14872
rect 15838 14832 15844 14844
rect 15896 14832 15902 14884
rect 16200 14875 16258 14881
rect 16200 14841 16212 14875
rect 16246 14872 16258 14875
rect 16666 14872 16672 14884
rect 16246 14844 16672 14872
rect 16246 14841 16258 14844
rect 16200 14835 16258 14841
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 18417 14875 18475 14881
rect 18417 14872 18429 14875
rect 17604 14844 18429 14872
rect 17218 14804 17224 14816
rect 13280 14776 17224 14804
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 17402 14764 17408 14816
rect 17460 14804 17466 14816
rect 17604 14813 17632 14844
rect 18417 14841 18429 14844
rect 18463 14841 18475 14875
rect 18417 14835 18475 14841
rect 17589 14807 17647 14813
rect 17589 14804 17601 14807
rect 17460 14776 17601 14804
rect 17460 14764 17466 14776
rect 17589 14773 17601 14776
rect 17635 14773 17647 14807
rect 18046 14804 18052 14816
rect 18007 14776 18052 14804
rect 17589 14767 17647 14773
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 18524 14804 18552 14912
rect 18598 14900 18604 14952
rect 18656 14940 18662 14952
rect 19981 14943 20039 14949
rect 19981 14940 19993 14943
rect 18656 14912 19993 14940
rect 18656 14900 18662 14912
rect 19981 14909 19993 14912
rect 20027 14909 20039 14943
rect 19981 14903 20039 14909
rect 20248 14943 20306 14949
rect 20248 14909 20260 14943
rect 20294 14940 20306 14943
rect 21358 14940 21364 14952
rect 20294 14912 21364 14940
rect 20294 14909 20306 14912
rect 20248 14903 20306 14909
rect 21358 14900 21364 14912
rect 21416 14900 21422 14952
rect 21361 14807 21419 14813
rect 21361 14804 21373 14807
rect 18524 14776 21373 14804
rect 21361 14773 21373 14776
rect 21407 14773 21419 14807
rect 21361 14767 21419 14773
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 2409 14603 2467 14609
rect 2409 14569 2421 14603
rect 2455 14600 2467 14603
rect 2961 14603 3019 14609
rect 2961 14600 2973 14603
rect 2455 14572 2973 14600
rect 2455 14569 2467 14572
rect 2409 14563 2467 14569
rect 2961 14569 2973 14572
rect 3007 14569 3019 14603
rect 3326 14600 3332 14612
rect 3287 14572 3332 14600
rect 2961 14563 3019 14569
rect 3326 14560 3332 14572
rect 3384 14560 3390 14612
rect 3421 14603 3479 14609
rect 3421 14569 3433 14603
rect 3467 14600 3479 14603
rect 4246 14600 4252 14612
rect 3467 14572 4252 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 5442 14600 5448 14612
rect 5403 14572 5448 14600
rect 5442 14560 5448 14572
rect 5500 14560 5506 14612
rect 5718 14600 5724 14612
rect 5679 14572 5724 14600
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 8941 14603 8999 14609
rect 8941 14600 8953 14603
rect 7708 14572 8953 14600
rect 7708 14560 7714 14572
rect 8941 14569 8953 14572
rect 8987 14569 8999 14603
rect 9674 14600 9680 14612
rect 9635 14572 9680 14600
rect 8941 14563 8999 14569
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 10502 14600 10508 14612
rect 10463 14572 10508 14600
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 13262 14600 13268 14612
rect 12176 14572 13268 14600
rect 5460 14532 5488 14560
rect 3528 14504 5488 14532
rect 6089 14535 6147 14541
rect 2317 14467 2375 14473
rect 2317 14433 2329 14467
rect 2363 14464 2375 14467
rect 2866 14464 2872 14476
rect 2363 14436 2872 14464
rect 2363 14433 2375 14436
rect 2317 14427 2375 14433
rect 2866 14424 2872 14436
rect 2924 14424 2930 14476
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 2501 14399 2559 14405
rect 2501 14396 2513 14399
rect 1719 14368 2513 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 2501 14365 2513 14368
rect 2547 14396 2559 14399
rect 3528 14396 3556 14504
rect 6089 14501 6101 14535
rect 6135 14532 6147 14535
rect 8481 14535 8539 14541
rect 8481 14532 8493 14535
rect 6135 14504 8493 14532
rect 6135 14501 6147 14504
rect 6089 14495 6147 14501
rect 8481 14501 8493 14504
rect 8527 14501 8539 14535
rect 10870 14532 10876 14544
rect 10831 14504 10876 14532
rect 8481 14495 8539 14501
rect 10870 14492 10876 14504
rect 10928 14492 10934 14544
rect 4321 14467 4379 14473
rect 4321 14464 4333 14467
rect 3804 14436 4333 14464
rect 3804 14408 3832 14436
rect 4321 14433 4333 14436
rect 4367 14433 4379 14467
rect 4321 14427 4379 14433
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14464 6239 14467
rect 6914 14464 6920 14476
rect 6227 14436 6920 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 7092 14467 7150 14473
rect 7092 14433 7104 14467
rect 7138 14464 7150 14467
rect 8386 14464 8392 14476
rect 7138 14436 8392 14464
rect 7138 14433 7150 14436
rect 7092 14427 7150 14433
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14433 9183 14467
rect 9125 14427 9183 14433
rect 2547 14368 3556 14396
rect 3605 14399 3663 14405
rect 2547 14365 2559 14368
rect 2501 14359 2559 14365
rect 3605 14365 3617 14399
rect 3651 14396 3663 14399
rect 3786 14396 3792 14408
rect 3651 14368 3792 14396
rect 3651 14365 3663 14368
rect 3605 14359 3663 14365
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 4062 14396 4068 14408
rect 4023 14368 4068 14396
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14365 6423 14399
rect 6822 14396 6828 14408
rect 6783 14368 6828 14396
rect 6365 14359 6423 14365
rect 6270 14328 6276 14340
rect 5368 14300 6276 14328
rect 1949 14263 2007 14269
rect 1949 14229 1961 14263
rect 1995 14260 2007 14263
rect 2774 14260 2780 14272
rect 1995 14232 2780 14260
rect 1995 14229 2007 14232
rect 1949 14223 2007 14229
rect 2774 14220 2780 14232
rect 2832 14220 2838 14272
rect 3326 14220 3332 14272
rect 3384 14260 3390 14272
rect 5368 14260 5396 14300
rect 6270 14288 6276 14300
rect 6328 14288 6334 14340
rect 3384 14232 5396 14260
rect 6380 14260 6408 14359
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 9140 14328 9168 14427
rect 12176 14337 12204 14572
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 13722 14600 13728 14612
rect 13596 14572 13728 14600
rect 13596 14560 13602 14572
rect 13722 14560 13728 14572
rect 13780 14600 13786 14612
rect 14277 14603 14335 14609
rect 14277 14600 14289 14603
rect 13780 14572 14289 14600
rect 13780 14560 13786 14572
rect 14277 14569 14289 14572
rect 14323 14569 14335 14603
rect 16666 14600 16672 14612
rect 16627 14572 16672 14600
rect 14277 14563 14335 14569
rect 16666 14560 16672 14572
rect 16724 14560 16730 14612
rect 12434 14492 12440 14544
rect 12492 14532 12498 14544
rect 13142 14535 13200 14541
rect 13142 14532 13154 14535
rect 12492 14504 13154 14532
rect 12492 14492 12498 14504
rect 13142 14501 13154 14504
rect 13188 14501 13200 14535
rect 17948 14535 18006 14541
rect 13142 14495 13200 14501
rect 15304 14504 15976 14532
rect 12897 14467 12955 14473
rect 12897 14433 12909 14467
rect 12943 14464 12955 14467
rect 13630 14464 13636 14476
rect 12943 14436 13636 14464
rect 12943 14433 12955 14436
rect 12897 14427 12955 14433
rect 13630 14424 13636 14436
rect 13688 14424 13694 14476
rect 15304 14473 15332 14504
rect 15948 14476 15976 14504
rect 17948 14501 17960 14535
rect 17994 14532 18006 14535
rect 19334 14532 19340 14544
rect 17994 14504 19340 14532
rect 17994 14501 18006 14504
rect 17948 14495 18006 14501
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 15556 14467 15614 14473
rect 15556 14433 15568 14467
rect 15602 14464 15614 14467
rect 15838 14464 15844 14476
rect 15602 14436 15844 14464
rect 15602 14433 15614 14436
rect 15556 14427 15614 14433
rect 15838 14424 15844 14436
rect 15896 14424 15902 14476
rect 15930 14424 15936 14476
rect 15988 14464 15994 14476
rect 17681 14467 17739 14473
rect 17681 14464 17693 14467
rect 15988 14436 17693 14464
rect 15988 14424 15994 14436
rect 17681 14433 17693 14436
rect 17727 14464 17739 14467
rect 18506 14464 18512 14476
rect 17727 14436 18512 14464
rect 17727 14433 17739 14436
rect 17681 14427 17739 14433
rect 18506 14424 18512 14436
rect 18564 14424 18570 14476
rect 16942 14396 16948 14408
rect 16903 14368 16948 14396
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 19334 14396 19340 14408
rect 19295 14368 19340 14396
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 12161 14331 12219 14337
rect 12161 14328 12173 14331
rect 9140 14300 12173 14328
rect 12161 14297 12173 14300
rect 12207 14297 12219 14331
rect 12161 14291 12219 14297
rect 7098 14260 7104 14272
rect 6380 14232 7104 14260
rect 3384 14220 3390 14232
rect 7098 14220 7104 14232
rect 7156 14260 7162 14272
rect 8018 14260 8024 14272
rect 7156 14232 8024 14260
rect 7156 14220 7162 14232
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 8202 14260 8208 14272
rect 8163 14232 8208 14260
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 14366 14260 14372 14272
rect 11940 14232 14372 14260
rect 11940 14220 11946 14232
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 14550 14260 14556 14272
rect 14511 14232 14556 14260
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 18690 14220 18696 14272
rect 18748 14260 18754 14272
rect 19061 14263 19119 14269
rect 19061 14260 19073 14263
rect 18748 14232 19073 14260
rect 18748 14220 18754 14232
rect 19061 14229 19073 14232
rect 19107 14229 19119 14263
rect 21358 14260 21364 14272
rect 21319 14232 21364 14260
rect 19061 14223 19119 14229
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 1486 14016 1492 14068
rect 1544 14056 1550 14068
rect 1673 14059 1731 14065
rect 1673 14056 1685 14059
rect 1544 14028 1685 14056
rect 1544 14016 1550 14028
rect 1673 14025 1685 14028
rect 1719 14025 1731 14059
rect 5902 14056 5908 14068
rect 1673 14019 1731 14025
rect 2056 14028 5672 14056
rect 5863 14028 5908 14056
rect 1486 13852 1492 13864
rect 1447 13824 1492 13852
rect 1486 13812 1492 13824
rect 1544 13812 1550 13864
rect 2056 13861 2084 14028
rect 5644 13988 5672 14028
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 7190 14056 7196 14068
rect 6012 14028 7196 14056
rect 6012 13988 6040 14028
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 8018 14016 8024 14068
rect 8076 14056 8082 14068
rect 8205 14059 8263 14065
rect 8205 14056 8217 14059
rect 8076 14028 8217 14056
rect 8076 14016 8082 14028
rect 8205 14025 8217 14028
rect 8251 14025 8263 14059
rect 8205 14019 8263 14025
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 12802 14056 12808 14068
rect 11379 14028 12808 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 14182 14056 14188 14068
rect 14143 14028 14188 14056
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 16209 14059 16267 14065
rect 16209 14025 16221 14059
rect 16255 14056 16267 14059
rect 16298 14056 16304 14068
rect 16255 14028 16304 14056
rect 16255 14025 16267 14028
rect 16209 14019 16267 14025
rect 16298 14016 16304 14028
rect 16356 14016 16362 14068
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 18049 14059 18107 14065
rect 18049 14056 18061 14059
rect 18012 14028 18061 14056
rect 18012 14016 18018 14028
rect 18049 14025 18061 14028
rect 18095 14025 18107 14059
rect 18049 14019 18107 14025
rect 5644 13960 6040 13988
rect 6270 13948 6276 14000
rect 6328 13988 6334 14000
rect 6365 13991 6423 13997
rect 6365 13988 6377 13991
rect 6328 13960 6377 13988
rect 6328 13948 6334 13960
rect 6365 13957 6377 13960
rect 6411 13957 6423 13991
rect 6365 13951 6423 13957
rect 2222 13920 2228 13932
rect 2183 13892 2228 13920
rect 2222 13880 2228 13892
rect 2280 13880 2286 13932
rect 2958 13920 2964 13932
rect 2919 13892 2964 13920
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13920 4215 13923
rect 4341 13923 4399 13929
rect 4341 13920 4353 13923
rect 4203 13892 4353 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 4341 13889 4353 13892
rect 4387 13889 4399 13923
rect 6380 13920 6408 13951
rect 9950 13948 9956 14000
rect 10008 13988 10014 14000
rect 10137 13991 10195 13997
rect 10137 13988 10149 13991
rect 10008 13960 10149 13988
rect 10008 13948 10014 13960
rect 10137 13957 10149 13960
rect 10183 13957 10195 13991
rect 10137 13951 10195 13957
rect 13446 13948 13452 14000
rect 13504 13988 13510 14000
rect 13817 13991 13875 13997
rect 13817 13988 13829 13991
rect 13504 13960 13829 13988
rect 13504 13948 13510 13960
rect 13817 13957 13829 13960
rect 13863 13957 13875 13991
rect 16022 13988 16028 14000
rect 13817 13951 13875 13957
rect 14844 13960 16028 13988
rect 11882 13920 11888 13932
rect 4341 13883 4399 13889
rect 4448 13892 4660 13920
rect 6380 13892 6960 13920
rect 11843 13892 11888 13920
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 3973 13855 4031 13861
rect 2832 13824 2877 13852
rect 2832 13812 2838 13824
rect 3973 13821 3985 13855
rect 4019 13852 4031 13855
rect 4448 13852 4476 13892
rect 4019 13824 4476 13852
rect 4525 13855 4583 13861
rect 4019 13821 4031 13824
rect 3973 13815 4031 13821
rect 4525 13821 4537 13855
rect 4571 13821 4583 13855
rect 4632 13852 4660 13892
rect 5718 13852 5724 13864
rect 4632 13824 5724 13852
rect 4525 13815 4583 13821
rect 3786 13744 3792 13796
rect 3844 13784 3850 13796
rect 4540 13784 4568 13815
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 6822 13852 6828 13864
rect 6783 13824 6828 13852
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 4792 13787 4850 13793
rect 4792 13784 4804 13787
rect 3844 13756 4568 13784
rect 4632 13756 4804 13784
rect 3844 13744 3850 13756
rect 3142 13676 3148 13728
rect 3200 13716 3206 13728
rect 3513 13719 3571 13725
rect 3513 13716 3525 13719
rect 3200 13688 3525 13716
rect 3200 13676 3206 13688
rect 3513 13685 3525 13688
rect 3559 13685 3571 13719
rect 3878 13716 3884 13728
rect 3839 13688 3884 13716
rect 3513 13679 3571 13685
rect 3878 13676 3884 13688
rect 3936 13676 3942 13728
rect 4341 13719 4399 13725
rect 4341 13685 4353 13719
rect 4387 13716 4399 13719
rect 4632 13716 4660 13756
rect 4792 13753 4804 13756
rect 4838 13784 4850 13787
rect 5442 13784 5448 13796
rect 4838 13756 5448 13784
rect 4838 13753 4850 13756
rect 4792 13747 4850 13753
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 6932 13784 6960 13892
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 14844 13929 14872 13960
rect 16022 13948 16028 13960
rect 16080 13948 16086 14000
rect 17313 13991 17371 13997
rect 17313 13988 17325 13991
rect 16500 13960 17325 13988
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13889 14887 13923
rect 15654 13920 15660 13932
rect 15615 13892 15660 13920
rect 14829 13883 14887 13889
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 15838 13920 15844 13932
rect 15751 13892 15844 13920
rect 15838 13880 15844 13892
rect 15896 13920 15902 13932
rect 16390 13920 16396 13932
rect 15896 13892 16396 13920
rect 15896 13880 15902 13892
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 7092 13855 7150 13861
rect 7092 13821 7104 13855
rect 7138 13852 7150 13855
rect 8202 13852 8208 13864
rect 7138 13824 8208 13852
rect 7138 13821 7150 13824
rect 7092 13815 7150 13821
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8754 13852 8760 13864
rect 8715 13824 8760 13852
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 11793 13855 11851 13861
rect 11793 13821 11805 13855
rect 11839 13852 11851 13855
rect 12342 13852 12348 13864
rect 11839 13824 12348 13852
rect 11839 13821 11851 13824
rect 11793 13815 11851 13821
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 12434 13812 12440 13864
rect 12492 13852 12498 13864
rect 12704 13855 12762 13861
rect 12492 13824 12537 13852
rect 12492 13812 12498 13824
rect 12704 13821 12716 13855
rect 12750 13852 12762 13855
rect 13722 13852 13728 13864
rect 12750 13824 13728 13852
rect 12750 13821 12762 13824
rect 12704 13815 12762 13821
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 14645 13855 14703 13861
rect 14645 13852 14657 13855
rect 14424 13824 14657 13852
rect 14424 13812 14430 13824
rect 14645 13821 14657 13824
rect 14691 13852 14703 13855
rect 16500 13852 16528 13960
rect 17313 13957 17325 13960
rect 17359 13988 17371 13991
rect 19242 13988 19248 14000
rect 17359 13960 19248 13988
rect 17359 13957 17371 13960
rect 17313 13951 17371 13957
rect 19242 13948 19248 13960
rect 19300 13948 19306 14000
rect 16666 13880 16672 13932
rect 16724 13920 16730 13932
rect 16761 13923 16819 13929
rect 16761 13920 16773 13923
rect 16724 13892 16773 13920
rect 16724 13880 16730 13892
rect 16761 13889 16773 13892
rect 16807 13889 16819 13923
rect 16761 13883 16819 13889
rect 18046 13880 18052 13932
rect 18104 13920 18110 13932
rect 18509 13923 18567 13929
rect 18509 13920 18521 13923
rect 18104 13892 18521 13920
rect 18104 13880 18110 13892
rect 18509 13889 18521 13892
rect 18555 13889 18567 13923
rect 18690 13920 18696 13932
rect 18651 13892 18696 13920
rect 18509 13883 18567 13889
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 14691 13824 16528 13852
rect 16577 13855 16635 13861
rect 14691 13821 14703 13824
rect 14645 13815 14703 13821
rect 16577 13821 16589 13855
rect 16623 13852 16635 13855
rect 16942 13852 16948 13864
rect 16623 13824 16948 13852
rect 16623 13821 16635 13824
rect 16577 13815 16635 13821
rect 16942 13812 16948 13824
rect 17000 13812 17006 13864
rect 7374 13784 7380 13796
rect 6932 13756 7380 13784
rect 7374 13744 7380 13756
rect 7432 13744 7438 13796
rect 9024 13787 9082 13793
rect 9024 13753 9036 13787
rect 9070 13784 9082 13787
rect 9582 13784 9588 13796
rect 9070 13756 9588 13784
rect 9070 13753 9082 13756
rect 9024 13747 9082 13753
rect 9582 13744 9588 13756
rect 9640 13744 9646 13796
rect 16669 13787 16727 13793
rect 16669 13784 16681 13787
rect 15212 13756 16681 13784
rect 4387 13688 4660 13716
rect 4387 13685 4399 13688
rect 4341 13679 4399 13685
rect 4706 13676 4712 13728
rect 4764 13716 4770 13728
rect 10410 13716 10416 13728
rect 4764 13688 10416 13716
rect 4764 13676 4770 13688
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 11698 13716 11704 13728
rect 11659 13688 11704 13716
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 14550 13716 14556 13728
rect 14511 13688 14556 13716
rect 14550 13676 14556 13688
rect 14608 13676 14614 13728
rect 15212 13725 15240 13756
rect 16669 13753 16681 13756
rect 16715 13753 16727 13787
rect 16669 13747 16727 13753
rect 18417 13787 18475 13793
rect 18417 13753 18429 13787
rect 18463 13784 18475 13787
rect 19334 13784 19340 13796
rect 18463 13756 19340 13784
rect 18463 13753 18475 13756
rect 18417 13747 18475 13753
rect 19334 13744 19340 13756
rect 19392 13744 19398 13796
rect 15197 13719 15255 13725
rect 15197 13685 15209 13719
rect 15243 13685 15255 13719
rect 15197 13679 15255 13685
rect 15286 13676 15292 13728
rect 15344 13716 15350 13728
rect 15565 13719 15623 13725
rect 15565 13716 15577 13719
rect 15344 13688 15577 13716
rect 15344 13676 15350 13688
rect 15565 13685 15577 13688
rect 15611 13685 15623 13719
rect 15565 13679 15623 13685
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 2961 13515 3019 13521
rect 2961 13512 2973 13515
rect 2924 13484 2973 13512
rect 2924 13472 2930 13484
rect 2961 13481 2973 13484
rect 3007 13481 3019 13515
rect 2961 13475 3019 13481
rect 3513 13515 3571 13521
rect 3513 13481 3525 13515
rect 3559 13512 3571 13515
rect 3878 13512 3884 13524
rect 3559 13484 3884 13512
rect 3559 13481 3571 13484
rect 3513 13475 3571 13481
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 5442 13512 5448 13524
rect 5403 13484 5448 13512
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7009 13515 7067 13521
rect 7009 13512 7021 13515
rect 6972 13484 7021 13512
rect 6972 13472 6978 13484
rect 7009 13481 7021 13484
rect 7055 13481 7067 13515
rect 7009 13475 7067 13481
rect 7190 13472 7196 13524
rect 7248 13512 7254 13524
rect 8573 13515 8631 13521
rect 8573 13512 8585 13515
rect 7248 13484 8585 13512
rect 7248 13472 7254 13484
rect 8573 13481 8585 13484
rect 8619 13481 8631 13515
rect 8573 13475 8631 13481
rect 9033 13515 9091 13521
rect 9033 13481 9045 13515
rect 9079 13512 9091 13515
rect 9677 13515 9735 13521
rect 9677 13512 9689 13515
rect 9079 13484 9689 13512
rect 9079 13481 9091 13484
rect 9033 13475 9091 13481
rect 9677 13481 9689 13484
rect 9723 13481 9735 13515
rect 9677 13475 9735 13481
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 10778 13512 10784 13524
rect 10183 13484 10784 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 12897 13515 12955 13521
rect 12897 13512 12909 13515
rect 11940 13484 12909 13512
rect 11940 13472 11946 13484
rect 12897 13481 12909 13484
rect 12943 13512 12955 13515
rect 13078 13512 13084 13524
rect 12943 13484 13084 13512
rect 12943 13481 12955 13484
rect 12897 13475 12955 13481
rect 13078 13472 13084 13484
rect 13136 13472 13142 13524
rect 13541 13515 13599 13521
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 14458 13512 14464 13524
rect 13587 13484 14464 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 1486 13404 1492 13456
rect 1544 13444 1550 13456
rect 2317 13447 2375 13453
rect 2317 13444 2329 13447
rect 1544 13416 2329 13444
rect 1544 13404 1550 13416
rect 2317 13413 2329 13416
rect 2363 13413 2375 13447
rect 2317 13407 2375 13413
rect 4332 13447 4390 13453
rect 4332 13413 4344 13447
rect 4378 13444 4390 13447
rect 5810 13444 5816 13456
rect 4378 13416 5816 13444
rect 4378 13413 4390 13416
rect 4332 13407 4390 13413
rect 5810 13404 5816 13416
rect 5868 13444 5874 13456
rect 7469 13447 7527 13453
rect 7469 13444 7481 13447
rect 5868 13416 6316 13444
rect 5868 13404 5874 13416
rect 2041 13379 2099 13385
rect 2041 13345 2053 13379
rect 2087 13376 2099 13379
rect 3142 13376 3148 13388
rect 2087 13348 3148 13376
rect 2087 13345 2099 13348
rect 2041 13339 2099 13345
rect 3142 13336 3148 13348
rect 3200 13336 3206 13388
rect 5902 13336 5908 13388
rect 5960 13376 5966 13388
rect 6089 13379 6147 13385
rect 6089 13376 6101 13379
rect 5960 13348 6101 13376
rect 5960 13336 5966 13348
rect 6089 13345 6101 13348
rect 6135 13345 6147 13379
rect 6089 13339 6147 13345
rect 3786 13268 3792 13320
rect 3844 13308 3850 13320
rect 6288 13317 6316 13416
rect 6932 13416 7481 13444
rect 6932 13388 6960 13416
rect 7469 13413 7481 13416
rect 7515 13444 7527 13447
rect 7558 13444 7564 13456
rect 7515 13416 7564 13444
rect 7515 13413 7527 13416
rect 7469 13407 7527 13413
rect 7558 13404 7564 13416
rect 7616 13404 7622 13456
rect 11241 13447 11299 13453
rect 11241 13413 11253 13447
rect 11287 13444 11299 13447
rect 13556 13444 13584 13475
rect 14458 13472 14464 13484
rect 14516 13512 14522 13524
rect 15749 13515 15807 13521
rect 15749 13512 15761 13515
rect 14516 13484 15761 13512
rect 14516 13472 14522 13484
rect 15749 13481 15761 13484
rect 15795 13481 15807 13515
rect 15749 13475 15807 13481
rect 11287 13416 13584 13444
rect 18040 13447 18098 13453
rect 11287 13413 11299 13416
rect 11241 13407 11299 13413
rect 18040 13413 18052 13447
rect 18086 13444 18098 13447
rect 18690 13444 18696 13456
rect 18086 13416 18696 13444
rect 18086 13413 18098 13416
rect 18040 13407 18098 13413
rect 18690 13404 18696 13416
rect 18748 13404 18754 13456
rect 6914 13336 6920 13388
rect 6972 13336 6978 13388
rect 7374 13376 7380 13388
rect 7335 13348 7380 13376
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13376 8999 13379
rect 9490 13376 9496 13388
rect 8987 13348 9496 13376
rect 8987 13345 8999 13348
rect 8941 13339 8999 13345
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 10042 13376 10048 13388
rect 10003 13348 10048 13376
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 11784 13379 11842 13385
rect 11784 13345 11796 13379
rect 11830 13376 11842 13379
rect 13446 13376 13452 13388
rect 11830 13348 13452 13376
rect 11830 13345 11842 13348
rect 11784 13339 11842 13345
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 14476 13348 15669 13376
rect 4065 13311 4123 13317
rect 4065 13308 4077 13311
rect 3844 13280 4077 13308
rect 3844 13268 3850 13280
rect 4065 13277 4077 13280
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 6181 13311 6239 13317
rect 6181 13277 6193 13311
rect 6227 13277 6239 13311
rect 6181 13271 6239 13277
rect 6273 13311 6331 13317
rect 6273 13277 6285 13311
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13308 7711 13311
rect 8202 13308 8208 13320
rect 7699 13280 8208 13308
rect 7699 13277 7711 13280
rect 7653 13271 7711 13277
rect 6196 13240 6224 13271
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 9950 13308 9956 13320
rect 9263 13280 9956 13308
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 9950 13268 9956 13280
rect 10008 13268 10014 13320
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 7282 13240 7288 13252
rect 6196 13212 7288 13240
rect 7282 13200 7288 13212
rect 7340 13240 7346 13252
rect 8021 13243 8079 13249
rect 8021 13240 8033 13243
rect 7340 13212 8033 13240
rect 7340 13200 7346 13212
rect 8021 13209 8033 13212
rect 8067 13209 8079 13243
rect 8021 13203 8079 13209
rect 9306 13200 9312 13252
rect 9364 13240 9370 13252
rect 9582 13240 9588 13252
rect 9364 13212 9588 13240
rect 9364 13200 9370 13212
rect 9582 13200 9588 13212
rect 9640 13240 9646 13252
rect 10244 13240 10272 13271
rect 9640 13212 10272 13240
rect 9640 13200 9646 13212
rect 3970 13132 3976 13184
rect 4028 13172 4034 13184
rect 10594 13172 10600 13184
rect 4028 13144 10600 13172
rect 4028 13132 4034 13144
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 11532 13172 11560 13271
rect 12986 13268 12992 13320
rect 13044 13308 13050 13320
rect 13538 13308 13544 13320
rect 13044 13280 13544 13308
rect 13044 13268 13050 13280
rect 13538 13268 13544 13280
rect 13596 13308 13602 13320
rect 13633 13311 13691 13317
rect 13633 13308 13645 13311
rect 13596 13280 13645 13308
rect 13596 13268 13602 13280
rect 13633 13277 13645 13280
rect 13679 13277 13691 13311
rect 13633 13271 13691 13277
rect 13722 13268 13728 13320
rect 13780 13308 13786 13320
rect 13780 13280 13825 13308
rect 13780 13268 13786 13280
rect 14090 13200 14096 13252
rect 14148 13240 14154 13252
rect 14476 13249 14504 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 15838 13268 15844 13320
rect 15896 13308 15902 13320
rect 16301 13311 16359 13317
rect 15896 13280 15941 13308
rect 15896 13268 15902 13280
rect 16301 13277 16313 13311
rect 16347 13308 16359 13311
rect 17034 13308 17040 13320
rect 16347 13280 17040 13308
rect 16347 13277 16359 13280
rect 16301 13271 16359 13277
rect 17034 13268 17040 13280
rect 17092 13268 17098 13320
rect 17770 13308 17776 13320
rect 17731 13280 17776 13308
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 14461 13243 14519 13249
rect 14461 13240 14473 13243
rect 14148 13212 14473 13240
rect 14148 13200 14154 13212
rect 14461 13209 14473 13212
rect 14507 13209 14519 13243
rect 14461 13203 14519 13209
rect 14918 13200 14924 13252
rect 14976 13240 14982 13252
rect 17405 13243 17463 13249
rect 17405 13240 17417 13243
rect 14976 13212 17417 13240
rect 14976 13200 14982 13212
rect 17405 13209 17417 13212
rect 17451 13240 17463 13243
rect 17678 13240 17684 13252
rect 17451 13212 17684 13240
rect 17451 13209 17463 13212
rect 17405 13203 17463 13209
rect 17678 13200 17684 13212
rect 17736 13200 17742 13252
rect 12434 13172 12440 13184
rect 11532 13144 12440 13172
rect 12434 13132 12440 13144
rect 12492 13172 12498 13184
rect 12710 13172 12716 13184
rect 12492 13144 12716 13172
rect 12492 13132 12498 13144
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 12986 13132 12992 13184
rect 13044 13172 13050 13184
rect 13173 13175 13231 13181
rect 13173 13172 13185 13175
rect 13044 13144 13185 13172
rect 13044 13132 13050 13144
rect 13173 13141 13185 13144
rect 13219 13141 13231 13175
rect 13173 13135 13231 13141
rect 13998 13132 14004 13184
rect 14056 13172 14062 13184
rect 14829 13175 14887 13181
rect 14829 13172 14841 13175
rect 14056 13144 14841 13172
rect 14056 13132 14062 13144
rect 14829 13141 14841 13144
rect 14875 13172 14887 13175
rect 15102 13172 15108 13184
rect 14875 13144 15108 13172
rect 14875 13141 14887 13144
rect 14829 13135 14887 13141
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 15289 13175 15347 13181
rect 15289 13141 15301 13175
rect 15335 13172 15347 13175
rect 17126 13172 17132 13184
rect 15335 13144 17132 13172
rect 15335 13141 15347 13144
rect 15289 13135 15347 13141
rect 17126 13132 17132 13144
rect 17184 13132 17190 13184
rect 19150 13172 19156 13184
rect 19111 13144 19156 13172
rect 19150 13132 19156 13144
rect 19208 13132 19214 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1946 12968 1952 12980
rect 1907 12940 1952 12968
rect 1946 12928 1952 12940
rect 2004 12928 2010 12980
rect 2501 12971 2559 12977
rect 2501 12937 2513 12971
rect 2547 12968 2559 12971
rect 3050 12968 3056 12980
rect 2547 12940 3056 12968
rect 2547 12937 2559 12940
rect 2501 12931 2559 12937
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 3602 12968 3608 12980
rect 3563 12940 3608 12968
rect 3602 12928 3608 12940
rect 3660 12928 3666 12980
rect 4154 12928 4160 12980
rect 4212 12968 4218 12980
rect 5810 12968 5816 12980
rect 4212 12940 5396 12968
rect 5771 12940 5816 12968
rect 4212 12928 4218 12940
rect 5368 12900 5396 12940
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 8481 12971 8539 12977
rect 8481 12968 8493 12971
rect 6196 12940 8493 12968
rect 6196 12900 6224 12940
rect 8481 12937 8493 12940
rect 8527 12937 8539 12971
rect 8481 12931 8539 12937
rect 11333 12971 11391 12977
rect 11333 12937 11345 12971
rect 11379 12968 11391 12971
rect 11698 12968 11704 12980
rect 11379 12940 11704 12968
rect 11379 12937 11391 12940
rect 11333 12931 11391 12937
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 12342 12928 12348 12980
rect 12400 12968 12406 12980
rect 12529 12971 12587 12977
rect 12529 12968 12541 12971
rect 12400 12940 12541 12968
rect 12400 12928 12406 12940
rect 12529 12937 12541 12940
rect 12575 12937 12587 12971
rect 13538 12968 13544 12980
rect 13499 12940 13544 12968
rect 12529 12931 12587 12937
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 14458 12928 14464 12980
rect 14516 12968 14522 12980
rect 14645 12971 14703 12977
rect 14645 12968 14657 12971
rect 14516 12940 14657 12968
rect 14516 12928 14522 12940
rect 14645 12937 14657 12940
rect 14691 12937 14703 12971
rect 16390 12968 16396 12980
rect 16351 12940 16396 12968
rect 14645 12931 14703 12937
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 16574 12928 16580 12980
rect 16632 12968 16638 12980
rect 16669 12971 16727 12977
rect 16669 12968 16681 12971
rect 16632 12940 16681 12968
rect 16632 12928 16638 12940
rect 16669 12937 16681 12940
rect 16715 12937 16727 12971
rect 16669 12931 16727 12937
rect 18874 12928 18880 12980
rect 18932 12968 18938 12980
rect 19061 12971 19119 12977
rect 19061 12968 19073 12971
rect 18932 12940 19073 12968
rect 18932 12928 18938 12940
rect 19061 12937 19073 12940
rect 19107 12937 19119 12971
rect 19061 12931 19119 12937
rect 5368 12872 6224 12900
rect 11992 12872 13216 12900
rect 9030 12832 9036 12844
rect 8991 12804 9036 12832
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 9490 12832 9496 12844
rect 9451 12804 9496 12832
rect 9490 12792 9496 12804
rect 9548 12792 9554 12844
rect 11992 12841 12020 12872
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12801 12035 12835
rect 12986 12832 12992 12844
rect 12947 12804 12992 12832
rect 11977 12795 12035 12801
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13188 12841 13216 12872
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12832 13231 12835
rect 13446 12832 13452 12844
rect 13219 12804 13452 12832
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 13446 12792 13452 12804
rect 13504 12792 13510 12844
rect 17126 12832 17132 12844
rect 17087 12804 17132 12832
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12801 17279 12835
rect 17221 12795 17279 12801
rect 1765 12767 1823 12773
rect 1765 12733 1777 12767
rect 1811 12764 1823 12767
rect 2038 12764 2044 12776
rect 1811 12736 2044 12764
rect 1811 12733 1823 12736
rect 1765 12727 1823 12733
rect 2038 12724 2044 12736
rect 2096 12724 2102 12776
rect 2317 12767 2375 12773
rect 2317 12733 2329 12767
rect 2363 12764 2375 12767
rect 2774 12764 2780 12776
rect 2363 12736 2780 12764
rect 2363 12733 2375 12736
rect 2317 12727 2375 12733
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 2869 12767 2927 12773
rect 2869 12733 2881 12767
rect 2915 12764 2927 12767
rect 3142 12764 3148 12776
rect 2915 12736 3148 12764
rect 2915 12733 2927 12736
rect 2869 12727 2927 12733
rect 3142 12724 3148 12736
rect 3200 12724 3206 12776
rect 3418 12764 3424 12776
rect 3379 12736 3424 12764
rect 3418 12724 3424 12736
rect 3476 12724 3482 12776
rect 3786 12724 3792 12776
rect 3844 12764 3850 12776
rect 7098 12773 7104 12776
rect 4433 12767 4491 12773
rect 4433 12764 4445 12767
rect 3844 12736 4445 12764
rect 3844 12724 3850 12736
rect 4433 12733 4445 12736
rect 4479 12764 4491 12767
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 4479 12736 6837 12764
rect 4479 12733 4491 12736
rect 4433 12727 4491 12733
rect 6825 12733 6837 12736
rect 6871 12733 6883 12767
rect 7092 12764 7104 12773
rect 7059 12736 7104 12764
rect 6825 12727 6883 12733
rect 7092 12727 7104 12736
rect 7098 12724 7104 12727
rect 7156 12724 7162 12776
rect 9953 12767 10011 12773
rect 9953 12764 9965 12767
rect 7668 12736 9965 12764
rect 4700 12699 4758 12705
rect 4700 12665 4712 12699
rect 4746 12696 4758 12699
rect 4798 12696 4804 12708
rect 4746 12668 4804 12696
rect 4746 12665 4758 12668
rect 4700 12659 4758 12665
rect 4798 12656 4804 12668
rect 4856 12656 4862 12708
rect 5902 12656 5908 12708
rect 5960 12696 5966 12708
rect 7668 12696 7696 12736
rect 9953 12733 9965 12736
rect 9999 12764 10011 12767
rect 10042 12764 10048 12776
rect 9999 12736 10048 12764
rect 9999 12733 10011 12736
rect 9953 12727 10011 12733
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12764 10747 12767
rect 11882 12764 11888 12776
rect 10735 12736 11888 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 12894 12764 12900 12776
rect 12855 12736 12900 12764
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 14274 12724 14280 12776
rect 14332 12764 14338 12776
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 14332 12736 14381 12764
rect 14332 12724 14338 12736
rect 14369 12733 14381 12736
rect 14415 12733 14427 12767
rect 14369 12727 14427 12733
rect 14642 12724 14648 12776
rect 14700 12764 14706 12776
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 14700 12736 15025 12764
rect 14700 12724 14706 12736
rect 15013 12733 15025 12736
rect 15059 12733 15071 12767
rect 17034 12764 17040 12776
rect 16995 12736 17040 12764
rect 15013 12727 15071 12733
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 17236 12764 17264 12795
rect 17678 12792 17684 12844
rect 17736 12832 17742 12844
rect 18509 12835 18567 12841
rect 18509 12832 18521 12835
rect 17736 12804 18521 12832
rect 17736 12792 17742 12804
rect 18509 12801 18521 12804
rect 18555 12801 18567 12835
rect 18690 12832 18696 12844
rect 18603 12804 18696 12832
rect 18509 12795 18567 12801
rect 18690 12792 18696 12804
rect 18748 12832 18754 12844
rect 19150 12832 19156 12844
rect 18748 12804 19156 12832
rect 18748 12792 18754 12804
rect 19150 12792 19156 12804
rect 19208 12792 19214 12844
rect 19613 12835 19671 12841
rect 19613 12801 19625 12835
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 17144 12736 17264 12764
rect 5960 12668 7696 12696
rect 5960 12656 5966 12668
rect 7742 12656 7748 12708
rect 7800 12696 7806 12708
rect 8849 12699 8907 12705
rect 8849 12696 8861 12699
rect 7800 12668 8861 12696
rect 7800 12656 7806 12668
rect 8849 12665 8861 12668
rect 8895 12665 8907 12699
rect 8849 12659 8907 12665
rect 11701 12699 11759 12705
rect 11701 12665 11713 12699
rect 11747 12696 11759 12699
rect 12802 12696 12808 12708
rect 11747 12668 12808 12696
rect 11747 12665 11759 12668
rect 11701 12659 11759 12665
rect 12802 12656 12808 12668
rect 12860 12656 12866 12708
rect 14918 12696 14924 12708
rect 14108 12668 14924 12696
rect 3053 12631 3111 12637
rect 3053 12597 3065 12631
rect 3099 12628 3111 12631
rect 3234 12628 3240 12640
rect 3099 12600 3240 12628
rect 3099 12597 3111 12600
rect 3053 12591 3111 12597
rect 3234 12588 3240 12600
rect 3292 12588 3298 12640
rect 6457 12631 6515 12637
rect 6457 12597 6469 12631
rect 6503 12628 6515 12631
rect 6914 12628 6920 12640
rect 6503 12600 6920 12628
rect 6503 12597 6515 12600
rect 6457 12591 6515 12597
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 7190 12588 7196 12640
rect 7248 12628 7254 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 7248 12600 8217 12628
rect 7248 12588 7254 12600
rect 8205 12597 8217 12600
rect 8251 12597 8263 12631
rect 8205 12591 8263 12597
rect 8938 12588 8944 12640
rect 8996 12628 9002 12640
rect 11054 12628 11060 12640
rect 8996 12600 9041 12628
rect 10967 12600 11060 12628
rect 8996 12588 9002 12600
rect 11054 12588 11060 12600
rect 11112 12628 11118 12640
rect 11793 12631 11851 12637
rect 11793 12628 11805 12631
rect 11112 12600 11805 12628
rect 11112 12588 11118 12600
rect 11793 12597 11805 12600
rect 11839 12597 11851 12631
rect 11793 12591 11851 12597
rect 11882 12588 11888 12640
rect 11940 12628 11946 12640
rect 12250 12628 12256 12640
rect 11940 12600 12256 12628
rect 11940 12588 11946 12600
rect 12250 12588 12256 12600
rect 12308 12628 12314 12640
rect 14108 12628 14136 12668
rect 14918 12656 14924 12668
rect 14976 12656 14982 12708
rect 15280 12699 15338 12705
rect 15280 12665 15292 12699
rect 15326 12696 15338 12699
rect 16758 12696 16764 12708
rect 15326 12668 16764 12696
rect 15326 12665 15338 12668
rect 15280 12659 15338 12665
rect 16758 12656 16764 12668
rect 16816 12696 16822 12708
rect 17144 12696 17172 12736
rect 18782 12724 18788 12776
rect 18840 12764 18846 12776
rect 19628 12764 19656 12795
rect 18840 12736 19656 12764
rect 18840 12724 18846 12736
rect 19521 12699 19579 12705
rect 19521 12696 19533 12699
rect 16816 12668 17172 12696
rect 18064 12668 19533 12696
rect 16816 12656 16822 12668
rect 12308 12600 14136 12628
rect 14185 12631 14243 12637
rect 12308 12588 12314 12600
rect 14185 12597 14197 12631
rect 14231 12628 14243 12631
rect 14274 12628 14280 12640
rect 14231 12600 14280 12628
rect 14231 12597 14243 12600
rect 14185 12591 14243 12597
rect 14274 12588 14280 12600
rect 14332 12588 14338 12640
rect 18064 12637 18092 12668
rect 19521 12665 19533 12668
rect 19567 12665 19579 12699
rect 19521 12659 19579 12665
rect 18049 12631 18107 12637
rect 18049 12597 18061 12631
rect 18095 12597 18107 12631
rect 18049 12591 18107 12597
rect 18417 12631 18475 12637
rect 18417 12597 18429 12631
rect 18463 12628 18475 12631
rect 19242 12628 19248 12640
rect 18463 12600 19248 12628
rect 18463 12597 18475 12600
rect 18417 12591 18475 12597
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 19426 12628 19432 12640
rect 19387 12600 19432 12628
rect 19426 12588 19432 12600
rect 19484 12588 19490 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 3510 12384 3516 12436
rect 3568 12424 3574 12436
rect 9306 12424 9312 12436
rect 3568 12396 9168 12424
rect 9267 12396 9312 12424
rect 3568 12384 3574 12396
rect 3142 12356 3148 12368
rect 3103 12328 3148 12356
rect 3142 12316 3148 12328
rect 3200 12316 3206 12368
rect 7650 12356 7656 12368
rect 6288 12328 7656 12356
rect 2130 12288 2136 12300
rect 2091 12260 2136 12288
rect 2130 12248 2136 12260
rect 2188 12248 2194 12300
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12288 2927 12291
rect 4154 12288 4160 12300
rect 2915 12260 4160 12288
rect 2915 12257 2927 12260
rect 2869 12251 2927 12257
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 4332 12291 4390 12297
rect 4332 12257 4344 12291
rect 4378 12288 4390 12291
rect 5442 12288 5448 12300
rect 4378 12260 5448 12288
rect 4378 12257 4390 12260
rect 4332 12251 4390 12257
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 6288 12297 6316 12328
rect 7650 12316 7656 12328
rect 7708 12316 7714 12368
rect 8196 12359 8254 12365
rect 8196 12325 8208 12359
rect 8242 12356 8254 12359
rect 8478 12356 8484 12368
rect 8242 12328 8484 12356
rect 8242 12325 8254 12328
rect 8196 12319 8254 12325
rect 8478 12316 8484 12328
rect 8536 12356 8542 12368
rect 9030 12356 9036 12368
rect 8536 12328 9036 12356
rect 8536 12316 8542 12328
rect 9030 12316 9036 12328
rect 9088 12316 9094 12368
rect 9140 12356 9168 12396
rect 9306 12384 9312 12396
rect 9364 12384 9370 12436
rect 11609 12427 11667 12433
rect 11609 12393 11621 12427
rect 11655 12424 11667 12427
rect 11882 12424 11888 12436
rect 11655 12396 11888 12424
rect 11655 12393 11667 12396
rect 11609 12387 11667 12393
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 14093 12427 14151 12433
rect 14093 12393 14105 12427
rect 14139 12424 14151 12427
rect 14734 12424 14740 12436
rect 14139 12396 14740 12424
rect 14139 12393 14151 12396
rect 14093 12387 14151 12393
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 16669 12427 16727 12433
rect 16669 12393 16681 12427
rect 16715 12424 16727 12427
rect 16758 12424 16764 12436
rect 16715 12396 16764 12424
rect 16715 12393 16727 12396
rect 16669 12387 16727 12393
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 19242 12384 19248 12436
rect 19300 12424 19306 12436
rect 19337 12427 19395 12433
rect 19337 12424 19349 12427
rect 19300 12396 19349 12424
rect 19300 12384 19306 12396
rect 19337 12393 19349 12396
rect 19383 12393 19395 12427
rect 19337 12387 19395 12393
rect 9677 12359 9735 12365
rect 9677 12356 9689 12359
rect 9140 12328 9689 12356
rect 9677 12325 9689 12328
rect 9723 12356 9735 12359
rect 10505 12359 10563 12365
rect 10505 12356 10517 12359
rect 9723 12328 10517 12356
rect 9723 12325 9735 12328
rect 9677 12319 9735 12325
rect 10505 12325 10517 12328
rect 10551 12325 10563 12359
rect 10505 12319 10563 12325
rect 11146 12316 11152 12368
rect 11204 12356 11210 12368
rect 11790 12356 11796 12368
rect 11204 12328 11796 12356
rect 11204 12316 11210 12328
rect 11790 12316 11796 12328
rect 11848 12316 11854 12368
rect 12428 12359 12486 12365
rect 12428 12325 12440 12359
rect 12474 12356 12486 12359
rect 13078 12356 13084 12368
rect 12474 12328 13084 12356
rect 12474 12325 12486 12328
rect 12428 12319 12486 12325
rect 13078 12316 13084 12328
rect 13136 12316 13142 12368
rect 15556 12359 15614 12365
rect 15556 12325 15568 12359
rect 15602 12356 15614 12359
rect 15838 12356 15844 12368
rect 15602 12328 15844 12356
rect 15602 12325 15614 12328
rect 15556 12319 15614 12325
rect 15838 12316 15844 12328
rect 15896 12316 15902 12368
rect 17586 12356 17592 12368
rect 17236 12328 17592 12356
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12257 6331 12291
rect 6273 12251 6331 12257
rect 6822 12248 6828 12300
rect 6880 12288 6886 12300
rect 6917 12291 6975 12297
rect 6917 12288 6929 12291
rect 6880 12260 6929 12288
rect 6880 12248 6886 12260
rect 6917 12257 6929 12260
rect 6963 12257 6975 12291
rect 6917 12251 6975 12257
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7561 12291 7619 12297
rect 7561 12288 7573 12291
rect 7064 12260 7573 12288
rect 7064 12248 7070 12260
rect 7561 12257 7573 12260
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8754 12288 8760 12300
rect 7975 12260 8760 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8754 12248 8760 12260
rect 8812 12288 8818 12300
rect 9490 12288 9496 12300
rect 8812 12260 9496 12288
rect 8812 12248 8818 12260
rect 9490 12248 9496 12260
rect 9548 12248 9554 12300
rect 10318 12248 10324 12300
rect 10376 12288 10382 12300
rect 10413 12291 10471 12297
rect 10413 12288 10425 12291
rect 10376 12260 10425 12288
rect 10376 12248 10382 12260
rect 10413 12257 10425 12260
rect 10459 12257 10471 12291
rect 10413 12251 10471 12257
rect 11517 12291 11575 12297
rect 11517 12257 11529 12291
rect 11563 12288 11575 12291
rect 11974 12288 11980 12300
rect 11563 12260 11980 12288
rect 11563 12257 11575 12260
rect 11517 12251 11575 12257
rect 11974 12248 11980 12260
rect 12032 12248 12038 12300
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12288 12219 12291
rect 12710 12288 12716 12300
rect 12207 12260 12716 12288
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 14458 12288 14464 12300
rect 14419 12260 14464 12288
rect 14458 12248 14464 12260
rect 14516 12248 14522 12300
rect 14642 12248 14648 12300
rect 14700 12288 14706 12300
rect 17236 12297 17264 12328
rect 17586 12316 17592 12328
rect 17644 12356 17650 12368
rect 17770 12356 17776 12368
rect 17644 12328 17776 12356
rect 17644 12316 17650 12328
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 14700 12260 15301 12288
rect 14700 12248 14706 12260
rect 15289 12257 15301 12260
rect 15335 12288 15347 12291
rect 17221 12291 17279 12297
rect 17221 12288 17233 12291
rect 15335 12260 17233 12288
rect 15335 12257 15347 12260
rect 15289 12251 15347 12257
rect 17221 12257 17233 12260
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 17488 12291 17546 12297
rect 17488 12257 17500 12291
rect 17534 12288 17546 12291
rect 18046 12288 18052 12300
rect 17534 12260 18052 12288
rect 17534 12257 17546 12260
rect 17488 12251 17546 12257
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 3418 12220 3424 12232
rect 2455 12192 3424 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3786 12180 3792 12232
rect 3844 12220 3850 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 3844 12192 4077 12220
rect 3844 12180 3850 12192
rect 4065 12189 4077 12192
rect 4111 12189 4123 12223
rect 5460 12220 5488 12248
rect 7101 12223 7159 12229
rect 7101 12220 7113 12223
rect 5460 12192 7113 12220
rect 4065 12183 4123 12189
rect 7101 12189 7113 12192
rect 7147 12220 7159 12223
rect 7190 12220 7196 12232
rect 7147 12192 7196 12220
rect 7147 12189 7159 12192
rect 7101 12183 7159 12189
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 11701 12223 11759 12229
rect 11701 12220 11713 12223
rect 10643 12192 11713 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 11701 12189 11713 12192
rect 11747 12189 11759 12223
rect 11701 12183 11759 12189
rect 10410 12112 10416 12164
rect 10468 12152 10474 12164
rect 10612 12152 10640 12183
rect 10468 12124 10640 12152
rect 11716 12152 11744 12183
rect 13630 12180 13636 12232
rect 13688 12220 13694 12232
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 13688 12192 14565 12220
rect 13688 12180 13694 12192
rect 14553 12189 14565 12192
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 11716 12124 11928 12152
rect 10468 12112 10474 12124
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 5445 12087 5503 12093
rect 5445 12084 5457 12087
rect 4856 12056 5457 12084
rect 4856 12044 4862 12056
rect 5445 12053 5457 12056
rect 5491 12053 5503 12087
rect 5445 12047 5503 12053
rect 5534 12044 5540 12096
rect 5592 12084 5598 12096
rect 5721 12087 5779 12093
rect 5721 12084 5733 12087
rect 5592 12056 5733 12084
rect 5592 12044 5598 12056
rect 5721 12053 5733 12056
rect 5767 12084 5779 12087
rect 5902 12084 5908 12096
rect 5767 12056 5908 12084
rect 5767 12053 5779 12056
rect 5721 12047 5779 12053
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 6086 12084 6092 12096
rect 6047 12056 6092 12084
rect 6086 12044 6092 12056
rect 6144 12044 6150 12096
rect 6546 12084 6552 12096
rect 6507 12056 6552 12084
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 10045 12087 10103 12093
rect 10045 12053 10057 12087
rect 10091 12084 10103 12087
rect 11054 12084 11060 12096
rect 10091 12056 11060 12084
rect 10091 12053 10103 12056
rect 10045 12047 10103 12053
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 11149 12087 11207 12093
rect 11149 12053 11161 12087
rect 11195 12084 11207 12087
rect 11790 12084 11796 12096
rect 11195 12056 11796 12084
rect 11195 12053 11207 12056
rect 11149 12047 11207 12053
rect 11790 12044 11796 12056
rect 11848 12044 11854 12096
rect 11900 12084 11928 12124
rect 14182 12112 14188 12164
rect 14240 12152 14246 12164
rect 14660 12152 14688 12248
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 15194 12220 15200 12232
rect 14783 12192 15200 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 15194 12180 15200 12192
rect 15252 12180 15258 12232
rect 18874 12220 18880 12232
rect 18835 12192 18880 12220
rect 18874 12180 18880 12192
rect 18932 12180 18938 12232
rect 14240 12124 14688 12152
rect 14240 12112 14246 12124
rect 13541 12087 13599 12093
rect 13541 12084 13553 12087
rect 11900 12056 13553 12084
rect 13541 12053 13553 12056
rect 13587 12053 13599 12087
rect 13541 12047 13599 12053
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 18601 12087 18659 12093
rect 18601 12084 18613 12087
rect 18196 12056 18613 12084
rect 18196 12044 18202 12056
rect 18601 12053 18613 12056
rect 18647 12084 18659 12087
rect 18782 12084 18788 12096
rect 18647 12056 18788 12084
rect 18647 12053 18659 12056
rect 18601 12047 18659 12053
rect 18782 12044 18788 12056
rect 18840 12044 18846 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 8478 11880 8484 11892
rect 4120 11852 8064 11880
rect 8439 11852 8484 11880
rect 4120 11840 4126 11852
rect 2130 11772 2136 11824
rect 2188 11812 2194 11824
rect 3881 11815 3939 11821
rect 3881 11812 3893 11815
rect 2188 11784 3893 11812
rect 2188 11772 2194 11784
rect 3881 11781 3893 11784
rect 3927 11781 3939 11815
rect 6546 11812 6552 11824
rect 3881 11775 3939 11781
rect 4356 11784 6552 11812
rect 2038 11744 2044 11756
rect 1999 11716 2044 11744
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 4356 11753 4384 11784
rect 6546 11772 6552 11784
rect 6604 11772 6610 11824
rect 8036 11812 8064 11852
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 11146 11880 11152 11892
rect 8588 11852 11152 11880
rect 8588 11812 8616 11852
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 11333 11883 11391 11889
rect 11333 11880 11345 11883
rect 11296 11852 11345 11880
rect 11296 11840 11302 11852
rect 11333 11849 11345 11852
rect 11379 11849 11391 11883
rect 13814 11880 13820 11892
rect 13775 11852 13820 11880
rect 11333 11843 11391 11849
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 15565 11883 15623 11889
rect 15565 11849 15577 11883
rect 15611 11880 15623 11883
rect 15838 11880 15844 11892
rect 15611 11852 15844 11880
rect 15611 11849 15623 11852
rect 15565 11843 15623 11849
rect 15838 11840 15844 11852
rect 15896 11840 15902 11892
rect 18049 11883 18107 11889
rect 18049 11849 18061 11883
rect 18095 11880 18107 11883
rect 19426 11880 19432 11892
rect 18095 11852 19432 11880
rect 18095 11849 18107 11852
rect 18049 11843 18107 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 8036 11784 8616 11812
rect 16117 11815 16175 11821
rect 16117 11781 16129 11815
rect 16163 11812 16175 11815
rect 17586 11812 17592 11824
rect 16163 11784 17592 11812
rect 16163 11781 16175 11784
rect 16117 11775 16175 11781
rect 17586 11772 17592 11784
rect 17644 11772 17650 11824
rect 4341 11747 4399 11753
rect 2832 11716 2877 11744
rect 2832 11704 2838 11716
rect 4341 11713 4353 11747
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11744 4583 11747
rect 4798 11744 4804 11756
rect 4571 11716 4804 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 5442 11744 5448 11756
rect 5403 11716 5448 11744
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 9677 11747 9735 11753
rect 9677 11744 9689 11747
rect 9548 11716 9689 11744
rect 9548 11704 9554 11716
rect 9677 11713 9689 11716
rect 9723 11713 9735 11747
rect 11790 11744 11796 11756
rect 11751 11716 11796 11744
rect 9677 11707 9735 11713
rect 11790 11704 11796 11716
rect 11848 11704 11854 11756
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11713 11943 11747
rect 12526 11744 12532 11756
rect 12487 11716 12532 11744
rect 11885 11707 11943 11713
rect 1765 11679 1823 11685
rect 1765 11645 1777 11679
rect 1811 11676 1823 11679
rect 1946 11676 1952 11688
rect 1811 11648 1952 11676
rect 1811 11645 1823 11648
rect 1765 11639 1823 11645
rect 1946 11636 1952 11648
rect 2004 11636 2010 11688
rect 2501 11679 2559 11685
rect 2501 11645 2513 11679
rect 2547 11676 2559 11679
rect 5718 11676 5724 11688
rect 2547 11648 5724 11676
rect 2547 11645 2559 11648
rect 2501 11639 2559 11645
rect 5718 11636 5724 11648
rect 5776 11636 5782 11688
rect 6178 11636 6184 11688
rect 6236 11676 6242 11688
rect 7101 11679 7159 11685
rect 7101 11676 7113 11679
rect 6236 11648 7113 11676
rect 6236 11636 6242 11648
rect 7101 11645 7113 11648
rect 7147 11645 7159 11679
rect 9766 11676 9772 11688
rect 7101 11639 7159 11645
rect 7208 11648 9772 11676
rect 4249 11611 4307 11617
rect 4249 11577 4261 11611
rect 4295 11608 4307 11611
rect 5261 11611 5319 11617
rect 4295 11580 4936 11608
rect 4295 11577 4307 11580
rect 4249 11571 4307 11577
rect 4908 11549 4936 11580
rect 5261 11577 5273 11611
rect 5307 11608 5319 11611
rect 5905 11611 5963 11617
rect 5905 11608 5917 11611
rect 5307 11580 5917 11608
rect 5307 11577 5319 11580
rect 5261 11571 5319 11577
rect 5905 11577 5917 11580
rect 5951 11577 5963 11611
rect 5905 11571 5963 11577
rect 6914 11568 6920 11620
rect 6972 11608 6978 11620
rect 7208 11608 7236 11648
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 9944 11679 10002 11685
rect 9944 11645 9956 11679
rect 9990 11676 10002 11679
rect 10410 11676 10416 11688
rect 9990 11648 10416 11676
rect 9990 11645 10002 11648
rect 9944 11639 10002 11645
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 11112 11648 11713 11676
rect 11112 11636 11118 11648
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11900 11676 11928 11707
rect 12526 11704 12532 11716
rect 12584 11704 12590 11756
rect 14182 11744 14188 11756
rect 14143 11716 14188 11744
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 18046 11704 18052 11756
rect 18104 11744 18110 11756
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 18104 11716 18613 11744
rect 18104 11704 18110 11716
rect 18601 11713 18613 11716
rect 18647 11744 18659 11747
rect 18690 11744 18696 11756
rect 18647 11716 18696 11744
rect 18647 11713 18659 11716
rect 18601 11707 18659 11713
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 11701 11639 11759 11645
rect 11808 11648 11928 11676
rect 13173 11679 13231 11685
rect 6972 11580 7236 11608
rect 6972 11568 6978 11580
rect 7282 11568 7288 11620
rect 7340 11617 7346 11620
rect 7340 11611 7404 11617
rect 7340 11577 7358 11611
rect 7392 11577 7404 11611
rect 7340 11571 7404 11577
rect 7340 11568 7346 11571
rect 8478 11568 8484 11620
rect 8536 11608 8542 11620
rect 8849 11611 8907 11617
rect 8849 11608 8861 11611
rect 8536 11580 8861 11608
rect 8536 11568 8542 11580
rect 8849 11577 8861 11580
rect 8895 11608 8907 11611
rect 10134 11608 10140 11620
rect 8895 11580 10140 11608
rect 8895 11577 8907 11580
rect 8849 11571 8907 11577
rect 10134 11568 10140 11580
rect 10192 11568 10198 11620
rect 11808 11608 11836 11648
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 11072 11580 11836 11608
rect 13188 11608 13216 11639
rect 14274 11636 14280 11688
rect 14332 11676 14338 11688
rect 16301 11679 16359 11685
rect 16301 11676 16313 11679
rect 14332 11648 16313 11676
rect 14332 11636 14338 11648
rect 16301 11645 16313 11648
rect 16347 11645 16359 11679
rect 16301 11639 16359 11645
rect 18417 11679 18475 11685
rect 18417 11645 18429 11679
rect 18463 11676 18475 11679
rect 18874 11676 18880 11688
rect 18463 11648 18880 11676
rect 18463 11645 18475 11648
rect 18417 11639 18475 11645
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 14292 11608 14320 11636
rect 13188 11580 14320 11608
rect 14452 11611 14510 11617
rect 11072 11552 11100 11580
rect 14452 11577 14464 11611
rect 14498 11608 14510 11611
rect 15194 11608 15200 11620
rect 14498 11580 15200 11608
rect 14498 11577 14510 11580
rect 14452 11571 14510 11577
rect 15194 11568 15200 11580
rect 15252 11608 15258 11620
rect 15470 11608 15476 11620
rect 15252 11580 15476 11608
rect 15252 11568 15258 11580
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 4893 11543 4951 11549
rect 4893 11509 4905 11543
rect 4939 11509 4951 11543
rect 4893 11503 4951 11509
rect 5353 11543 5411 11549
rect 5353 11509 5365 11543
rect 5399 11540 5411 11543
rect 5626 11540 5632 11552
rect 5399 11512 5632 11540
rect 5399 11509 5411 11512
rect 5353 11503 5411 11509
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 5994 11500 6000 11552
rect 6052 11540 6058 11552
rect 6365 11543 6423 11549
rect 6365 11540 6377 11543
rect 6052 11512 6377 11540
rect 6052 11500 6058 11512
rect 6365 11509 6377 11512
rect 6411 11540 6423 11543
rect 6822 11540 6828 11552
rect 6411 11512 6828 11540
rect 6411 11509 6423 11512
rect 6365 11503 6423 11509
rect 6822 11500 6828 11512
rect 6880 11540 6886 11552
rect 7466 11540 7472 11552
rect 6880 11512 7472 11540
rect 6880 11500 6886 11512
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 9125 11543 9183 11549
rect 9125 11540 9137 11543
rect 8444 11512 9137 11540
rect 8444 11500 8450 11512
rect 9125 11509 9137 11512
rect 9171 11509 9183 11543
rect 11054 11540 11060 11552
rect 11015 11512 11060 11540
rect 9125 11503 9183 11509
rect 11054 11500 11060 11512
rect 11112 11500 11118 11552
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12710 11540 12716 11552
rect 12492 11512 12716 11540
rect 12492 11500 12498 11512
rect 12710 11500 12716 11512
rect 12768 11540 12774 11552
rect 12989 11543 13047 11549
rect 12989 11540 13001 11543
rect 12768 11512 13001 11540
rect 12768 11500 12774 11512
rect 12989 11509 13001 11512
rect 13035 11509 13047 11543
rect 13446 11540 13452 11552
rect 13407 11512 13452 11540
rect 12989 11503 13047 11509
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 17494 11500 17500 11552
rect 17552 11540 17558 11552
rect 17589 11543 17647 11549
rect 17589 11540 17601 11543
rect 17552 11512 17601 11540
rect 17552 11500 17558 11512
rect 17589 11509 17601 11512
rect 17635 11540 17647 11543
rect 18509 11543 18567 11549
rect 18509 11540 18521 11543
rect 17635 11512 18521 11540
rect 17635 11509 17647 11512
rect 17589 11503 17647 11509
rect 18509 11509 18521 11512
rect 18555 11509 18567 11543
rect 18509 11503 18567 11509
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 1946 11336 1952 11348
rect 1907 11308 1952 11336
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 2961 11339 3019 11345
rect 2961 11336 2973 11339
rect 2455 11308 2973 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 2961 11305 2973 11308
rect 3007 11305 3019 11339
rect 2961 11299 3019 11305
rect 3421 11339 3479 11345
rect 3421 11305 3433 11339
rect 3467 11336 3479 11339
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 3467 11308 4077 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 4065 11305 4077 11308
rect 4111 11305 4123 11339
rect 4065 11299 4123 11305
rect 4525 11339 4583 11345
rect 4525 11305 4537 11339
rect 4571 11336 4583 11339
rect 4890 11336 4896 11348
rect 4571 11308 4896 11336
rect 4571 11305 4583 11308
rect 4525 11299 4583 11305
rect 4890 11296 4896 11308
rect 4948 11296 4954 11348
rect 6641 11339 6699 11345
rect 6641 11305 6653 11339
rect 6687 11336 6699 11339
rect 7558 11336 7564 11348
rect 6687 11308 7564 11336
rect 6687 11305 6699 11308
rect 6641 11299 6699 11305
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 8938 11336 8944 11348
rect 7699 11308 8944 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 9033 11339 9091 11345
rect 9033 11305 9045 11339
rect 9079 11336 9091 11339
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 9079 11308 9137 11336
rect 9079 11305 9091 11308
rect 9033 11299 9091 11305
rect 9125 11305 9137 11308
rect 9171 11336 9183 11339
rect 9490 11336 9496 11348
rect 9171 11308 9496 11336
rect 9171 11305 9183 11308
rect 9125 11299 9183 11305
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 10318 11336 10324 11348
rect 10279 11308 10324 11336
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 12618 11336 12624 11348
rect 12579 11308 12624 11336
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 13630 11336 13636 11348
rect 13591 11308 13636 11336
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 13872 11308 14105 11336
rect 13872 11296 13878 11308
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 14093 11299 14151 11305
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 14645 11339 14703 11345
rect 14645 11336 14657 11339
rect 14516 11308 14657 11336
rect 14516 11296 14522 11308
rect 14645 11305 14657 11308
rect 14691 11305 14703 11339
rect 18877 11339 18935 11345
rect 18877 11336 18889 11339
rect 14645 11299 14703 11305
rect 16684 11308 18889 11336
rect 3970 11228 3976 11280
rect 4028 11268 4034 11280
rect 6914 11268 6920 11280
rect 4028 11240 6920 11268
rect 4028 11228 4034 11240
rect 6914 11228 6920 11240
rect 6972 11228 6978 11280
rect 7006 11228 7012 11280
rect 7064 11268 7070 11280
rect 8113 11271 8171 11277
rect 7064 11240 7109 11268
rect 7064 11228 7070 11240
rect 8113 11237 8125 11271
rect 8159 11268 8171 11271
rect 8478 11268 8484 11280
rect 8159 11240 8484 11268
rect 8159 11237 8171 11240
rect 8113 11231 8171 11237
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 8570 11228 8576 11280
rect 8628 11268 8634 11280
rect 8665 11271 8723 11277
rect 8665 11268 8677 11271
rect 8628 11240 8677 11268
rect 8628 11228 8634 11240
rect 8665 11237 8677 11240
rect 8711 11237 8723 11271
rect 12434 11268 12440 11280
rect 8665 11231 8723 11237
rect 10980 11240 12440 11268
rect 2314 11200 2320 11212
rect 2275 11172 2320 11200
rect 2314 11160 2320 11172
rect 2372 11160 2378 11212
rect 3329 11203 3387 11209
rect 3329 11169 3341 11203
rect 3375 11200 3387 11203
rect 4062 11200 4068 11212
rect 3375 11172 4068 11200
rect 3375 11169 3387 11172
rect 3329 11163 3387 11169
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4338 11160 4344 11212
rect 4396 11200 4402 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4396 11172 4445 11200
rect 4396 11160 4402 11172
rect 4433 11169 4445 11172
rect 4479 11200 4491 11203
rect 5445 11203 5503 11209
rect 5445 11200 5457 11203
rect 4479 11172 5457 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 5445 11169 5457 11172
rect 5491 11200 5503 11203
rect 5994 11200 6000 11212
rect 5491 11172 6000 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 6086 11160 6092 11212
rect 6144 11200 6150 11212
rect 6365 11203 6423 11209
rect 6365 11200 6377 11203
rect 6144 11172 6377 11200
rect 6144 11160 6150 11172
rect 6365 11169 6377 11172
rect 6411 11200 6423 11203
rect 6411 11172 7411 11200
rect 6411 11169 6423 11172
rect 6365 11163 6423 11169
rect 2593 11135 2651 11141
rect 2593 11101 2605 11135
rect 2639 11132 2651 11135
rect 2682 11132 2688 11144
rect 2639 11104 2688 11132
rect 2639 11101 2651 11104
rect 2593 11095 2651 11101
rect 2682 11092 2688 11104
rect 2740 11092 2746 11144
rect 3513 11135 3571 11141
rect 3513 11101 3525 11135
rect 3559 11101 3571 11135
rect 3513 11095 3571 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11132 5227 11135
rect 5626 11132 5632 11144
rect 5215 11104 5632 11132
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 2406 11024 2412 11076
rect 2464 11064 2470 11076
rect 3528 11064 3556 11095
rect 4154 11064 4160 11076
rect 2464 11036 4160 11064
rect 2464 11024 2470 11036
rect 4154 11024 4160 11036
rect 4212 11024 4218 11076
rect 4724 10996 4752 11095
rect 5626 11092 5632 11104
rect 5684 11132 5690 11144
rect 5813 11135 5871 11141
rect 5813 11132 5825 11135
rect 5684 11104 5825 11132
rect 5684 11092 5690 11104
rect 5813 11101 5825 11104
rect 5859 11132 5871 11135
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 5859 11104 7113 11132
rect 5859 11101 5871 11104
rect 5813 11095 5871 11101
rect 7101 11101 7113 11104
rect 7147 11101 7159 11135
rect 7282 11132 7288 11144
rect 7195 11104 7288 11132
rect 7101 11095 7159 11101
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 7383 11132 7411 11172
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 8018 11200 8024 11212
rect 7524 11172 8024 11200
rect 7524 11160 7530 11172
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 10980 11209 11008 11240
rect 12434 11228 12440 11240
rect 12492 11228 12498 11280
rect 15924 11271 15982 11277
rect 15924 11237 15936 11271
rect 15970 11268 15982 11271
rect 16114 11268 16120 11280
rect 15970 11240 16120 11268
rect 15970 11237 15982 11240
rect 15924 11231 15982 11237
rect 16114 11228 16120 11240
rect 16172 11268 16178 11280
rect 16684 11268 16712 11308
rect 18877 11305 18889 11308
rect 18923 11305 18935 11339
rect 18877 11299 18935 11305
rect 16172 11240 16712 11268
rect 17764 11271 17822 11277
rect 16172 11228 16178 11240
rect 17764 11237 17776 11271
rect 17810 11268 17822 11271
rect 18138 11268 18144 11280
rect 17810 11240 18144 11268
rect 17810 11237 17822 11240
rect 17764 11231 17822 11237
rect 18138 11228 18144 11240
rect 18196 11228 18202 11280
rect 11238 11209 11244 11212
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 8128 11172 9321 11200
rect 8128 11132 8156 11172
rect 9309 11169 9321 11172
rect 9355 11169 9367 11203
rect 9309 11163 9367 11169
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11232 11163 11244 11209
rect 11296 11200 11302 11212
rect 11296 11172 11332 11200
rect 11238 11160 11244 11163
rect 11296 11160 11302 11172
rect 12526 11160 12532 11212
rect 12584 11200 12590 11212
rect 12989 11203 13047 11209
rect 12989 11200 13001 11203
rect 12584 11172 13001 11200
rect 12584 11160 12590 11172
rect 12989 11169 13001 11172
rect 13035 11169 13047 11203
rect 12989 11163 13047 11169
rect 13446 11160 13452 11212
rect 13504 11200 13510 11212
rect 14001 11203 14059 11209
rect 14001 11200 14013 11203
rect 13504 11172 14013 11200
rect 13504 11160 13510 11172
rect 14001 11169 14013 11172
rect 14047 11169 14059 11203
rect 14001 11163 14059 11169
rect 15657 11203 15715 11209
rect 15657 11169 15669 11203
rect 15703 11200 15715 11203
rect 16298 11200 16304 11212
rect 15703 11172 16304 11200
rect 15703 11169 15715 11172
rect 15657 11163 15715 11169
rect 16298 11160 16304 11172
rect 16356 11200 16362 11212
rect 17497 11203 17555 11209
rect 17497 11200 17509 11203
rect 16356 11172 17509 11200
rect 16356 11160 16362 11172
rect 17497 11169 17509 11172
rect 17543 11200 17555 11203
rect 17586 11200 17592 11212
rect 17543 11172 17592 11200
rect 17543 11169 17555 11172
rect 17497 11163 17555 11169
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 7383 11104 8156 11132
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 6178 11064 6184 11076
rect 6139 11036 6184 11064
rect 6178 11024 6184 11036
rect 6236 11024 6242 11076
rect 7300 11064 7328 11092
rect 8110 11064 8116 11076
rect 7300 11036 8116 11064
rect 8110 11024 8116 11036
rect 8168 11064 8174 11076
rect 8211 11064 8239 11095
rect 12158 11092 12164 11144
rect 12216 11132 12222 11144
rect 13081 11135 13139 11141
rect 13081 11132 13093 11135
rect 12216 11104 13093 11132
rect 12216 11092 12222 11104
rect 13081 11101 13093 11104
rect 13127 11101 13139 11135
rect 13081 11095 13139 11101
rect 13173 11135 13231 11141
rect 13173 11101 13185 11135
rect 13219 11101 13231 11135
rect 13173 11095 13231 11101
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 14366 11132 14372 11144
rect 14323 11104 14372 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 8168 11036 8239 11064
rect 8168 11024 8174 11036
rect 8478 11024 8484 11076
rect 8536 11064 8542 11076
rect 9033 11067 9091 11073
rect 9033 11064 9045 11067
rect 8536 11036 9045 11064
rect 8536 11024 8542 11036
rect 9033 11033 9045 11036
rect 9079 11033 9091 11067
rect 9398 11064 9404 11076
rect 9033 11027 9091 11033
rect 9140 11036 9404 11064
rect 4798 10996 4804 11008
rect 4711 10968 4804 10996
rect 4798 10956 4804 10968
rect 4856 10996 4862 11008
rect 9140 10996 9168 11036
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 12345 11067 12403 11073
rect 12345 11033 12357 11067
rect 12391 11064 12403 11067
rect 12710 11064 12716 11076
rect 12391 11036 12716 11064
rect 12391 11033 12403 11036
rect 12345 11027 12403 11033
rect 12710 11024 12716 11036
rect 12768 11064 12774 11076
rect 13188 11064 13216 11095
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 12768 11036 13216 11064
rect 12768 11024 12774 11036
rect 4856 10968 9168 10996
rect 4856 10956 4862 10968
rect 9214 10956 9220 11008
rect 9272 10996 9278 11008
rect 13998 10996 14004 11008
rect 9272 10968 14004 10996
rect 9272 10956 9278 10968
rect 13998 10956 14004 10968
rect 14056 10956 14062 11008
rect 17034 10996 17040 11008
rect 16995 10968 17040 10996
rect 17034 10956 17040 10968
rect 17092 10956 17098 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 2314 10792 2320 10804
rect 1811 10764 2320 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 2314 10752 2320 10764
rect 2372 10752 2378 10804
rect 4154 10792 4160 10804
rect 4115 10764 4160 10792
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4525 10795 4583 10801
rect 4525 10761 4537 10795
rect 4571 10792 4583 10795
rect 4890 10792 4896 10804
rect 4571 10764 4896 10792
rect 4571 10761 4583 10764
rect 4525 10755 4583 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 5718 10792 5724 10804
rect 5679 10764 5724 10792
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 5828 10764 7788 10792
rect 3878 10684 3884 10736
rect 3936 10724 3942 10736
rect 5828 10724 5856 10764
rect 6454 10724 6460 10736
rect 3936 10696 5856 10724
rect 6288 10696 6460 10724
rect 3936 10684 3942 10696
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 2409 10659 2467 10665
rect 2409 10656 2421 10659
rect 2372 10628 2421 10656
rect 2372 10616 2378 10628
rect 2409 10625 2421 10628
rect 2455 10625 2467 10659
rect 2409 10619 2467 10625
rect 4522 10616 4528 10668
rect 4580 10656 4586 10668
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4580 10628 4905 10656
rect 4580 10616 4586 10628
rect 4893 10625 4905 10628
rect 4939 10656 4951 10659
rect 6288 10656 6316 10696
rect 6454 10684 6460 10696
rect 6512 10684 6518 10736
rect 7760 10724 7788 10764
rect 8110 10752 8116 10804
rect 8168 10792 8174 10804
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 8168 10764 8217 10792
rect 8168 10752 8174 10764
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 9214 10792 9220 10804
rect 8205 10755 8263 10761
rect 8312 10764 9220 10792
rect 8312 10724 8340 10764
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 9398 10752 9404 10804
rect 9456 10792 9462 10804
rect 10870 10792 10876 10804
rect 9456 10764 10876 10792
rect 9456 10752 9462 10764
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 11296 10764 11529 10792
rect 11296 10752 11302 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 13817 10795 13875 10801
rect 13817 10761 13829 10795
rect 13863 10792 13875 10795
rect 14366 10792 14372 10804
rect 13863 10764 14372 10792
rect 13863 10761 13875 10764
rect 13817 10755 13875 10761
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 15470 10792 15476 10804
rect 15431 10764 15476 10792
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 17678 10724 17684 10736
rect 7760 10696 8340 10724
rect 17639 10696 17684 10724
rect 17678 10684 17684 10696
rect 17736 10684 17742 10736
rect 4939 10628 6316 10656
rect 6365 10659 6423 10665
rect 4939 10625 4951 10628
rect 4893 10619 4951 10625
rect 6365 10625 6377 10659
rect 6411 10656 6423 10659
rect 6730 10656 6736 10668
rect 6411 10628 6736 10656
rect 6411 10625 6423 10628
rect 6365 10619 6423 10625
rect 6730 10616 6736 10628
rect 6788 10656 6794 10668
rect 6788 10628 6960 10656
rect 6788 10616 6794 10628
rect 2774 10588 2780 10600
rect 2735 10560 2780 10588
rect 2774 10548 2780 10560
rect 2832 10548 2838 10600
rect 5258 10588 5264 10600
rect 5171 10560 5264 10588
rect 5258 10548 5264 10560
rect 5316 10588 5322 10600
rect 6638 10588 6644 10600
rect 5316 10560 6644 10588
rect 5316 10548 5322 10560
rect 6638 10548 6644 10560
rect 6696 10548 6702 10600
rect 6822 10588 6828 10600
rect 6783 10560 6828 10588
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 6932 10588 6960 10628
rect 9490 10616 9496 10668
rect 9548 10656 9554 10668
rect 10137 10659 10195 10665
rect 10137 10656 10149 10659
rect 9548 10628 10149 10656
rect 9548 10616 9554 10628
rect 10137 10625 10149 10628
rect 10183 10625 10195 10659
rect 16298 10656 16304 10668
rect 16259 10628 16304 10656
rect 10137 10619 10195 10625
rect 16298 10616 16304 10628
rect 16356 10616 16362 10668
rect 7081 10591 7139 10597
rect 7081 10588 7093 10591
rect 6932 10560 7093 10588
rect 7081 10557 7093 10560
rect 7127 10557 7139 10591
rect 7081 10551 7139 10557
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 8478 10588 8484 10600
rect 7708 10560 8484 10588
rect 7708 10548 7714 10560
rect 8478 10548 8484 10560
rect 8536 10548 8542 10600
rect 8588 10560 9996 10588
rect 3044 10523 3102 10529
rect 3044 10489 3056 10523
rect 3090 10520 3102 10523
rect 3510 10520 3516 10532
rect 3090 10492 3516 10520
rect 3090 10489 3102 10492
rect 3044 10483 3102 10489
rect 3510 10480 3516 10492
rect 3568 10480 3574 10532
rect 3970 10480 3976 10532
rect 4028 10520 4034 10532
rect 8588 10520 8616 10560
rect 4028 10492 8616 10520
rect 8748 10523 8806 10529
rect 4028 10480 4034 10492
rect 8748 10489 8760 10523
rect 8794 10520 8806 10523
rect 8938 10520 8944 10532
rect 8794 10492 8944 10520
rect 8794 10489 8806 10492
rect 8748 10483 8806 10489
rect 8938 10480 8944 10492
rect 8996 10480 9002 10532
rect 2130 10452 2136 10464
rect 2091 10424 2136 10452
rect 2130 10412 2136 10424
rect 2188 10412 2194 10464
rect 2225 10455 2283 10461
rect 2225 10421 2237 10455
rect 2271 10452 2283 10455
rect 2866 10452 2872 10464
rect 2271 10424 2872 10452
rect 2271 10421 2283 10424
rect 2225 10415 2283 10421
rect 2866 10412 2872 10424
rect 2924 10412 2930 10464
rect 6086 10452 6092 10464
rect 6047 10424 6092 10452
rect 6086 10412 6092 10424
rect 6144 10412 6150 10464
rect 6181 10455 6239 10461
rect 6181 10421 6193 10455
rect 6227 10452 6239 10455
rect 7374 10452 7380 10464
rect 6227 10424 7380 10452
rect 6227 10421 6239 10424
rect 6181 10415 6239 10421
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 9861 10455 9919 10461
rect 9861 10452 9873 10455
rect 8260 10424 9873 10452
rect 8260 10412 8266 10424
rect 9861 10421 9873 10424
rect 9907 10421 9919 10455
rect 9968 10452 9996 10560
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12710 10597 12716 10600
rect 12704 10588 12716 10597
rect 12492 10560 12537 10588
rect 12671 10560 12716 10588
rect 12492 10548 12498 10560
rect 12704 10551 12716 10560
rect 12710 10548 12716 10551
rect 12768 10548 12774 10600
rect 14366 10597 14372 10600
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10588 13967 10591
rect 14093 10591 14151 10597
rect 14093 10588 14105 10591
rect 13955 10560 14105 10588
rect 13955 10557 13967 10560
rect 13909 10551 13967 10557
rect 14093 10557 14105 10560
rect 14139 10557 14151 10591
rect 14360 10588 14372 10597
rect 14327 10560 14372 10588
rect 14093 10551 14151 10557
rect 14360 10551 14372 10560
rect 14366 10548 14372 10551
rect 14424 10548 14430 10600
rect 16568 10591 16626 10597
rect 16568 10557 16580 10591
rect 16614 10588 16626 10591
rect 17034 10588 17040 10600
rect 16614 10560 17040 10588
rect 16614 10557 16626 10560
rect 16568 10551 16626 10557
rect 17034 10548 17040 10560
rect 17092 10548 17098 10600
rect 10404 10523 10462 10529
rect 10404 10489 10416 10523
rect 10450 10520 10462 10523
rect 11054 10520 11060 10532
rect 10450 10492 11060 10520
rect 10450 10489 10462 10492
rect 10404 10483 10462 10489
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 11885 10523 11943 10529
rect 11885 10489 11897 10523
rect 11931 10520 11943 10523
rect 12526 10520 12532 10532
rect 11931 10492 12532 10520
rect 11931 10489 11943 10492
rect 11885 10483 11943 10489
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 12250 10452 12256 10464
rect 9968 10424 12256 10452
rect 9861 10415 9919 10421
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 13909 10455 13967 10461
rect 13909 10452 13921 10455
rect 12492 10424 13921 10452
rect 12492 10412 12498 10424
rect 13909 10421 13921 10424
rect 13955 10421 13967 10455
rect 18046 10452 18052 10464
rect 18007 10424 18052 10452
rect 13909 10415 13967 10421
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 2130 10208 2136 10260
rect 2188 10248 2194 10260
rect 3421 10251 3479 10257
rect 3421 10248 3433 10251
rect 2188 10220 3433 10248
rect 2188 10208 2194 10220
rect 3421 10217 3433 10220
rect 3467 10217 3479 10251
rect 4062 10248 4068 10260
rect 4023 10220 4068 10248
rect 3421 10211 3479 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4522 10248 4528 10260
rect 4483 10220 4528 10248
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 4982 10208 4988 10260
rect 5040 10248 5046 10260
rect 6730 10248 6736 10260
rect 5040 10220 6592 10248
rect 6691 10220 6736 10248
rect 5040 10208 5046 10220
rect 2032 10183 2090 10189
rect 2032 10149 2044 10183
rect 2078 10180 2090 10183
rect 2314 10180 2320 10192
rect 2078 10152 2320 10180
rect 2078 10149 2090 10152
rect 2032 10143 2090 10149
rect 2314 10140 2320 10152
rect 2372 10140 2378 10192
rect 3786 10180 3792 10192
rect 3252 10152 3792 10180
rect 3252 10124 3280 10152
rect 3786 10140 3792 10152
rect 3844 10180 3850 10192
rect 6178 10180 6184 10192
rect 3844 10152 6184 10180
rect 3844 10140 3850 10152
rect 1765 10115 1823 10121
rect 1765 10081 1777 10115
rect 1811 10112 1823 10115
rect 2774 10112 2780 10124
rect 1811 10084 2780 10112
rect 1811 10081 1823 10084
rect 1765 10075 1823 10081
rect 2774 10072 2780 10084
rect 2832 10112 2838 10124
rect 3234 10112 3240 10124
rect 2832 10084 3240 10112
rect 2832 10072 2838 10084
rect 3234 10072 3240 10084
rect 3292 10072 3298 10124
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10112 4491 10115
rect 5258 10112 5264 10124
rect 4479 10084 5264 10112
rect 4479 10081 4491 10084
rect 4433 10075 4491 10081
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 5368 10121 5396 10152
rect 6178 10140 6184 10152
rect 6236 10140 6242 10192
rect 6564 10180 6592 10220
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 7374 10248 7380 10260
rect 7335 10220 7380 10248
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 7745 10251 7803 10257
rect 7745 10217 7757 10251
rect 7791 10248 7803 10251
rect 8389 10251 8447 10257
rect 8389 10248 8401 10251
rect 7791 10220 8401 10248
rect 7791 10217 7803 10220
rect 7745 10211 7803 10217
rect 8389 10217 8401 10220
rect 8435 10217 8447 10251
rect 8389 10211 8447 10217
rect 9677 10251 9735 10257
rect 9677 10217 9689 10251
rect 9723 10248 9735 10251
rect 9858 10248 9864 10260
rect 9723 10220 9864 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 10042 10248 10048 10260
rect 10003 10220 10048 10248
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10217 10931 10251
rect 10873 10211 10931 10217
rect 7009 10183 7067 10189
rect 7009 10180 7021 10183
rect 6564 10152 7021 10180
rect 7009 10149 7021 10152
rect 7055 10180 7067 10183
rect 8757 10183 8815 10189
rect 8757 10180 8769 10183
rect 7055 10152 8769 10180
rect 7055 10149 7067 10152
rect 7009 10143 7067 10149
rect 8757 10149 8769 10152
rect 8803 10149 8815 10183
rect 10888 10180 10916 10211
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 12253 10251 12311 10257
rect 12253 10248 12265 10251
rect 12032 10220 12265 10248
rect 12032 10208 12038 10220
rect 12253 10217 12265 10220
rect 12299 10217 12311 10251
rect 12253 10211 12311 10217
rect 15473 10251 15531 10257
rect 15473 10217 15485 10251
rect 15519 10217 15531 10251
rect 15473 10211 15531 10217
rect 16577 10251 16635 10257
rect 16577 10217 16589 10251
rect 16623 10248 16635 10251
rect 16850 10248 16856 10260
rect 16623 10220 16856 10248
rect 16623 10217 16635 10220
rect 16577 10211 16635 10217
rect 12158 10180 12164 10192
rect 10888 10152 12164 10180
rect 8757 10143 8815 10149
rect 12158 10140 12164 10152
rect 12216 10140 12222 10192
rect 15488 10180 15516 10211
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 16945 10251 17003 10257
rect 16945 10217 16957 10251
rect 16991 10248 17003 10251
rect 18046 10248 18052 10260
rect 16991 10220 18052 10248
rect 16991 10217 17003 10220
rect 16945 10211 17003 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 17037 10183 17095 10189
rect 17037 10180 17049 10183
rect 15488 10152 17049 10180
rect 17037 10149 17049 10152
rect 17083 10149 17095 10183
rect 17037 10143 17095 10149
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10081 5411 10115
rect 5353 10075 5411 10081
rect 5620 10115 5678 10121
rect 5620 10081 5632 10115
rect 5666 10112 5678 10115
rect 5666 10084 7972 10112
rect 5666 10081 5678 10084
rect 5620 10075 5678 10081
rect 7944 10056 7972 10084
rect 8956 10084 10272 10112
rect 8956 10056 8984 10084
rect 3510 10004 3516 10056
rect 3568 10044 3574 10056
rect 4709 10047 4767 10053
rect 4709 10044 4721 10047
rect 3568 10016 4721 10044
rect 3568 10004 3574 10016
rect 4709 10013 4721 10016
rect 4755 10044 4767 10047
rect 4798 10044 4804 10056
rect 4755 10016 4804 10044
rect 4755 10013 4767 10016
rect 4709 10007 4767 10013
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10013 7895 10047
rect 7837 10007 7895 10013
rect 7852 9976 7880 10007
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 8021 10047 8079 10053
rect 8021 10044 8033 10047
rect 7984 10016 8033 10044
rect 7984 10004 7990 10016
rect 8021 10013 8033 10016
rect 8067 10044 8079 10047
rect 8202 10044 8208 10056
rect 8067 10016 8208 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 8846 10044 8852 10056
rect 8807 10016 8852 10044
rect 8846 10004 8852 10016
rect 8904 10004 8910 10056
rect 8938 10004 8944 10056
rect 8996 10044 9002 10056
rect 10244 10053 10272 10084
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 10744 10084 11253 10112
rect 10744 10072 10750 10084
rect 11241 10081 11253 10084
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 11333 10115 11391 10121
rect 11333 10081 11345 10115
rect 11379 10112 11391 10115
rect 11379 10084 12020 10112
rect 11379 10081 11391 10084
rect 11333 10075 11391 10081
rect 11992 10053 12020 10084
rect 12250 10072 12256 10124
rect 12308 10112 12314 10124
rect 13446 10112 13452 10124
rect 12308 10084 13452 10112
rect 12308 10072 12314 10084
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 14734 10072 14740 10124
rect 14792 10112 14798 10124
rect 14921 10115 14979 10121
rect 14921 10112 14933 10115
rect 14792 10084 14933 10112
rect 14792 10072 14798 10084
rect 14921 10081 14933 10084
rect 14967 10112 14979 10115
rect 15841 10115 15899 10121
rect 15841 10112 15853 10115
rect 14967 10084 15853 10112
rect 14967 10081 14979 10084
rect 14921 10075 14979 10081
rect 15841 10081 15853 10084
rect 15887 10081 15899 10115
rect 15841 10075 15899 10081
rect 10137 10047 10195 10053
rect 8996 10016 9041 10044
rect 8996 10004 9002 10016
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 11977 10047 12035 10053
rect 11977 10013 11989 10047
rect 12023 10044 12035 10047
rect 13538 10044 13544 10056
rect 12023 10016 13544 10044
rect 12023 10013 12035 10016
rect 11977 10007 12035 10013
rect 9858 9976 9864 9988
rect 7852 9948 9864 9976
rect 9858 9936 9864 9948
rect 9916 9936 9922 9988
rect 10152 9976 10180 10007
rect 11146 9976 11152 9988
rect 10152 9948 11152 9976
rect 11146 9936 11152 9948
rect 11204 9936 11210 9988
rect 11238 9936 11244 9988
rect 11296 9976 11302 9988
rect 11440 9976 11468 10007
rect 13538 10004 13544 10016
rect 13596 10044 13602 10056
rect 15102 10044 15108 10056
rect 13596 10016 15108 10044
rect 13596 10004 13602 10016
rect 15102 10004 15108 10016
rect 15160 10044 15166 10056
rect 15933 10047 15991 10053
rect 15933 10044 15945 10047
rect 15160 10016 15945 10044
rect 15160 10004 15166 10016
rect 15933 10013 15945 10016
rect 15979 10013 15991 10047
rect 16114 10044 16120 10056
rect 16075 10016 16120 10044
rect 15933 10007 15991 10013
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 17126 10044 17132 10056
rect 17087 10016 17132 10044
rect 17126 10004 17132 10016
rect 17184 10004 17190 10056
rect 11296 9948 11468 9976
rect 11296 9936 11302 9948
rect 2682 9868 2688 9920
rect 2740 9908 2746 9920
rect 3145 9911 3203 9917
rect 3145 9908 3157 9911
rect 2740 9880 3157 9908
rect 2740 9868 2746 9880
rect 3145 9877 3157 9880
rect 3191 9877 3203 9911
rect 3145 9871 3203 9877
rect 9582 9868 9588 9920
rect 9640 9908 9646 9920
rect 14090 9908 14096 9920
rect 9640 9880 14096 9908
rect 9640 9868 9646 9880
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 2866 9704 2872 9716
rect 2827 9676 2872 9704
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 6144 9676 6837 9704
rect 6144 9664 6150 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 6825 9667 6883 9673
rect 8938 9664 8944 9716
rect 8996 9704 9002 9716
rect 9401 9707 9459 9713
rect 9401 9704 9413 9707
rect 8996 9676 9413 9704
rect 8996 9664 9002 9676
rect 9401 9673 9413 9676
rect 9447 9673 9459 9707
rect 9401 9667 9459 9673
rect 9769 9707 9827 9713
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 10042 9704 10048 9716
rect 9815 9676 10048 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 15102 9704 15108 9716
rect 15063 9676 15108 9704
rect 15102 9664 15108 9676
rect 15160 9664 15166 9716
rect 1854 9596 1860 9648
rect 1912 9636 1918 9648
rect 1949 9639 2007 9645
rect 1949 9636 1961 9639
rect 1912 9608 1961 9636
rect 1912 9596 1918 9608
rect 1949 9605 1961 9608
rect 1995 9605 2007 9639
rect 11146 9636 11152 9648
rect 11107 9608 11152 9636
rect 1949 9599 2007 9605
rect 11146 9596 11152 9608
rect 11204 9596 11210 9648
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9568 2651 9571
rect 2774 9568 2780 9580
rect 2639 9540 2780 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 2774 9528 2780 9540
rect 2832 9568 2838 9580
rect 3326 9568 3332 9580
rect 2832 9540 3332 9568
rect 2832 9528 2838 9540
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 3510 9568 3516 9580
rect 3471 9540 3516 9568
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 4798 9568 4804 9580
rect 4759 9540 4804 9568
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 7469 9571 7527 9577
rect 6972 9540 7420 9568
rect 6972 9528 6978 9540
rect 7392 9512 7420 9540
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 7926 9568 7932 9580
rect 7515 9540 7932 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 10686 9568 10692 9580
rect 9824 9540 10692 9568
rect 9824 9528 9830 9540
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 1762 9500 1768 9512
rect 1723 9472 1768 9500
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 4028 9472 7328 9500
rect 4028 9460 4034 9472
rect 3881 9435 3939 9441
rect 3881 9432 3893 9435
rect 3252 9404 3893 9432
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 3252 9373 3280 9404
rect 3881 9401 3893 9404
rect 3927 9432 3939 9435
rect 5626 9432 5632 9444
rect 3927 9404 5632 9432
rect 3927 9401 3939 9404
rect 3881 9395 3939 9401
rect 5626 9392 5632 9404
rect 5684 9392 5690 9444
rect 6273 9435 6331 9441
rect 6273 9401 6285 9435
rect 6319 9432 6331 9435
rect 7193 9435 7251 9441
rect 7193 9432 7205 9435
rect 6319 9404 7205 9432
rect 6319 9401 6331 9404
rect 6273 9395 6331 9401
rect 7193 9401 7205 9404
rect 7239 9401 7251 9435
rect 7300 9432 7328 9472
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 7650 9500 7656 9512
rect 7432 9472 7656 9500
rect 7432 9460 7438 9472
rect 7650 9460 7656 9472
rect 7708 9500 7714 9512
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7708 9472 8033 9500
rect 7708 9460 7714 9472
rect 8021 9469 8033 9472
rect 8067 9469 8079 9503
rect 17402 9500 17408 9512
rect 8021 9463 8079 9469
rect 8128 9472 17408 9500
rect 8128 9432 8156 9472
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 7300 9404 8156 9432
rect 8288 9435 8346 9441
rect 7193 9395 7251 9401
rect 8288 9401 8300 9435
rect 8334 9432 8346 9435
rect 8662 9432 8668 9444
rect 8334 9404 8668 9432
rect 8334 9401 8346 9404
rect 8288 9395 8346 9401
rect 8662 9392 8668 9404
rect 8720 9392 8726 9444
rect 3237 9367 3295 9373
rect 3237 9364 3249 9367
rect 3108 9336 3249 9364
rect 3108 9324 3114 9336
rect 3237 9333 3249 9336
rect 3283 9333 3295 9367
rect 4246 9364 4252 9376
rect 4207 9336 4252 9364
rect 3237 9327 3295 9333
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 4614 9364 4620 9376
rect 4575 9336 4620 9364
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 4709 9367 4767 9373
rect 4709 9333 4721 9367
rect 4755 9364 4767 9367
rect 4890 9364 4896 9376
rect 4755 9336 4896 9364
rect 4755 9333 4767 9336
rect 4709 9327 4767 9333
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 7282 9364 7288 9376
rect 7243 9336 7288 9364
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 11146 9324 11152 9376
rect 11204 9364 11210 9376
rect 13354 9364 13360 9376
rect 11204 9336 13360 9364
rect 11204 9324 11210 9336
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 1949 9163 2007 9169
rect 1949 9160 1961 9163
rect 1452 9132 1961 9160
rect 1452 9120 1458 9132
rect 1949 9129 1961 9132
rect 1995 9129 2007 9163
rect 4614 9160 4620 9172
rect 4575 9132 4620 9160
rect 1949 9123 2007 9129
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 7929 9163 7987 9169
rect 7929 9129 7941 9163
rect 7975 9160 7987 9163
rect 8202 9160 8208 9172
rect 7975 9132 8208 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 8386 9120 8392 9172
rect 8444 9160 8450 9172
rect 8573 9163 8631 9169
rect 8573 9160 8585 9163
rect 8444 9132 8585 9160
rect 8444 9120 8450 9132
rect 8573 9129 8585 9132
rect 8619 9129 8631 9163
rect 8573 9123 8631 9129
rect 2332 9064 2728 9092
rect 1765 9027 1823 9033
rect 1765 8993 1777 9027
rect 1811 9024 1823 9027
rect 2222 9024 2228 9036
rect 1811 8996 2228 9024
rect 1811 8993 1823 8996
rect 1765 8987 1823 8993
rect 2222 8984 2228 8996
rect 2280 8984 2286 9036
rect 2332 9033 2360 9064
rect 2590 9033 2596 9036
rect 2317 9027 2375 9033
rect 2317 8993 2329 9027
rect 2363 8993 2375 9027
rect 2584 9024 2596 9033
rect 2551 8996 2596 9024
rect 2317 8987 2375 8993
rect 2584 8987 2596 8996
rect 2590 8984 2596 8987
rect 2648 8984 2654 9036
rect 2700 9024 2728 9064
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 17310 9092 17316 9104
rect 4120 9064 17316 9092
rect 4120 9052 4126 9064
rect 17310 9052 17316 9064
rect 17368 9052 17374 9104
rect 3142 9024 3148 9036
rect 2700 8996 3148 9024
rect 3142 8984 3148 8996
rect 3200 8984 3206 9036
rect 4525 9027 4583 9033
rect 4525 8993 4537 9027
rect 4571 9024 4583 9027
rect 4982 9024 4988 9036
rect 4571 8996 4988 9024
rect 4571 8993 4583 8996
rect 4525 8987 4583 8993
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 5092 8996 5641 9024
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 5092 8965 5120 8996
rect 5629 8993 5641 8996
rect 5675 9024 5687 9027
rect 7193 9027 7251 9033
rect 7193 9024 7205 9027
rect 5675 8996 7205 9024
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 7193 8993 7205 8996
rect 7239 8993 7251 9027
rect 8018 9024 8024 9036
rect 7979 8996 8024 9024
rect 7193 8987 7251 8993
rect 5077 8959 5135 8965
rect 5077 8956 5089 8959
rect 3936 8928 5089 8956
rect 3936 8916 3942 8928
rect 5077 8925 5089 8928
rect 5123 8925 5135 8959
rect 5077 8919 5135 8925
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8925 5227 8959
rect 5169 8919 5227 8925
rect 5184 8888 5212 8919
rect 3712 8860 5212 8888
rect 7208 8888 7236 8987
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 7708 8928 8125 8956
rect 7708 8916 7714 8928
rect 8113 8925 8125 8928
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 8846 8888 8852 8900
rect 7208 8860 8852 8888
rect 3712 8832 3740 8860
rect 8846 8848 8852 8860
rect 8904 8848 8910 8900
rect 3694 8820 3700 8832
rect 3655 8792 3700 8820
rect 3694 8780 3700 8792
rect 3752 8780 3758 8832
rect 3786 8780 3792 8832
rect 3844 8820 3850 8832
rect 4249 8823 4307 8829
rect 4249 8820 4261 8823
rect 3844 8792 4261 8820
rect 3844 8780 3850 8792
rect 4249 8789 4261 8792
rect 4295 8820 4307 8823
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4295 8792 4537 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 4525 8783 4583 8789
rect 6270 8780 6276 8832
rect 6328 8820 6334 8832
rect 6641 8823 6699 8829
rect 6641 8820 6653 8823
rect 6328 8792 6653 8820
rect 6328 8780 6334 8792
rect 6641 8789 6653 8792
rect 6687 8820 6699 8823
rect 7282 8820 7288 8832
rect 6687 8792 7288 8820
rect 6687 8789 6699 8792
rect 6641 8783 6699 8789
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 7561 8823 7619 8829
rect 7561 8789 7573 8823
rect 7607 8820 7619 8823
rect 8478 8820 8484 8832
rect 7607 8792 8484 8820
rect 7607 8789 7619 8792
rect 7561 8783 7619 8789
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 4890 8616 4896 8628
rect 4851 8588 4896 8616
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5997 8619 6055 8625
rect 5997 8616 6009 8619
rect 5368 8588 6009 8616
rect 4525 8551 4583 8557
rect 4525 8517 4537 8551
rect 4571 8548 4583 8551
rect 4798 8548 4804 8560
rect 4571 8520 4804 8548
rect 4571 8517 4583 8520
rect 4525 8511 4583 8517
rect 4798 8508 4804 8520
rect 4856 8508 4862 8560
rect 2222 8480 2228 8492
rect 2183 8452 2228 8480
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 5368 8489 5396 8588
rect 5997 8585 6009 8588
rect 6043 8616 6055 8619
rect 6043 8588 7880 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 7852 8548 7880 8588
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 8076 8588 8493 8616
rect 8076 8576 8082 8588
rect 8481 8585 8493 8588
rect 8527 8585 8539 8619
rect 8481 8579 8539 8585
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9585 8619 9643 8625
rect 9585 8616 9597 8619
rect 9355 8588 9597 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9585 8585 9597 8588
rect 9631 8616 9643 8619
rect 11882 8616 11888 8628
rect 9631 8588 11888 8616
rect 9631 8585 9643 8588
rect 9585 8579 9643 8585
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 11146 8548 11152 8560
rect 7852 8520 11152 8548
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8449 5503 8483
rect 5445 8443 5503 8449
rect 2041 8415 2099 8421
rect 2041 8381 2053 8415
rect 2087 8412 2099 8415
rect 2958 8412 2964 8424
rect 2087 8384 2964 8412
rect 2087 8381 2099 8384
rect 2041 8375 2099 8381
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 3142 8372 3148 8424
rect 3200 8412 3206 8424
rect 3412 8415 3470 8421
rect 3200 8384 3293 8412
rect 3200 8372 3206 8384
rect 3412 8381 3424 8415
rect 3458 8412 3470 8415
rect 3694 8412 3700 8424
rect 3458 8384 3700 8412
rect 3458 8381 3470 8384
rect 3412 8375 3470 8381
rect 3694 8372 3700 8384
rect 3752 8412 3758 8424
rect 5460 8412 5488 8443
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 9033 8483 9091 8489
rect 9033 8480 9045 8483
rect 8812 8452 9045 8480
rect 8812 8440 8818 8452
rect 9033 8449 9045 8452
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 3752 8384 5488 8412
rect 6825 8415 6883 8421
rect 3752 8372 3758 8384
rect 6825 8381 6837 8415
rect 6871 8412 6883 8415
rect 7374 8412 7380 8424
rect 6871 8384 7380 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 8849 8415 8907 8421
rect 8849 8412 8861 8415
rect 8444 8384 8861 8412
rect 8444 8372 8450 8384
rect 8849 8381 8861 8384
rect 8895 8381 8907 8415
rect 8849 8375 8907 8381
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8412 8999 8415
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 8987 8384 9321 8412
rect 8987 8381 8999 8384
rect 8941 8375 8999 8381
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 3160 8276 3188 8372
rect 5261 8347 5319 8353
rect 5261 8313 5273 8347
rect 5307 8344 5319 8347
rect 5534 8344 5540 8356
rect 5307 8316 5540 8344
rect 5307 8313 5319 8316
rect 5261 8307 5319 8313
rect 5534 8304 5540 8316
rect 5592 8344 5598 8356
rect 7098 8353 7104 8356
rect 6273 8347 6331 8353
rect 6273 8344 6285 8347
rect 5592 8316 6285 8344
rect 5592 8304 5598 8316
rect 6273 8313 6285 8316
rect 6319 8313 6331 8347
rect 7092 8344 7104 8353
rect 7059 8316 7104 8344
rect 6273 8307 6331 8313
rect 7092 8307 7104 8316
rect 7098 8304 7104 8307
rect 7156 8304 7162 8356
rect 7576 8316 8340 8344
rect 3970 8276 3976 8288
rect 3160 8248 3976 8276
rect 3970 8236 3976 8248
rect 4028 8276 4034 8288
rect 5718 8276 5724 8288
rect 4028 8248 5724 8276
rect 4028 8236 4034 8248
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 5810 8236 5816 8288
rect 5868 8276 5874 8288
rect 7576 8276 7604 8316
rect 5868 8248 7604 8276
rect 5868 8236 5874 8248
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 7708 8248 8217 8276
rect 7708 8236 7714 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 8312 8276 8340 8316
rect 17494 8276 17500 8288
rect 8312 8248 17500 8276
rect 8205 8239 8263 8245
rect 17494 8236 17500 8248
rect 17552 8236 17558 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 2958 8072 2964 8084
rect 1688 8044 2728 8072
rect 2919 8044 2964 8072
rect 1688 7936 1716 8044
rect 1762 7964 1768 8016
rect 1820 8004 1826 8016
rect 2225 8007 2283 8013
rect 2225 8004 2237 8007
rect 1820 7976 2237 8004
rect 1820 7964 1826 7976
rect 2225 7973 2237 7976
rect 2271 7973 2283 8007
rect 2700 8004 2728 8044
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 4246 8072 4252 8084
rect 3467 8044 4252 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4430 8032 4436 8084
rect 4488 8072 4494 8084
rect 5810 8072 5816 8084
rect 4488 8044 5816 8072
rect 4488 8032 4494 8044
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 7098 8072 7104 8084
rect 7011 8044 7104 8072
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 8478 8032 8484 8084
rect 8536 8072 8542 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 8536 8044 10149 8072
rect 8536 8032 8542 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 14734 8072 14740 8084
rect 10137 8035 10195 8041
rect 12176 8044 14740 8072
rect 4332 8007 4390 8013
rect 2700 7976 4292 8004
rect 2225 7967 2283 7973
rect 1938 7939 1996 7945
rect 1938 7936 1950 7939
rect 1688 7908 1950 7936
rect 1938 7905 1950 7908
rect 1984 7905 1996 7939
rect 1938 7899 1996 7905
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7936 3387 7939
rect 4154 7936 4160 7948
rect 3375 7908 4160 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 4154 7896 4160 7908
rect 4212 7896 4218 7948
rect 4264 7936 4292 7976
rect 4332 7973 4344 8007
rect 4378 8004 4390 8007
rect 4798 8004 4804 8016
rect 4378 7976 4804 8004
rect 4378 7973 4390 7976
rect 4332 7967 4390 7973
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 7116 8004 7144 8032
rect 8754 8004 8760 8016
rect 4908 7976 6776 8004
rect 7116 7976 8760 8004
rect 4908 7936 4936 7976
rect 5977 7939 6035 7945
rect 5977 7936 5989 7939
rect 4264 7908 4936 7936
rect 5460 7908 5989 7936
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 3605 7831 3663 7837
rect 3620 7732 3648 7831
rect 3970 7828 3976 7880
rect 4028 7868 4034 7880
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 4028 7840 4077 7868
rect 4028 7828 4034 7840
rect 4065 7837 4077 7840
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 5460 7741 5488 7908
rect 5977 7905 5989 7908
rect 6023 7905 6035 7939
rect 5977 7899 6035 7905
rect 5718 7868 5724 7880
rect 5679 7840 5724 7868
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 5445 7735 5503 7741
rect 5445 7732 5457 7735
rect 3620 7704 5457 7732
rect 5445 7701 5457 7704
rect 5491 7701 5503 7735
rect 6748 7732 6776 7976
rect 8754 7964 8760 7976
rect 8812 7964 8818 8016
rect 8846 7964 8852 8016
rect 8904 8004 8910 8016
rect 12176 8004 12204 8044
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 8904 7976 12204 8004
rect 8904 7964 8910 7976
rect 7374 7936 7380 7948
rect 7335 7908 7380 7936
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 7650 7945 7656 7948
rect 7644 7936 7656 7945
rect 7611 7908 7656 7936
rect 7644 7899 7656 7908
rect 7650 7896 7656 7899
rect 7708 7896 7714 7948
rect 8478 7896 8484 7948
rect 8536 7936 8542 7948
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 8536 7908 10057 7936
rect 8536 7896 8542 7908
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 10045 7899 10103 7905
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 8662 7760 8668 7812
rect 8720 7800 8726 7812
rect 8757 7803 8815 7809
rect 8757 7800 8769 7803
rect 8720 7772 8769 7800
rect 8720 7760 8726 7772
rect 8757 7769 8769 7772
rect 8803 7800 8815 7803
rect 10244 7800 10272 7831
rect 8803 7772 10272 7800
rect 8803 7769 8815 7772
rect 8757 7763 8815 7769
rect 9677 7735 9735 7741
rect 9677 7732 9689 7735
rect 6748 7704 9689 7732
rect 5445 7695 5503 7701
rect 9677 7701 9689 7704
rect 9723 7701 9735 7735
rect 9677 7695 9735 7701
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 4154 7528 4160 7540
rect 4115 7500 4160 7528
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 8113 7531 8171 7537
rect 8113 7497 8125 7531
rect 8159 7528 8171 7531
rect 8202 7528 8208 7540
rect 8159 7500 8208 7528
rect 8159 7497 8171 7500
rect 8113 7491 8171 7497
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 19429 7531 19487 7537
rect 19429 7497 19441 7531
rect 19475 7528 19487 7531
rect 19702 7528 19708 7540
rect 19475 7500 19708 7528
rect 19475 7497 19487 7500
rect 19429 7491 19487 7497
rect 19702 7488 19708 7500
rect 19760 7488 19766 7540
rect 7098 7420 7104 7472
rect 7156 7460 7162 7472
rect 18877 7463 18935 7469
rect 7156 7432 7201 7460
rect 7156 7420 7162 7432
rect 18877 7429 18889 7463
rect 18923 7460 18935 7463
rect 19518 7460 19524 7472
rect 18923 7432 19524 7460
rect 18923 7429 18935 7432
rect 18877 7423 18935 7429
rect 19518 7420 19524 7432
rect 19576 7420 19582 7472
rect 4706 7392 4712 7404
rect 4667 7364 4712 7392
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 7745 7395 7803 7401
rect 6512 7364 7687 7392
rect 6512 7352 6518 7364
rect 4525 7259 4583 7265
rect 4525 7225 4537 7259
rect 4571 7256 4583 7259
rect 5169 7259 5227 7265
rect 5169 7256 5181 7259
rect 4571 7228 5181 7256
rect 4571 7225 4583 7228
rect 4525 7219 4583 7225
rect 5169 7225 5181 7228
rect 5215 7225 5227 7259
rect 5169 7219 5227 7225
rect 6730 7216 6736 7268
rect 6788 7256 6794 7268
rect 7469 7259 7527 7265
rect 7469 7256 7481 7259
rect 6788 7228 7481 7256
rect 6788 7216 6794 7228
rect 7469 7225 7481 7228
rect 7515 7225 7527 7259
rect 7659 7256 7687 7364
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 8754 7392 8760 7404
rect 7791 7364 8760 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 7834 7284 7840 7336
rect 7892 7324 7898 7336
rect 18325 7327 18383 7333
rect 18325 7324 18337 7327
rect 7892 7296 18337 7324
rect 7892 7284 7898 7296
rect 18325 7293 18337 7296
rect 18371 7324 18383 7327
rect 18693 7327 18751 7333
rect 18693 7324 18705 7327
rect 18371 7296 18705 7324
rect 18371 7293 18383 7296
rect 18325 7287 18383 7293
rect 18693 7293 18705 7296
rect 18739 7293 18751 7327
rect 18693 7287 18751 7293
rect 18782 7284 18788 7336
rect 18840 7324 18846 7336
rect 19245 7327 19303 7333
rect 19245 7324 19257 7327
rect 18840 7296 19257 7324
rect 18840 7284 18846 7296
rect 19245 7293 19257 7296
rect 19291 7324 19303 7327
rect 19797 7327 19855 7333
rect 19797 7324 19809 7327
rect 19291 7296 19809 7324
rect 19291 7293 19303 7296
rect 19245 7287 19303 7293
rect 19797 7293 19809 7296
rect 19843 7293 19855 7327
rect 19797 7287 19855 7293
rect 8573 7259 8631 7265
rect 8573 7256 8585 7259
rect 7659 7228 8585 7256
rect 7469 7219 7527 7225
rect 8573 7225 8585 7228
rect 8619 7256 8631 7259
rect 9125 7259 9183 7265
rect 9125 7256 9137 7259
rect 8619 7228 9137 7256
rect 8619 7225 8631 7228
rect 8573 7219 8631 7225
rect 9125 7225 9137 7228
rect 9171 7225 9183 7259
rect 9125 7219 9183 7225
rect 3786 7188 3792 7200
rect 3747 7160 3792 7188
rect 3786 7148 3792 7160
rect 3844 7188 3850 7200
rect 4617 7191 4675 7197
rect 4617 7188 4629 7191
rect 3844 7160 4629 7188
rect 3844 7148 3850 7160
rect 4617 7157 4629 7160
rect 4663 7188 4675 7191
rect 6270 7188 6276 7200
rect 4663 7160 6276 7188
rect 4663 7157 4675 7160
rect 4617 7151 4675 7157
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 6362 7148 6368 7200
rect 6420 7188 6426 7200
rect 7561 7191 7619 7197
rect 7561 7188 7573 7191
rect 6420 7160 7573 7188
rect 6420 7148 6426 7160
rect 7561 7157 7573 7160
rect 7607 7157 7619 7191
rect 7561 7151 7619 7157
rect 7742 7148 7748 7200
rect 7800 7188 7806 7200
rect 8481 7191 8539 7197
rect 8481 7188 8493 7191
rect 7800 7160 8493 7188
rect 7800 7148 7806 7160
rect 8481 7157 8493 7160
rect 8527 7188 8539 7191
rect 9493 7191 9551 7197
rect 9493 7188 9505 7191
rect 8527 7160 9505 7188
rect 8527 7157 8539 7160
rect 8481 7151 8539 7157
rect 9493 7157 9505 7160
rect 9539 7157 9551 7191
rect 9493 7151 9551 7157
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 2774 6944 2780 6996
rect 2832 6984 2838 6996
rect 6362 6984 6368 6996
rect 2832 6956 6368 6984
rect 2832 6944 2838 6956
rect 6362 6944 6368 6956
rect 6420 6944 6426 6996
rect 7098 6944 7104 6996
rect 7156 6984 7162 6996
rect 7653 6987 7711 6993
rect 7653 6984 7665 6987
rect 7156 6956 7665 6984
rect 7156 6944 7162 6956
rect 7653 6953 7665 6956
rect 7699 6953 7711 6987
rect 7653 6947 7711 6953
rect 7484 6888 8340 6916
rect 3970 6808 3976 6860
rect 4028 6848 4034 6860
rect 7484 6848 7512 6888
rect 4028 6820 7512 6848
rect 7561 6851 7619 6857
rect 4028 6808 4034 6820
rect 7561 6817 7573 6851
rect 7607 6848 7619 6851
rect 8205 6851 8263 6857
rect 8205 6848 8217 6851
rect 7607 6820 8217 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 8205 6817 8217 6820
rect 8251 6817 8263 6851
rect 8312 6848 8340 6888
rect 19613 6851 19671 6857
rect 19613 6848 19625 6851
rect 8312 6820 19625 6848
rect 8205 6811 8263 6817
rect 19613 6817 19625 6820
rect 19659 6848 19671 6851
rect 20165 6851 20223 6857
rect 20165 6848 20177 6851
rect 19659 6820 20177 6848
rect 19659 6817 19671 6820
rect 19613 6811 19671 6817
rect 20165 6817 20177 6820
rect 20211 6817 20223 6851
rect 20165 6811 20223 6817
rect 5626 6740 5632 6792
rect 5684 6780 5690 6792
rect 6730 6780 6736 6792
rect 5684 6752 6736 6780
rect 5684 6740 5690 6752
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 7708 6752 7757 6780
rect 7708 6740 7714 6752
rect 7745 6749 7757 6752
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 19797 6715 19855 6721
rect 19797 6681 19809 6715
rect 19843 6712 19855 6715
rect 20438 6712 20444 6724
rect 19843 6684 20444 6712
rect 19843 6681 19855 6684
rect 19797 6675 19855 6681
rect 20438 6672 20444 6684
rect 20496 6672 20502 6724
rect 7193 6647 7251 6653
rect 7193 6613 7205 6647
rect 7239 6644 7251 6647
rect 8478 6644 8484 6656
rect 7239 6616 8484 6644
rect 7239 6613 7251 6616
rect 7193 6607 7251 6613
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 18782 6644 18788 6656
rect 8628 6616 18788 6644
rect 8628 6604 8634 6616
rect 18782 6604 18788 6616
rect 18840 6604 18846 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 20165 6443 20223 6449
rect 20165 6409 20177 6443
rect 20211 6440 20223 6443
rect 20898 6440 20904 6452
rect 20211 6412 20904 6440
rect 20211 6409 20223 6412
rect 20165 6403 20223 6409
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 19981 6239 20039 6245
rect 19981 6205 19993 6239
rect 20027 6205 20039 6239
rect 19981 6199 20039 6205
rect 19996 6168 20024 6199
rect 20533 6171 20591 6177
rect 20533 6168 20545 6171
rect 19996 6140 20545 6168
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 19996 6100 20024 6140
rect 20533 6137 20545 6140
rect 20579 6137 20591 6171
rect 20533 6131 20591 6137
rect 4120 6072 20024 6100
rect 4120 6060 4126 6072
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 21082 5896 21088 5908
rect 21043 5868 21088 5896
rect 21082 5856 21088 5868
rect 21140 5856 21146 5908
rect 20438 5720 20444 5772
rect 20496 5760 20502 5772
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20496 5732 20913 5760
rect 20496 5720 20502 5732
rect 20901 5729 20913 5732
rect 20947 5729 20959 5763
rect 20901 5723 20959 5729
rect 20438 5556 20444 5568
rect 20399 5528 20444 5556
rect 20438 5516 20444 5528
rect 20496 5516 20502 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 20438 5352 20444 5364
rect 4120 5324 20444 5352
rect 4120 5312 4126 5324
rect 20438 5312 20444 5324
rect 20496 5312 20502 5364
rect 20990 5352 20996 5364
rect 20951 5324 20996 5352
rect 20990 5312 20996 5324
rect 21048 5312 21054 5364
rect 3970 5244 3976 5296
rect 4028 5284 4034 5296
rect 14642 5284 14648 5296
rect 4028 5256 14648 5284
rect 4028 5244 4034 5256
rect 14642 5244 14648 5256
rect 14700 5244 14706 5296
rect 20809 5151 20867 5157
rect 20809 5148 20821 5151
rect 20456 5120 20821 5148
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 20456 5021 20484 5120
rect 20809 5117 20821 5120
rect 20855 5117 20867 5151
rect 20809 5111 20867 5117
rect 20441 5015 20499 5021
rect 20441 5012 20453 5015
rect 4120 4984 20453 5012
rect 4120 4972 4126 4984
rect 20441 4981 20453 4984
rect 20487 4981 20499 5015
rect 20441 4975 20499 4981
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 11698 4768 11704 4820
rect 11756 4808 11762 4820
rect 12066 4808 12072 4820
rect 11756 4780 12072 4808
rect 11756 4768 11762 4780
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 3510 2048 3516 2100
rect 3568 2088 3574 2100
rect 6822 2088 6828 2100
rect 3568 2060 6828 2088
rect 3568 2048 3574 2060
rect 6822 2048 6828 2060
rect 6880 2048 6886 2100
rect 3326 1300 3332 1352
rect 3384 1340 3390 1352
rect 5534 1340 5540 1352
rect 3384 1312 5540 1340
rect 3384 1300 3390 1312
rect 5534 1300 5540 1312
rect 5592 1300 5598 1352
<< via1 >>
rect 2964 21904 3016 21956
rect 3976 21904 4028 21956
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 1952 20587 2004 20596
rect 1952 20553 1961 20587
rect 1961 20553 1995 20587
rect 1995 20553 2004 20587
rect 1952 20544 2004 20553
rect 2780 20544 2832 20596
rect 8944 20544 8996 20596
rect 14924 20544 14976 20596
rect 8760 20451 8812 20460
rect 8760 20417 8769 20451
rect 8769 20417 8803 20451
rect 8803 20417 8812 20451
rect 8760 20408 8812 20417
rect 1768 20383 1820 20392
rect 1768 20349 1777 20383
rect 1777 20349 1811 20383
rect 1811 20349 1820 20383
rect 1768 20340 1820 20349
rect 1860 20340 1912 20392
rect 12808 20383 12860 20392
rect 12808 20349 12817 20383
rect 12817 20349 12851 20383
rect 12851 20349 12860 20383
rect 12808 20340 12860 20349
rect 14096 20383 14148 20392
rect 14096 20349 14105 20383
rect 14105 20349 14139 20383
rect 14139 20349 14148 20383
rect 14096 20340 14148 20349
rect 4160 20272 4212 20324
rect 14556 20272 14608 20324
rect 3148 20247 3200 20256
rect 3148 20213 3157 20247
rect 3157 20213 3191 20247
rect 3191 20213 3200 20247
rect 3148 20204 3200 20213
rect 4896 20247 4948 20256
rect 4896 20213 4905 20247
rect 4905 20213 4939 20247
rect 4939 20213 4948 20247
rect 4896 20204 4948 20213
rect 8208 20204 8260 20256
rect 11060 20204 11112 20256
rect 12164 20204 12216 20256
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 4160 20043 4212 20052
rect 4160 20009 4169 20043
rect 4169 20009 4203 20043
rect 4203 20009 4212 20043
rect 4160 20000 4212 20009
rect 4896 20043 4948 20052
rect 4896 20009 4905 20043
rect 4905 20009 4939 20043
rect 4939 20009 4948 20043
rect 4896 20000 4948 20009
rect 9404 20000 9456 20052
rect 2872 19932 2924 19984
rect 8760 19932 8812 19984
rect 13544 20000 13596 20052
rect 14464 20000 14516 20052
rect 15384 20000 15436 20052
rect 15844 20000 15896 20052
rect 16304 20000 16356 20052
rect 16764 20000 16816 20052
rect 18604 20000 18656 20052
rect 1860 19907 1912 19916
rect 1860 19873 1869 19907
rect 1869 19873 1903 19907
rect 1903 19873 1912 19907
rect 1860 19864 1912 19873
rect 4344 19864 4396 19916
rect 5724 19864 5776 19916
rect 6460 19864 6512 19916
rect 8300 19864 8352 19916
rect 9772 19864 9824 19916
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 14556 19907 14608 19916
rect 2688 19660 2740 19712
rect 3700 19703 3752 19712
rect 3700 19669 3709 19703
rect 3709 19669 3743 19703
rect 3743 19669 3752 19703
rect 3700 19660 3752 19669
rect 4160 19660 4212 19712
rect 4804 19660 4856 19712
rect 5448 19796 5500 19848
rect 10140 19839 10192 19848
rect 10140 19805 10149 19839
rect 10149 19805 10183 19839
rect 10183 19805 10192 19839
rect 10140 19796 10192 19805
rect 14556 19873 14565 19907
rect 14565 19873 14599 19907
rect 14599 19873 14608 19907
rect 14556 19864 14608 19873
rect 14648 19864 14700 19916
rect 15384 19864 15436 19916
rect 16396 19907 16448 19916
rect 16396 19873 16405 19907
rect 16405 19873 16439 19907
rect 16439 19873 16448 19907
rect 16396 19864 16448 19873
rect 16948 19907 17000 19916
rect 16948 19873 16957 19907
rect 16957 19873 16991 19907
rect 16991 19873 17000 19907
rect 16948 19864 17000 19873
rect 18880 19932 18932 19984
rect 18144 19864 18196 19916
rect 14188 19796 14240 19848
rect 10048 19728 10100 19780
rect 14004 19728 14056 19780
rect 17684 19728 17736 19780
rect 8300 19703 8352 19712
rect 8300 19669 8309 19703
rect 8309 19669 8343 19703
rect 8343 19669 8352 19703
rect 8300 19660 8352 19669
rect 9036 19660 9088 19712
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 1768 19320 1820 19372
rect 1400 19295 1452 19304
rect 1400 19261 1409 19295
rect 1409 19261 1443 19295
rect 1443 19261 1452 19295
rect 1400 19252 1452 19261
rect 2688 19252 2740 19304
rect 4344 19456 4396 19508
rect 5448 19456 5500 19508
rect 6460 19499 6512 19508
rect 6460 19465 6469 19499
rect 6469 19465 6503 19499
rect 6503 19465 6512 19499
rect 6460 19456 6512 19465
rect 4068 19320 4120 19372
rect 4988 19320 5040 19372
rect 9680 19320 9732 19372
rect 10140 19456 10192 19508
rect 14096 19388 14148 19440
rect 16396 19320 16448 19372
rect 16948 19320 17000 19372
rect 4160 19252 4212 19304
rect 4804 19252 4856 19304
rect 5080 19295 5132 19304
rect 5080 19261 5089 19295
rect 5089 19261 5123 19295
rect 5123 19261 5132 19295
rect 5080 19252 5132 19261
rect 7380 19295 7432 19304
rect 7380 19261 7389 19295
rect 7389 19261 7423 19295
rect 7423 19261 7432 19295
rect 7380 19252 7432 19261
rect 8760 19252 8812 19304
rect 11244 19252 11296 19304
rect 12624 19252 12676 19304
rect 13360 19295 13412 19304
rect 13360 19261 13369 19295
rect 13369 19261 13403 19295
rect 13403 19261 13412 19295
rect 13360 19252 13412 19261
rect 14740 19295 14792 19304
rect 14740 19261 14749 19295
rect 14749 19261 14783 19295
rect 14783 19261 14792 19295
rect 14740 19252 14792 19261
rect 15384 19252 15436 19304
rect 16304 19295 16356 19304
rect 6092 19184 6144 19236
rect 10048 19227 10100 19236
rect 10048 19193 10082 19227
rect 10082 19193 10100 19227
rect 10048 19184 10100 19193
rect 14648 19184 14700 19236
rect 16304 19261 16313 19295
rect 16313 19261 16347 19295
rect 16347 19261 16356 19295
rect 16304 19252 16356 19261
rect 17040 19295 17092 19304
rect 17040 19261 17049 19295
rect 17049 19261 17083 19295
rect 17083 19261 17092 19295
rect 17040 19252 17092 19261
rect 17960 19252 18012 19304
rect 20720 19252 20772 19304
rect 16580 19184 16632 19236
rect 18236 19184 18288 19236
rect 21180 19227 21232 19236
rect 21180 19193 21189 19227
rect 21189 19193 21223 19227
rect 21223 19193 21232 19227
rect 21180 19184 21232 19193
rect 1676 19116 1728 19168
rect 2596 19116 2648 19168
rect 4528 19116 4580 19168
rect 5264 19116 5316 19168
rect 6736 19116 6788 19168
rect 7748 19116 7800 19168
rect 8944 19116 8996 19168
rect 9772 19116 9824 19168
rect 13084 19116 13136 19168
rect 18052 19116 18104 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 2872 18955 2924 18964
rect 2872 18921 2881 18955
rect 2881 18921 2915 18955
rect 2915 18921 2924 18955
rect 2872 18912 2924 18921
rect 3148 18912 3200 18964
rect 4988 18912 5040 18964
rect 5724 18912 5776 18964
rect 6736 18912 6788 18964
rect 1400 18844 1452 18896
rect 3424 18844 3476 18896
rect 4528 18819 4580 18828
rect 4528 18785 4537 18819
rect 4537 18785 4571 18819
rect 4571 18785 4580 18819
rect 4528 18776 4580 18785
rect 5172 18776 5224 18828
rect 5816 18844 5868 18896
rect 7288 18844 7340 18896
rect 8208 18912 8260 18964
rect 8944 18955 8996 18964
rect 8944 18921 8953 18955
rect 8953 18921 8987 18955
rect 8987 18921 8996 18955
rect 8944 18912 8996 18921
rect 9036 18955 9088 18964
rect 9036 18921 9045 18955
rect 9045 18921 9079 18955
rect 9079 18921 9088 18955
rect 9036 18912 9088 18921
rect 10048 18912 10100 18964
rect 14648 18912 14700 18964
rect 17132 18912 17184 18964
rect 17224 18912 17276 18964
rect 19064 18912 19116 18964
rect 20720 18912 20772 18964
rect 22284 18912 22336 18964
rect 8300 18844 8352 18896
rect 7840 18819 7892 18828
rect 3700 18708 3752 18760
rect 4344 18708 4396 18760
rect 5540 18751 5592 18760
rect 5540 18717 5549 18751
rect 5549 18717 5583 18751
rect 5583 18717 5592 18751
rect 5540 18708 5592 18717
rect 6092 18708 6144 18760
rect 6460 18640 6512 18692
rect 7840 18785 7849 18819
rect 7849 18785 7883 18819
rect 7883 18785 7892 18819
rect 7840 18776 7892 18785
rect 7932 18776 7984 18828
rect 10508 18844 10560 18896
rect 14280 18844 14332 18896
rect 7748 18708 7800 18760
rect 9772 18776 9824 18828
rect 9956 18819 10008 18828
rect 9956 18785 9990 18819
rect 9990 18785 10008 18819
rect 9956 18776 10008 18785
rect 12532 18776 12584 18828
rect 13544 18819 13596 18828
rect 13544 18785 13553 18819
rect 13553 18785 13587 18819
rect 13587 18785 13596 18819
rect 13544 18776 13596 18785
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 12900 18708 12952 18760
rect 14648 18751 14700 18760
rect 14188 18683 14240 18692
rect 2044 18572 2096 18624
rect 7932 18572 7984 18624
rect 8300 18572 8352 18624
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 14188 18649 14197 18683
rect 14197 18649 14231 18683
rect 14231 18649 14240 18683
rect 14188 18640 14240 18649
rect 14648 18717 14657 18751
rect 14657 18717 14691 18751
rect 14691 18717 14700 18751
rect 14648 18708 14700 18717
rect 16948 18776 17000 18828
rect 18236 18819 18288 18828
rect 18236 18785 18245 18819
rect 18245 18785 18279 18819
rect 18279 18785 18288 18819
rect 18236 18776 18288 18785
rect 15752 18751 15804 18760
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 16764 18751 16816 18760
rect 15384 18640 15436 18692
rect 16764 18717 16773 18751
rect 16773 18717 16807 18751
rect 16807 18717 16816 18751
rect 16764 18708 16816 18717
rect 16672 18640 16724 18692
rect 14556 18572 14608 18624
rect 15292 18615 15344 18624
rect 15292 18581 15301 18615
rect 15301 18581 15335 18615
rect 15335 18581 15344 18615
rect 15292 18572 15344 18581
rect 15476 18572 15528 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 1860 18164 1912 18216
rect 4160 18368 4212 18420
rect 12440 18368 12492 18420
rect 13636 18368 13688 18420
rect 14280 18411 14332 18420
rect 14280 18377 14289 18411
rect 14289 18377 14323 18411
rect 14323 18377 14332 18411
rect 14280 18368 14332 18377
rect 14648 18368 14700 18420
rect 15384 18368 15436 18420
rect 2688 18232 2740 18284
rect 6092 18300 6144 18352
rect 6552 18300 6604 18352
rect 664 18096 716 18148
rect 5080 18207 5132 18216
rect 3700 18096 3752 18148
rect 3884 18096 3936 18148
rect 4804 18096 4856 18148
rect 5080 18173 5089 18207
rect 5089 18173 5123 18207
rect 5123 18173 5132 18207
rect 5080 18164 5132 18173
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 10416 18300 10468 18352
rect 12900 18300 12952 18352
rect 8668 18232 8720 18284
rect 12348 18232 12400 18284
rect 7288 18164 7340 18216
rect 8300 18207 8352 18216
rect 8300 18173 8309 18207
rect 8309 18173 8343 18207
rect 8343 18173 8352 18207
rect 8300 18164 8352 18173
rect 8392 18164 8444 18216
rect 12072 18164 12124 18216
rect 12256 18164 12308 18216
rect 12532 18164 12584 18216
rect 15292 18275 15344 18284
rect 15292 18241 15301 18275
rect 15301 18241 15335 18275
rect 15335 18241 15344 18275
rect 15292 18232 15344 18241
rect 18144 18232 18196 18284
rect 15476 18164 15528 18216
rect 18052 18207 18104 18216
rect 5172 18096 5224 18148
rect 6184 18096 6236 18148
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 2504 18071 2556 18080
rect 2504 18037 2513 18071
rect 2513 18037 2547 18071
rect 2547 18037 2556 18071
rect 2504 18028 2556 18037
rect 2596 18028 2648 18080
rect 7012 18028 7064 18080
rect 7564 18028 7616 18080
rect 7932 18096 7984 18148
rect 15292 18096 15344 18148
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 18052 18164 18104 18173
rect 19248 18164 19300 18216
rect 22744 18164 22796 18216
rect 16672 18096 16724 18148
rect 8392 18028 8444 18080
rect 10876 18028 10928 18080
rect 21180 18096 21232 18148
rect 17224 18028 17276 18080
rect 20996 18028 21048 18080
rect 21824 18028 21876 18080
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 1768 17867 1820 17876
rect 1768 17833 1777 17867
rect 1777 17833 1811 17867
rect 1811 17833 1820 17867
rect 1768 17824 1820 17833
rect 2964 17824 3016 17876
rect 4896 17824 4948 17876
rect 5540 17824 5592 17876
rect 6276 17824 6328 17876
rect 2044 17756 2096 17808
rect 11980 17824 12032 17876
rect 12440 17824 12492 17876
rect 12900 17824 12952 17876
rect 13544 17867 13596 17876
rect 10048 17756 10100 17808
rect 10140 17756 10192 17808
rect 11888 17756 11940 17808
rect 12348 17799 12400 17808
rect 12348 17765 12357 17799
rect 12357 17765 12391 17799
rect 12391 17765 12400 17799
rect 12348 17756 12400 17765
rect 12532 17756 12584 17808
rect 13544 17833 13553 17867
rect 13553 17833 13587 17867
rect 13587 17833 13596 17867
rect 13544 17824 13596 17833
rect 14556 17867 14608 17876
rect 14556 17833 14565 17867
rect 14565 17833 14599 17867
rect 14599 17833 14608 17867
rect 14556 17824 14608 17833
rect 16672 17867 16724 17876
rect 16672 17833 16681 17867
rect 16681 17833 16715 17867
rect 16715 17833 16724 17867
rect 16672 17824 16724 17833
rect 18052 17824 18104 17876
rect 15752 17756 15804 17808
rect 1584 17731 1636 17740
rect 1584 17697 1593 17731
rect 1593 17697 1627 17731
rect 1627 17697 1636 17731
rect 1584 17688 1636 17697
rect 2136 17731 2188 17740
rect 2136 17697 2145 17731
rect 2145 17697 2179 17731
rect 2179 17697 2188 17731
rect 2136 17688 2188 17697
rect 3424 17484 3476 17536
rect 6000 17731 6052 17740
rect 6000 17697 6009 17731
rect 6009 17697 6043 17731
rect 6043 17697 6052 17731
rect 6000 17688 6052 17697
rect 8300 17731 8352 17740
rect 8300 17697 8309 17731
rect 8309 17697 8343 17731
rect 8343 17697 8352 17731
rect 8300 17688 8352 17697
rect 8944 17731 8996 17740
rect 8944 17697 8953 17731
rect 8953 17697 8987 17731
rect 8987 17697 8996 17731
rect 8944 17688 8996 17697
rect 9680 17731 9732 17740
rect 4160 17620 4212 17672
rect 6184 17663 6236 17672
rect 6184 17629 6193 17663
rect 6193 17629 6227 17663
rect 6227 17629 6236 17663
rect 7196 17663 7248 17672
rect 6184 17620 6236 17629
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 9036 17663 9088 17672
rect 9036 17629 9045 17663
rect 9045 17629 9079 17663
rect 9079 17629 9088 17663
rect 9036 17620 9088 17629
rect 3976 17552 4028 17604
rect 4068 17527 4120 17536
rect 4068 17493 4077 17527
rect 4077 17493 4111 17527
rect 4111 17493 4120 17527
rect 4068 17484 4120 17493
rect 7380 17552 7432 17604
rect 8668 17552 8720 17604
rect 9680 17697 9689 17731
rect 9689 17697 9723 17731
rect 9723 17697 9732 17731
rect 9680 17688 9732 17697
rect 11704 17731 11756 17740
rect 11704 17697 11713 17731
rect 11713 17697 11747 17731
rect 11747 17697 11756 17731
rect 11704 17688 11756 17697
rect 15108 17688 15160 17740
rect 11796 17663 11848 17672
rect 9312 17484 9364 17536
rect 11796 17629 11805 17663
rect 11805 17629 11839 17663
rect 11839 17629 11848 17663
rect 11796 17620 11848 17629
rect 12440 17620 12492 17672
rect 15292 17663 15344 17672
rect 15292 17629 15301 17663
rect 15301 17629 15335 17663
rect 15335 17629 15344 17663
rect 15292 17620 15344 17629
rect 18052 17620 18104 17672
rect 18788 17663 18840 17672
rect 18788 17629 18797 17663
rect 18797 17629 18831 17663
rect 18831 17629 18840 17663
rect 18788 17620 18840 17629
rect 9956 17484 10008 17536
rect 13176 17484 13228 17536
rect 14280 17484 14332 17536
rect 16672 17484 16724 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 1584 17212 1636 17264
rect 5080 17280 5132 17332
rect 4804 17212 4856 17264
rect 6920 17144 6972 17196
rect 7380 17280 7432 17332
rect 8484 17280 8536 17332
rect 9036 17280 9088 17332
rect 11796 17280 11848 17332
rect 11980 17280 12032 17332
rect 12256 17280 12308 17332
rect 8944 17212 8996 17264
rect 10048 17144 10100 17196
rect 2044 17119 2096 17128
rect 2044 17085 2053 17119
rect 2053 17085 2087 17119
rect 2087 17085 2096 17119
rect 2044 17076 2096 17085
rect 3148 17076 3200 17128
rect 4160 17076 4212 17128
rect 7748 17076 7800 17128
rect 1676 16983 1728 16992
rect 1676 16949 1685 16983
rect 1685 16949 1719 16983
rect 1719 16949 1728 16983
rect 1676 16940 1728 16949
rect 4160 16940 4212 16992
rect 6000 16940 6052 16992
rect 8852 17076 8904 17128
rect 9864 17076 9916 17128
rect 11888 17076 11940 17128
rect 12256 17144 12308 17196
rect 12348 17076 12400 17128
rect 12532 17144 12584 17196
rect 12716 17144 12768 17196
rect 17040 17280 17092 17332
rect 13728 17144 13780 17196
rect 17776 17144 17828 17196
rect 12532 17008 12584 17060
rect 14096 17076 14148 17128
rect 18144 17119 18196 17128
rect 18144 17085 18153 17119
rect 18153 17085 18187 17119
rect 18187 17085 18196 17119
rect 18144 17076 18196 17085
rect 14004 17008 14056 17060
rect 14648 17008 14700 17060
rect 15108 17008 15160 17060
rect 18604 17008 18656 17060
rect 8208 16940 8260 16992
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 9496 16940 9548 16949
rect 13176 16940 13228 16992
rect 14188 16940 14240 16992
rect 17316 16983 17368 16992
rect 17316 16949 17325 16983
rect 17325 16949 17359 16983
rect 17359 16949 17368 16983
rect 17316 16940 17368 16949
rect 17408 16983 17460 16992
rect 17408 16949 17417 16983
rect 17417 16949 17451 16983
rect 17451 16949 17460 16983
rect 17408 16940 17460 16949
rect 18788 16940 18840 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 2136 16736 2188 16788
rect 4068 16736 4120 16788
rect 6184 16736 6236 16788
rect 7196 16736 7248 16788
rect 9312 16736 9364 16788
rect 10232 16779 10284 16788
rect 10232 16745 10241 16779
rect 10241 16745 10275 16779
rect 10275 16745 10284 16779
rect 10232 16736 10284 16745
rect 11152 16736 11204 16788
rect 12348 16779 12400 16788
rect 12348 16745 12357 16779
rect 12357 16745 12391 16779
rect 12391 16745 12400 16779
rect 12348 16736 12400 16745
rect 13360 16736 13412 16788
rect 14004 16736 14056 16788
rect 17776 16779 17828 16788
rect 17776 16745 17785 16779
rect 17785 16745 17819 16779
rect 17819 16745 17828 16779
rect 17776 16736 17828 16745
rect 18604 16736 18656 16788
rect 3056 16668 3108 16720
rect 3148 16668 3200 16720
rect 2228 16600 2280 16652
rect 5448 16600 5500 16652
rect 6920 16643 6972 16652
rect 6920 16609 6929 16643
rect 6929 16609 6963 16643
rect 6963 16609 6972 16643
rect 6920 16600 6972 16609
rect 8208 16600 8260 16652
rect 12716 16668 12768 16720
rect 13912 16668 13964 16720
rect 16764 16668 16816 16720
rect 4160 16532 4212 16584
rect 4804 16532 4856 16584
rect 8852 16600 8904 16652
rect 9496 16600 9548 16652
rect 10600 16643 10652 16652
rect 10600 16609 10609 16643
rect 10609 16609 10643 16643
rect 10643 16609 10652 16643
rect 10600 16600 10652 16609
rect 10968 16643 11020 16652
rect 10968 16609 10977 16643
rect 10977 16609 11011 16643
rect 11011 16609 11020 16643
rect 10968 16600 11020 16609
rect 11980 16600 12032 16652
rect 14004 16600 14056 16652
rect 14280 16643 14332 16652
rect 14280 16609 14289 16643
rect 14289 16609 14323 16643
rect 14323 16609 14332 16643
rect 14280 16600 14332 16609
rect 15292 16600 15344 16652
rect 18144 16600 18196 16652
rect 9036 16575 9088 16584
rect 9036 16541 9045 16575
rect 9045 16541 9079 16575
rect 9079 16541 9088 16575
rect 9036 16532 9088 16541
rect 14188 16532 14240 16584
rect 15200 16532 15252 16584
rect 16028 16532 16080 16584
rect 8392 16396 8444 16448
rect 14556 16396 14608 16448
rect 15660 16439 15712 16448
rect 15660 16405 15669 16439
rect 15669 16405 15703 16439
rect 15703 16405 15712 16439
rect 15660 16396 15712 16405
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 1676 16235 1728 16244
rect 1676 16201 1685 16235
rect 1685 16201 1719 16235
rect 1719 16201 1728 16235
rect 1676 16192 1728 16201
rect 9036 16192 9088 16244
rect 10048 16235 10100 16244
rect 10048 16201 10057 16235
rect 10057 16201 10091 16235
rect 10091 16201 10100 16235
rect 10048 16192 10100 16201
rect 11704 16192 11756 16244
rect 12532 16192 12584 16244
rect 14648 16192 14700 16244
rect 18052 16235 18104 16244
rect 18052 16201 18061 16235
rect 18061 16201 18095 16235
rect 18095 16201 18104 16235
rect 18052 16192 18104 16201
rect 1584 15988 1636 16040
rect 10232 16124 10284 16176
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 5448 16099 5500 16108
rect 5448 16065 5457 16099
rect 5457 16065 5491 16099
rect 5491 16065 5500 16099
rect 5448 16056 5500 16065
rect 8208 16056 8260 16108
rect 8668 16099 8720 16108
rect 8668 16065 8677 16099
rect 8677 16065 8711 16099
rect 8711 16065 8720 16099
rect 8668 16056 8720 16065
rect 11152 16056 11204 16108
rect 3424 15988 3476 16040
rect 8300 15988 8352 16040
rect 9220 15988 9272 16040
rect 12716 16056 12768 16108
rect 8484 15920 8536 15972
rect 9404 15920 9456 15972
rect 10600 15920 10652 15972
rect 18144 16124 18196 16176
rect 13636 16031 13688 16040
rect 13636 15997 13645 16031
rect 13645 15997 13679 16031
rect 13679 15997 13688 16031
rect 13636 15988 13688 15997
rect 15660 16056 15712 16108
rect 16028 16056 16080 16108
rect 17316 16056 17368 16108
rect 18604 16099 18656 16108
rect 18604 16065 18613 16099
rect 18613 16065 18647 16099
rect 18647 16065 18656 16099
rect 18604 16056 18656 16065
rect 13452 15920 13504 15972
rect 15200 15920 15252 15972
rect 15384 15988 15436 16040
rect 15476 15920 15528 15972
rect 5356 15895 5408 15904
rect 5356 15861 5365 15895
rect 5365 15861 5399 15895
rect 5399 15861 5408 15895
rect 5356 15852 5408 15861
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 6828 15852 6880 15861
rect 10692 15895 10744 15904
rect 10692 15861 10701 15895
rect 10701 15861 10735 15895
rect 10735 15861 10744 15895
rect 10692 15852 10744 15861
rect 11888 15852 11940 15904
rect 12532 15852 12584 15904
rect 13544 15852 13596 15904
rect 15292 15895 15344 15904
rect 15292 15861 15301 15895
rect 15301 15861 15335 15895
rect 15335 15861 15344 15895
rect 15292 15852 15344 15861
rect 17316 15852 17368 15904
rect 18512 15895 18564 15904
rect 18512 15861 18521 15895
rect 18521 15861 18555 15895
rect 18555 15861 18564 15895
rect 18512 15852 18564 15861
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 2780 15648 2832 15700
rect 3240 15648 3292 15700
rect 5356 15648 5408 15700
rect 6644 15648 6696 15700
rect 8300 15648 8352 15700
rect 10324 15648 10376 15700
rect 10692 15648 10744 15700
rect 14004 15691 14056 15700
rect 14004 15657 14013 15691
rect 14013 15657 14047 15691
rect 14047 15657 14056 15691
rect 14004 15648 14056 15657
rect 15292 15648 15344 15700
rect 17408 15648 17460 15700
rect 11152 15623 11204 15632
rect 1952 15512 2004 15564
rect 11152 15589 11186 15623
rect 11186 15589 11204 15623
rect 11152 15580 11204 15589
rect 14556 15580 14608 15632
rect 2964 15512 3016 15564
rect 4804 15512 4856 15564
rect 1584 15444 1636 15496
rect 6276 15512 6328 15564
rect 5908 15376 5960 15428
rect 7656 15512 7708 15564
rect 9404 15444 9456 15496
rect 9680 15376 9732 15428
rect 10968 15512 11020 15564
rect 13268 15555 13320 15564
rect 13268 15521 13277 15555
rect 13277 15521 13311 15555
rect 13311 15521 13320 15555
rect 13268 15512 13320 15521
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 14280 15512 14332 15564
rect 18788 15623 18840 15632
rect 18788 15589 18822 15623
rect 18822 15589 18840 15623
rect 18788 15580 18840 15589
rect 18144 15512 18196 15564
rect 18604 15512 18656 15564
rect 14372 15444 14424 15496
rect 14648 15487 14700 15496
rect 14648 15453 14657 15487
rect 14657 15453 14691 15487
rect 14691 15453 14700 15487
rect 14648 15444 14700 15453
rect 15844 15444 15896 15496
rect 16672 15487 16724 15496
rect 16672 15453 16681 15487
rect 16681 15453 16715 15487
rect 16715 15453 16724 15487
rect 16672 15444 16724 15453
rect 16764 15487 16816 15496
rect 16764 15453 16773 15487
rect 16773 15453 16807 15487
rect 16807 15453 16816 15487
rect 16764 15444 16816 15453
rect 14096 15376 14148 15428
rect 15384 15376 15436 15428
rect 15568 15376 15620 15428
rect 18512 15376 18564 15428
rect 3332 15351 3384 15360
rect 3332 15317 3341 15351
rect 3341 15317 3375 15351
rect 3375 15317 3384 15351
rect 3332 15308 3384 15317
rect 5448 15308 5500 15360
rect 12440 15308 12492 15360
rect 13452 15308 13504 15360
rect 19892 15351 19944 15360
rect 19892 15317 19901 15351
rect 19901 15317 19935 15351
rect 19935 15317 19944 15351
rect 19892 15308 19944 15317
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 1676 15147 1728 15156
rect 1676 15113 1685 15147
rect 1685 15113 1719 15147
rect 1719 15113 1728 15147
rect 1676 15104 1728 15113
rect 1952 14968 2004 15020
rect 4252 15104 4304 15156
rect 6276 15147 6328 15156
rect 6276 15113 6285 15147
rect 6285 15113 6319 15147
rect 6319 15113 6328 15147
rect 6276 15104 6328 15113
rect 6644 15104 6696 15156
rect 9404 15147 9456 15156
rect 9404 15113 9413 15147
rect 9413 15113 9447 15147
rect 9447 15113 9456 15147
rect 9404 15104 9456 15113
rect 10324 15104 10376 15156
rect 12532 15147 12584 15156
rect 12532 15113 12541 15147
rect 12541 15113 12575 15147
rect 12575 15113 12584 15147
rect 12532 15104 12584 15113
rect 13912 15104 13964 15156
rect 15476 15147 15528 15156
rect 15476 15113 15485 15147
rect 15485 15113 15519 15147
rect 15519 15113 15528 15147
rect 15476 15104 15528 15113
rect 16856 15104 16908 15156
rect 4804 15036 4856 15088
rect 6828 15036 6880 15088
rect 12072 15079 12124 15088
rect 12072 15045 12081 15079
rect 12081 15045 12115 15079
rect 12115 15045 12124 15079
rect 12072 15036 12124 15045
rect 15660 15036 15712 15088
rect 4344 14968 4396 15020
rect 13544 15011 13596 15020
rect 2228 14832 2280 14884
rect 4160 14900 4212 14952
rect 8668 14900 8720 14952
rect 5724 14832 5776 14884
rect 3792 14764 3844 14816
rect 5448 14764 5500 14816
rect 10232 14900 10284 14952
rect 10508 14900 10560 14952
rect 9956 14875 10008 14884
rect 9956 14841 9990 14875
rect 9990 14841 10008 14875
rect 9956 14832 10008 14841
rect 12072 14832 12124 14884
rect 10232 14764 10284 14816
rect 12900 14807 12952 14816
rect 12900 14773 12909 14807
rect 12909 14773 12943 14807
rect 12943 14773 12952 14807
rect 12900 14764 12952 14773
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 14648 15011 14700 15020
rect 14648 14977 14657 15011
rect 14657 14977 14691 15011
rect 14691 14977 14700 15011
rect 14648 14968 14700 14977
rect 17224 14968 17276 15020
rect 19340 14968 19392 15020
rect 19892 14968 19944 15020
rect 14188 14900 14240 14952
rect 14372 14943 14424 14952
rect 14372 14909 14381 14943
rect 14381 14909 14415 14943
rect 14415 14909 14424 14943
rect 14372 14900 14424 14909
rect 15936 14943 15988 14952
rect 15936 14909 15945 14943
rect 15945 14909 15979 14943
rect 15979 14909 15988 14943
rect 15936 14900 15988 14909
rect 16028 14900 16080 14952
rect 15844 14832 15896 14884
rect 16672 14832 16724 14884
rect 17224 14764 17276 14816
rect 17408 14764 17460 14816
rect 18052 14807 18104 14816
rect 18052 14773 18061 14807
rect 18061 14773 18095 14807
rect 18095 14773 18104 14807
rect 18052 14764 18104 14773
rect 18604 14900 18656 14952
rect 21364 14900 21416 14952
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 3332 14603 3384 14612
rect 3332 14569 3341 14603
rect 3341 14569 3375 14603
rect 3375 14569 3384 14603
rect 3332 14560 3384 14569
rect 4252 14560 4304 14612
rect 5448 14603 5500 14612
rect 5448 14569 5457 14603
rect 5457 14569 5491 14603
rect 5491 14569 5500 14603
rect 5448 14560 5500 14569
rect 5724 14603 5776 14612
rect 5724 14569 5733 14603
rect 5733 14569 5767 14603
rect 5767 14569 5776 14603
rect 5724 14560 5776 14569
rect 7656 14560 7708 14612
rect 9680 14603 9732 14612
rect 9680 14569 9689 14603
rect 9689 14569 9723 14603
rect 9723 14569 9732 14603
rect 9680 14560 9732 14569
rect 10508 14603 10560 14612
rect 10508 14569 10517 14603
rect 10517 14569 10551 14603
rect 10551 14569 10560 14603
rect 10508 14560 10560 14569
rect 2872 14424 2924 14476
rect 10876 14535 10928 14544
rect 10876 14501 10885 14535
rect 10885 14501 10919 14535
rect 10919 14501 10928 14535
rect 10876 14492 10928 14501
rect 6920 14424 6972 14476
rect 8392 14424 8444 14476
rect 3792 14356 3844 14408
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 6828 14399 6880 14408
rect 2780 14220 2832 14272
rect 3332 14220 3384 14272
rect 6276 14288 6328 14340
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 13268 14560 13320 14612
rect 13544 14560 13596 14612
rect 13728 14560 13780 14612
rect 16672 14603 16724 14612
rect 16672 14569 16681 14603
rect 16681 14569 16715 14603
rect 16715 14569 16724 14603
rect 16672 14560 16724 14569
rect 12440 14492 12492 14544
rect 13636 14424 13688 14476
rect 19340 14492 19392 14544
rect 15844 14424 15896 14476
rect 15936 14424 15988 14476
rect 18512 14424 18564 14476
rect 16948 14399 17000 14408
rect 16948 14365 16957 14399
rect 16957 14365 16991 14399
rect 16991 14365 17000 14399
rect 16948 14356 17000 14365
rect 19340 14399 19392 14408
rect 19340 14365 19349 14399
rect 19349 14365 19383 14399
rect 19383 14365 19392 14399
rect 19340 14356 19392 14365
rect 7104 14220 7156 14272
rect 8024 14220 8076 14272
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 11888 14220 11940 14272
rect 14372 14220 14424 14272
rect 14556 14263 14608 14272
rect 14556 14229 14565 14263
rect 14565 14229 14599 14263
rect 14599 14229 14608 14263
rect 14556 14220 14608 14229
rect 18696 14220 18748 14272
rect 21364 14263 21416 14272
rect 21364 14229 21373 14263
rect 21373 14229 21407 14263
rect 21407 14229 21416 14263
rect 21364 14220 21416 14229
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 1492 14016 1544 14068
rect 5908 14059 5960 14068
rect 1492 13855 1544 13864
rect 1492 13821 1501 13855
rect 1501 13821 1535 13855
rect 1535 13821 1544 13855
rect 1492 13812 1544 13821
rect 5908 14025 5917 14059
rect 5917 14025 5951 14059
rect 5951 14025 5960 14059
rect 5908 14016 5960 14025
rect 7196 14016 7248 14068
rect 8024 14016 8076 14068
rect 12808 14016 12860 14068
rect 14188 14059 14240 14068
rect 14188 14025 14197 14059
rect 14197 14025 14231 14059
rect 14231 14025 14240 14059
rect 14188 14016 14240 14025
rect 16304 14016 16356 14068
rect 17960 14016 18012 14068
rect 6276 13948 6328 14000
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 2964 13923 3016 13932
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 9956 13948 10008 14000
rect 13452 13948 13504 14000
rect 11888 13923 11940 13932
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 3792 13744 3844 13796
rect 5724 13812 5776 13864
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 3148 13676 3200 13728
rect 3884 13719 3936 13728
rect 3884 13685 3893 13719
rect 3893 13685 3927 13719
rect 3927 13685 3936 13719
rect 3884 13676 3936 13685
rect 5448 13744 5500 13796
rect 11888 13889 11897 13923
rect 11897 13889 11931 13923
rect 11931 13889 11940 13923
rect 11888 13880 11940 13889
rect 16028 13948 16080 14000
rect 15660 13923 15712 13932
rect 15660 13889 15669 13923
rect 15669 13889 15703 13923
rect 15703 13889 15712 13923
rect 15660 13880 15712 13889
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 16396 13880 16448 13932
rect 8208 13812 8260 13864
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 8760 13812 8812 13821
rect 12348 13812 12400 13864
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 13728 13812 13780 13864
rect 14372 13812 14424 13864
rect 19248 13948 19300 14000
rect 16672 13880 16724 13932
rect 18052 13880 18104 13932
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 16948 13812 17000 13864
rect 7380 13744 7432 13796
rect 9588 13744 9640 13796
rect 4712 13676 4764 13728
rect 10416 13676 10468 13728
rect 11704 13719 11756 13728
rect 11704 13685 11713 13719
rect 11713 13685 11747 13719
rect 11747 13685 11756 13719
rect 11704 13676 11756 13685
rect 14556 13719 14608 13728
rect 14556 13685 14565 13719
rect 14565 13685 14599 13719
rect 14599 13685 14608 13719
rect 14556 13676 14608 13685
rect 19340 13744 19392 13796
rect 15292 13676 15344 13728
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 2872 13472 2924 13524
rect 3884 13472 3936 13524
rect 5448 13515 5500 13524
rect 5448 13481 5457 13515
rect 5457 13481 5491 13515
rect 5491 13481 5500 13515
rect 5448 13472 5500 13481
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 6920 13472 6972 13524
rect 7196 13472 7248 13524
rect 10784 13515 10836 13524
rect 10784 13481 10793 13515
rect 10793 13481 10827 13515
rect 10827 13481 10836 13515
rect 10784 13472 10836 13481
rect 11888 13472 11940 13524
rect 13084 13472 13136 13524
rect 1492 13404 1544 13456
rect 5816 13404 5868 13456
rect 3148 13336 3200 13388
rect 5908 13336 5960 13388
rect 3792 13268 3844 13320
rect 7564 13404 7616 13456
rect 14464 13472 14516 13524
rect 18696 13404 18748 13456
rect 6920 13336 6972 13388
rect 7380 13379 7432 13388
rect 7380 13345 7389 13379
rect 7389 13345 7423 13379
rect 7423 13345 7432 13379
rect 7380 13336 7432 13345
rect 9496 13336 9548 13388
rect 10048 13379 10100 13388
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 13452 13336 13504 13388
rect 8208 13268 8260 13320
rect 9956 13268 10008 13320
rect 7288 13200 7340 13252
rect 9312 13200 9364 13252
rect 9588 13200 9640 13252
rect 3976 13132 4028 13184
rect 10600 13132 10652 13184
rect 12992 13268 13044 13320
rect 13544 13268 13596 13320
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 14096 13200 14148 13252
rect 15844 13311 15896 13320
rect 15844 13277 15853 13311
rect 15853 13277 15887 13311
rect 15887 13277 15896 13311
rect 15844 13268 15896 13277
rect 17040 13268 17092 13320
rect 17776 13311 17828 13320
rect 17776 13277 17785 13311
rect 17785 13277 17819 13311
rect 17819 13277 17828 13311
rect 17776 13268 17828 13277
rect 14924 13200 14976 13252
rect 17684 13200 17736 13252
rect 12440 13132 12492 13184
rect 12716 13132 12768 13184
rect 12992 13132 13044 13184
rect 14004 13132 14056 13184
rect 15108 13132 15160 13184
rect 17132 13132 17184 13184
rect 19156 13175 19208 13184
rect 19156 13141 19165 13175
rect 19165 13141 19199 13175
rect 19199 13141 19208 13175
rect 19156 13132 19208 13141
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 1952 12971 2004 12980
rect 1952 12937 1961 12971
rect 1961 12937 1995 12971
rect 1995 12937 2004 12971
rect 1952 12928 2004 12937
rect 3056 12928 3108 12980
rect 3608 12971 3660 12980
rect 3608 12937 3617 12971
rect 3617 12937 3651 12971
rect 3651 12937 3660 12971
rect 3608 12928 3660 12937
rect 4160 12928 4212 12980
rect 5816 12971 5868 12980
rect 5816 12937 5825 12971
rect 5825 12937 5859 12971
rect 5859 12937 5868 12971
rect 5816 12928 5868 12937
rect 11704 12928 11756 12980
rect 12348 12928 12400 12980
rect 13544 12971 13596 12980
rect 13544 12937 13553 12971
rect 13553 12937 13587 12971
rect 13587 12937 13596 12971
rect 13544 12928 13596 12937
rect 14464 12928 14516 12980
rect 16396 12971 16448 12980
rect 16396 12937 16405 12971
rect 16405 12937 16439 12971
rect 16439 12937 16448 12971
rect 16396 12928 16448 12937
rect 16580 12928 16632 12980
rect 18880 12928 18932 12980
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 9496 12835 9548 12844
rect 9496 12801 9505 12835
rect 9505 12801 9539 12835
rect 9539 12801 9548 12835
rect 9496 12792 9548 12801
rect 12992 12835 13044 12844
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 13452 12792 13504 12844
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 2044 12724 2096 12776
rect 2780 12724 2832 12776
rect 3148 12724 3200 12776
rect 3424 12767 3476 12776
rect 3424 12733 3433 12767
rect 3433 12733 3467 12767
rect 3467 12733 3476 12767
rect 3424 12724 3476 12733
rect 3792 12724 3844 12776
rect 7104 12767 7156 12776
rect 7104 12733 7138 12767
rect 7138 12733 7156 12767
rect 7104 12724 7156 12733
rect 4804 12656 4856 12708
rect 5908 12656 5960 12708
rect 10048 12724 10100 12776
rect 11888 12724 11940 12776
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 14280 12724 14332 12776
rect 14648 12724 14700 12776
rect 17040 12767 17092 12776
rect 17040 12733 17049 12767
rect 17049 12733 17083 12767
rect 17083 12733 17092 12767
rect 17040 12724 17092 12733
rect 17684 12792 17736 12844
rect 18696 12835 18748 12844
rect 18696 12801 18705 12835
rect 18705 12801 18739 12835
rect 18739 12801 18748 12835
rect 18696 12792 18748 12801
rect 19156 12792 19208 12844
rect 7748 12656 7800 12708
rect 12808 12656 12860 12708
rect 3240 12588 3292 12640
rect 6920 12588 6972 12640
rect 7196 12588 7248 12640
rect 8944 12631 8996 12640
rect 8944 12597 8953 12631
rect 8953 12597 8987 12631
rect 8987 12597 8996 12631
rect 11060 12631 11112 12640
rect 8944 12588 8996 12597
rect 11060 12597 11069 12631
rect 11069 12597 11103 12631
rect 11103 12597 11112 12631
rect 11060 12588 11112 12597
rect 11888 12588 11940 12640
rect 12256 12588 12308 12640
rect 14924 12656 14976 12708
rect 16764 12656 16816 12708
rect 18788 12724 18840 12776
rect 14280 12588 14332 12640
rect 19248 12588 19300 12640
rect 19432 12631 19484 12640
rect 19432 12597 19441 12631
rect 19441 12597 19475 12631
rect 19475 12597 19484 12631
rect 19432 12588 19484 12597
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 3516 12384 3568 12436
rect 9312 12427 9364 12436
rect 3148 12359 3200 12368
rect 3148 12325 3157 12359
rect 3157 12325 3191 12359
rect 3191 12325 3200 12359
rect 3148 12316 3200 12325
rect 2136 12291 2188 12300
rect 2136 12257 2145 12291
rect 2145 12257 2179 12291
rect 2179 12257 2188 12291
rect 2136 12248 2188 12257
rect 4160 12248 4212 12300
rect 5448 12248 5500 12300
rect 7656 12316 7708 12368
rect 8484 12316 8536 12368
rect 9036 12316 9088 12368
rect 9312 12393 9321 12427
rect 9321 12393 9355 12427
rect 9355 12393 9364 12427
rect 9312 12384 9364 12393
rect 11888 12384 11940 12436
rect 14740 12384 14792 12436
rect 16764 12384 16816 12436
rect 19248 12384 19300 12436
rect 11152 12316 11204 12368
rect 11796 12316 11848 12368
rect 13084 12316 13136 12368
rect 15844 12316 15896 12368
rect 6828 12248 6880 12300
rect 7012 12291 7064 12300
rect 7012 12257 7021 12291
rect 7021 12257 7055 12291
rect 7055 12257 7064 12291
rect 7012 12248 7064 12257
rect 8760 12248 8812 12300
rect 9496 12248 9548 12300
rect 10324 12248 10376 12300
rect 11980 12248 12032 12300
rect 12716 12248 12768 12300
rect 14464 12291 14516 12300
rect 14464 12257 14473 12291
rect 14473 12257 14507 12291
rect 14507 12257 14516 12291
rect 14464 12248 14516 12257
rect 14648 12248 14700 12300
rect 17592 12316 17644 12368
rect 17776 12316 17828 12368
rect 18052 12248 18104 12300
rect 3424 12180 3476 12232
rect 3792 12180 3844 12232
rect 7196 12180 7248 12232
rect 10416 12112 10468 12164
rect 13636 12180 13688 12232
rect 4804 12044 4856 12096
rect 5540 12044 5592 12096
rect 5908 12044 5960 12096
rect 6092 12087 6144 12096
rect 6092 12053 6101 12087
rect 6101 12053 6135 12087
rect 6135 12053 6144 12087
rect 6092 12044 6144 12053
rect 6552 12087 6604 12096
rect 6552 12053 6561 12087
rect 6561 12053 6595 12087
rect 6595 12053 6604 12087
rect 6552 12044 6604 12053
rect 11060 12044 11112 12096
rect 11796 12044 11848 12096
rect 14188 12112 14240 12164
rect 15200 12180 15252 12232
rect 18880 12223 18932 12232
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 18144 12044 18196 12096
rect 18788 12044 18840 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 4068 11840 4120 11892
rect 8484 11883 8536 11892
rect 2136 11772 2188 11824
rect 2044 11747 2096 11756
rect 2044 11713 2053 11747
rect 2053 11713 2087 11747
rect 2087 11713 2096 11747
rect 2044 11704 2096 11713
rect 2780 11747 2832 11756
rect 2780 11713 2789 11747
rect 2789 11713 2823 11747
rect 2823 11713 2832 11747
rect 6552 11772 6604 11824
rect 8484 11849 8493 11883
rect 8493 11849 8527 11883
rect 8527 11849 8536 11883
rect 8484 11840 8536 11849
rect 11152 11840 11204 11892
rect 11244 11840 11296 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 15844 11840 15896 11892
rect 19432 11840 19484 11892
rect 17592 11772 17644 11824
rect 2780 11704 2832 11713
rect 4804 11704 4856 11756
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 9496 11704 9548 11756
rect 11796 11747 11848 11756
rect 11796 11713 11805 11747
rect 11805 11713 11839 11747
rect 11839 11713 11848 11747
rect 11796 11704 11848 11713
rect 12532 11747 12584 11756
rect 1952 11636 2004 11688
rect 5724 11636 5776 11688
rect 6184 11636 6236 11688
rect 6920 11568 6972 11620
rect 9772 11636 9824 11688
rect 10416 11636 10468 11688
rect 11060 11636 11112 11688
rect 12532 11713 12541 11747
rect 12541 11713 12575 11747
rect 12575 11713 12584 11747
rect 12532 11704 12584 11713
rect 14188 11747 14240 11756
rect 14188 11713 14197 11747
rect 14197 11713 14231 11747
rect 14231 11713 14240 11747
rect 14188 11704 14240 11713
rect 18052 11704 18104 11756
rect 18696 11704 18748 11756
rect 7288 11568 7340 11620
rect 8484 11568 8536 11620
rect 10140 11568 10192 11620
rect 14280 11636 14332 11688
rect 18880 11636 18932 11688
rect 15200 11568 15252 11620
rect 15476 11568 15528 11620
rect 5632 11500 5684 11552
rect 6000 11500 6052 11552
rect 6828 11500 6880 11552
rect 7472 11500 7524 11552
rect 8392 11500 8444 11552
rect 11060 11543 11112 11552
rect 11060 11509 11069 11543
rect 11069 11509 11103 11543
rect 11103 11509 11112 11543
rect 11060 11500 11112 11509
rect 12440 11500 12492 11552
rect 12716 11500 12768 11552
rect 13452 11543 13504 11552
rect 13452 11509 13461 11543
rect 13461 11509 13495 11543
rect 13495 11509 13504 11543
rect 13452 11500 13504 11509
rect 17500 11500 17552 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 1952 11339 2004 11348
rect 1952 11305 1961 11339
rect 1961 11305 1995 11339
rect 1995 11305 2004 11339
rect 1952 11296 2004 11305
rect 4896 11296 4948 11348
rect 7564 11296 7616 11348
rect 8944 11296 8996 11348
rect 9496 11296 9548 11348
rect 10324 11339 10376 11348
rect 10324 11305 10333 11339
rect 10333 11305 10367 11339
rect 10367 11305 10376 11339
rect 10324 11296 10376 11305
rect 12624 11339 12676 11348
rect 12624 11305 12633 11339
rect 12633 11305 12667 11339
rect 12667 11305 12676 11339
rect 12624 11296 12676 11305
rect 13636 11339 13688 11348
rect 13636 11305 13645 11339
rect 13645 11305 13679 11339
rect 13679 11305 13688 11339
rect 13636 11296 13688 11305
rect 13820 11296 13872 11348
rect 14464 11296 14516 11348
rect 3976 11228 4028 11280
rect 6920 11228 6972 11280
rect 7012 11271 7064 11280
rect 7012 11237 7021 11271
rect 7021 11237 7055 11271
rect 7055 11237 7064 11271
rect 7012 11228 7064 11237
rect 8484 11228 8536 11280
rect 8576 11228 8628 11280
rect 2320 11203 2372 11212
rect 2320 11169 2329 11203
rect 2329 11169 2363 11203
rect 2363 11169 2372 11203
rect 2320 11160 2372 11169
rect 4068 11160 4120 11212
rect 4344 11160 4396 11212
rect 6000 11160 6052 11212
rect 6092 11160 6144 11212
rect 2688 11092 2740 11144
rect 2412 11024 2464 11076
rect 4160 11024 4212 11076
rect 5632 11092 5684 11144
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 7472 11160 7524 11212
rect 8024 11203 8076 11212
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 8024 11160 8076 11169
rect 12440 11228 12492 11280
rect 16120 11228 16172 11280
rect 18144 11228 18196 11280
rect 11244 11203 11296 11212
rect 11244 11169 11278 11203
rect 11278 11169 11296 11203
rect 11244 11160 11296 11169
rect 12532 11160 12584 11212
rect 13452 11160 13504 11212
rect 16304 11160 16356 11212
rect 17592 11160 17644 11212
rect 6184 11067 6236 11076
rect 6184 11033 6193 11067
rect 6193 11033 6227 11067
rect 6227 11033 6236 11067
rect 6184 11024 6236 11033
rect 8116 11024 8168 11076
rect 12164 11092 12216 11144
rect 8484 11024 8536 11076
rect 4804 10956 4856 11008
rect 9404 11024 9456 11076
rect 12716 11024 12768 11076
rect 14372 11092 14424 11144
rect 9220 10956 9272 11008
rect 14004 10956 14056 11008
rect 17040 10999 17092 11008
rect 17040 10965 17049 10999
rect 17049 10965 17083 10999
rect 17083 10965 17092 10999
rect 17040 10956 17092 10965
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 2320 10752 2372 10804
rect 4160 10795 4212 10804
rect 4160 10761 4169 10795
rect 4169 10761 4203 10795
rect 4203 10761 4212 10795
rect 4160 10752 4212 10761
rect 4896 10752 4948 10804
rect 5724 10795 5776 10804
rect 5724 10761 5733 10795
rect 5733 10761 5767 10795
rect 5767 10761 5776 10795
rect 5724 10752 5776 10761
rect 3884 10684 3936 10736
rect 2320 10616 2372 10668
rect 4528 10616 4580 10668
rect 6460 10684 6512 10736
rect 8116 10752 8168 10804
rect 9220 10752 9272 10804
rect 9404 10752 9456 10804
rect 10876 10752 10928 10804
rect 11244 10752 11296 10804
rect 14372 10752 14424 10804
rect 15476 10795 15528 10804
rect 15476 10761 15485 10795
rect 15485 10761 15519 10795
rect 15519 10761 15528 10795
rect 15476 10752 15528 10761
rect 17684 10727 17736 10736
rect 17684 10693 17693 10727
rect 17693 10693 17727 10727
rect 17727 10693 17736 10727
rect 17684 10684 17736 10693
rect 6736 10616 6788 10668
rect 2780 10591 2832 10600
rect 2780 10557 2789 10591
rect 2789 10557 2823 10591
rect 2823 10557 2832 10591
rect 2780 10548 2832 10557
rect 5264 10591 5316 10600
rect 5264 10557 5273 10591
rect 5273 10557 5307 10591
rect 5307 10557 5316 10591
rect 5264 10548 5316 10557
rect 6644 10548 6696 10600
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 9496 10616 9548 10668
rect 16304 10659 16356 10668
rect 16304 10625 16313 10659
rect 16313 10625 16347 10659
rect 16347 10625 16356 10659
rect 16304 10616 16356 10625
rect 7656 10548 7708 10600
rect 8484 10591 8536 10600
rect 8484 10557 8493 10591
rect 8493 10557 8527 10591
rect 8527 10557 8536 10591
rect 8484 10548 8536 10557
rect 3516 10480 3568 10532
rect 3976 10480 4028 10532
rect 8944 10480 8996 10532
rect 2136 10455 2188 10464
rect 2136 10421 2145 10455
rect 2145 10421 2179 10455
rect 2179 10421 2188 10455
rect 2136 10412 2188 10421
rect 2872 10412 2924 10464
rect 6092 10455 6144 10464
rect 6092 10421 6101 10455
rect 6101 10421 6135 10455
rect 6135 10421 6144 10455
rect 6092 10412 6144 10421
rect 7380 10412 7432 10464
rect 8208 10412 8260 10464
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12716 10591 12768 10600
rect 12440 10548 12492 10557
rect 12716 10557 12750 10591
rect 12750 10557 12768 10591
rect 12716 10548 12768 10557
rect 14372 10591 14424 10600
rect 14372 10557 14406 10591
rect 14406 10557 14424 10591
rect 14372 10548 14424 10557
rect 17040 10548 17092 10600
rect 11060 10480 11112 10532
rect 12532 10480 12584 10532
rect 12256 10412 12308 10464
rect 12440 10412 12492 10464
rect 18052 10455 18104 10464
rect 18052 10421 18061 10455
rect 18061 10421 18095 10455
rect 18095 10421 18104 10455
rect 18052 10412 18104 10421
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 2136 10208 2188 10260
rect 4068 10251 4120 10260
rect 4068 10217 4077 10251
rect 4077 10217 4111 10251
rect 4111 10217 4120 10251
rect 4068 10208 4120 10217
rect 4528 10251 4580 10260
rect 4528 10217 4537 10251
rect 4537 10217 4571 10251
rect 4571 10217 4580 10251
rect 4528 10208 4580 10217
rect 4988 10208 5040 10260
rect 6736 10251 6788 10260
rect 2320 10140 2372 10192
rect 3792 10140 3844 10192
rect 2780 10072 2832 10124
rect 3240 10072 3292 10124
rect 5264 10072 5316 10124
rect 6184 10140 6236 10192
rect 6736 10217 6745 10251
rect 6745 10217 6779 10251
rect 6779 10217 6788 10251
rect 6736 10208 6788 10217
rect 7380 10251 7432 10260
rect 7380 10217 7389 10251
rect 7389 10217 7423 10251
rect 7423 10217 7432 10251
rect 7380 10208 7432 10217
rect 9864 10208 9916 10260
rect 10048 10251 10100 10260
rect 10048 10217 10057 10251
rect 10057 10217 10091 10251
rect 10091 10217 10100 10251
rect 10048 10208 10100 10217
rect 11980 10208 12032 10260
rect 12164 10140 12216 10192
rect 16856 10208 16908 10260
rect 18052 10208 18104 10260
rect 3516 10004 3568 10056
rect 4804 10004 4856 10056
rect 7932 10004 7984 10056
rect 8208 10004 8260 10056
rect 8852 10047 8904 10056
rect 8852 10013 8861 10047
rect 8861 10013 8895 10047
rect 8895 10013 8904 10047
rect 8852 10004 8904 10013
rect 8944 10047 8996 10056
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 10692 10072 10744 10124
rect 12256 10072 12308 10124
rect 13452 10072 13504 10124
rect 14740 10072 14792 10124
rect 8944 10004 8996 10013
rect 9864 9936 9916 9988
rect 11152 9936 11204 9988
rect 11244 9936 11296 9988
rect 13544 10004 13596 10056
rect 15108 10004 15160 10056
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 17132 10047 17184 10056
rect 17132 10013 17141 10047
rect 17141 10013 17175 10047
rect 17175 10013 17184 10047
rect 17132 10004 17184 10013
rect 2688 9868 2740 9920
rect 9588 9868 9640 9920
rect 14096 9868 14148 9920
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 2872 9707 2924 9716
rect 2872 9673 2881 9707
rect 2881 9673 2915 9707
rect 2915 9673 2924 9707
rect 2872 9664 2924 9673
rect 6092 9664 6144 9716
rect 8944 9664 8996 9716
rect 10048 9664 10100 9716
rect 15108 9707 15160 9716
rect 15108 9673 15117 9707
rect 15117 9673 15151 9707
rect 15151 9673 15160 9707
rect 15108 9664 15160 9673
rect 1860 9596 1912 9648
rect 11152 9639 11204 9648
rect 11152 9605 11161 9639
rect 11161 9605 11195 9639
rect 11195 9605 11204 9639
rect 11152 9596 11204 9605
rect 2780 9528 2832 9580
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 3516 9571 3568 9580
rect 3516 9537 3525 9571
rect 3525 9537 3559 9571
rect 3559 9537 3568 9571
rect 3516 9528 3568 9537
rect 4804 9571 4856 9580
rect 4804 9537 4813 9571
rect 4813 9537 4847 9571
rect 4847 9537 4856 9571
rect 4804 9528 4856 9537
rect 6920 9528 6972 9580
rect 7932 9528 7984 9580
rect 9772 9528 9824 9580
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 3976 9460 4028 9512
rect 3056 9324 3108 9376
rect 5632 9392 5684 9444
rect 7380 9460 7432 9512
rect 7656 9460 7708 9512
rect 17408 9460 17460 9512
rect 8668 9392 8720 9444
rect 4252 9367 4304 9376
rect 4252 9333 4261 9367
rect 4261 9333 4295 9367
rect 4295 9333 4304 9367
rect 4252 9324 4304 9333
rect 4620 9367 4672 9376
rect 4620 9333 4629 9367
rect 4629 9333 4663 9367
rect 4663 9333 4672 9367
rect 4620 9324 4672 9333
rect 4896 9324 4948 9376
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 11152 9324 11204 9376
rect 13360 9324 13412 9376
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 1400 9120 1452 9172
rect 4620 9163 4672 9172
rect 4620 9129 4629 9163
rect 4629 9129 4663 9163
rect 4663 9129 4672 9163
rect 4620 9120 4672 9129
rect 8208 9120 8260 9172
rect 8392 9120 8444 9172
rect 2228 8984 2280 9036
rect 2596 9027 2648 9036
rect 2596 8993 2630 9027
rect 2630 8993 2648 9027
rect 2596 8984 2648 8993
rect 4068 9052 4120 9104
rect 17316 9052 17368 9104
rect 3148 8984 3200 9036
rect 4988 9027 5040 9036
rect 4988 8993 4997 9027
rect 4997 8993 5031 9027
rect 5031 8993 5040 9027
rect 4988 8984 5040 8993
rect 3884 8916 3936 8968
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 7656 8916 7708 8968
rect 8852 8848 8904 8900
rect 3700 8823 3752 8832
rect 3700 8789 3709 8823
rect 3709 8789 3743 8823
rect 3743 8789 3752 8823
rect 3700 8780 3752 8789
rect 3792 8780 3844 8832
rect 6276 8780 6328 8832
rect 7288 8780 7340 8832
rect 8484 8780 8536 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 4804 8508 4856 8560
rect 2228 8483 2280 8492
rect 2228 8449 2237 8483
rect 2237 8449 2271 8483
rect 2271 8449 2280 8483
rect 2228 8440 2280 8449
rect 8024 8576 8076 8628
rect 11888 8576 11940 8628
rect 11152 8508 11204 8560
rect 2964 8372 3016 8424
rect 3148 8415 3200 8424
rect 3148 8381 3157 8415
rect 3157 8381 3191 8415
rect 3191 8381 3200 8415
rect 3148 8372 3200 8381
rect 3700 8372 3752 8424
rect 8760 8440 8812 8492
rect 7380 8372 7432 8424
rect 8392 8372 8444 8424
rect 5540 8304 5592 8356
rect 7104 8347 7156 8356
rect 7104 8313 7138 8347
rect 7138 8313 7156 8347
rect 7104 8304 7156 8313
rect 3976 8236 4028 8288
rect 5724 8236 5776 8288
rect 5816 8236 5868 8288
rect 7656 8236 7708 8288
rect 17500 8236 17552 8288
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 2964 8075 3016 8084
rect 1768 7964 1820 8016
rect 2964 8041 2973 8075
rect 2973 8041 3007 8075
rect 3007 8041 3016 8075
rect 2964 8032 3016 8041
rect 4252 8032 4304 8084
rect 4436 8032 4488 8084
rect 5816 8032 5868 8084
rect 7104 8075 7156 8084
rect 7104 8041 7113 8075
rect 7113 8041 7147 8075
rect 7147 8041 7156 8075
rect 7104 8032 7156 8041
rect 8484 8032 8536 8084
rect 4160 7896 4212 7948
rect 4804 7964 4856 8016
rect 3976 7828 4028 7880
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 8760 7964 8812 8016
rect 8852 7964 8904 8016
rect 14740 8032 14792 8084
rect 7380 7939 7432 7948
rect 7380 7905 7389 7939
rect 7389 7905 7423 7939
rect 7423 7905 7432 7939
rect 7380 7896 7432 7905
rect 7656 7939 7708 7948
rect 7656 7905 7690 7939
rect 7690 7905 7708 7939
rect 7656 7896 7708 7905
rect 8484 7896 8536 7948
rect 8668 7760 8720 7812
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 4160 7531 4212 7540
rect 4160 7497 4169 7531
rect 4169 7497 4203 7531
rect 4203 7497 4212 7531
rect 4160 7488 4212 7497
rect 8208 7488 8260 7540
rect 19708 7488 19760 7540
rect 7104 7463 7156 7472
rect 7104 7429 7113 7463
rect 7113 7429 7147 7463
rect 7147 7429 7156 7463
rect 7104 7420 7156 7429
rect 19524 7420 19576 7472
rect 4712 7395 4764 7404
rect 4712 7361 4721 7395
rect 4721 7361 4755 7395
rect 4755 7361 4764 7395
rect 4712 7352 4764 7361
rect 6460 7352 6512 7404
rect 6736 7216 6788 7268
rect 8760 7395 8812 7404
rect 8760 7361 8769 7395
rect 8769 7361 8803 7395
rect 8803 7361 8812 7395
rect 8760 7352 8812 7361
rect 7840 7284 7892 7336
rect 18788 7284 18840 7336
rect 3792 7191 3844 7200
rect 3792 7157 3801 7191
rect 3801 7157 3835 7191
rect 3835 7157 3844 7191
rect 3792 7148 3844 7157
rect 6276 7148 6328 7200
rect 6368 7191 6420 7200
rect 6368 7157 6377 7191
rect 6377 7157 6411 7191
rect 6411 7157 6420 7191
rect 6368 7148 6420 7157
rect 7748 7148 7800 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 2780 6944 2832 6996
rect 6368 6944 6420 6996
rect 7104 6944 7156 6996
rect 3976 6808 4028 6860
rect 5632 6740 5684 6792
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 7656 6740 7708 6792
rect 20444 6672 20496 6724
rect 8484 6604 8536 6656
rect 8576 6604 8628 6656
rect 18788 6604 18840 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 20904 6400 20956 6452
rect 4068 6060 4120 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 21088 5899 21140 5908
rect 21088 5865 21097 5899
rect 21097 5865 21131 5899
rect 21131 5865 21140 5899
rect 21088 5856 21140 5865
rect 20444 5720 20496 5772
rect 20444 5559 20496 5568
rect 20444 5525 20453 5559
rect 20453 5525 20487 5559
rect 20487 5525 20496 5559
rect 20444 5516 20496 5525
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 4068 5312 4120 5364
rect 20444 5312 20496 5364
rect 20996 5355 21048 5364
rect 20996 5321 21005 5355
rect 21005 5321 21039 5355
rect 21039 5321 21048 5355
rect 20996 5312 21048 5321
rect 3976 5244 4028 5296
rect 14648 5244 14700 5296
rect 4068 4972 4120 5024
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 11704 4768 11756 4820
rect 12072 4768 12124 4820
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 3516 2048 3568 2100
rect 6828 2048 6880 2100
rect 3332 1300 3384 1352
rect 5540 1300 5592 1352
<< metal2 >>
rect 202 22200 258 23000
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2870 22264 2926 22273
rect 216 19145 244 22200
rect 202 19136 258 19145
rect 202 19071 258 19080
rect 676 18154 704 22200
rect 1136 18737 1164 22200
rect 1596 20890 1624 22200
rect 1950 21312 2006 21321
rect 1950 21247 2006 21256
rect 1596 20862 1716 20890
rect 1582 20768 1638 20777
rect 1582 20703 1638 20712
rect 1490 19816 1546 19825
rect 1490 19751 1546 19760
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1412 18902 1440 19246
rect 1400 18896 1452 18902
rect 1400 18838 1452 18844
rect 1122 18728 1178 18737
rect 1122 18663 1178 18672
rect 664 18148 716 18154
rect 664 18090 716 18096
rect 1398 14240 1454 14249
rect 1398 14175 1454 14184
rect 1412 9178 1440 14175
rect 1504 14074 1532 19751
rect 1596 19514 1624 20703
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1688 19174 1716 20862
rect 1964 20602 1992 21247
rect 1952 20596 2004 20602
rect 1952 20538 2004 20544
rect 1768 20392 1820 20398
rect 1768 20334 1820 20340
rect 1860 20392 1912 20398
rect 1860 20334 1912 20340
rect 1780 19378 1808 20334
rect 1872 19922 1900 20334
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1676 19168 1728 19174
rect 1676 19110 1728 19116
rect 2056 18630 2084 22200
rect 2516 18748 2544 22200
rect 2870 22199 2926 22208
rect 2962 22200 3018 23000
rect 3238 22672 3294 22681
rect 3238 22607 3294 22616
rect 2884 21842 2912 22199
rect 2976 21962 3004 22200
rect 2964 21956 3016 21962
rect 2964 21898 3016 21904
rect 2884 21814 3004 21842
rect 2778 21720 2834 21729
rect 2778 21655 2834 21664
rect 2792 20602 2820 21655
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2872 19984 2924 19990
rect 2872 19926 2924 19932
rect 2688 19712 2740 19718
rect 2688 19654 2740 19660
rect 2700 19310 2728 19654
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 2596 19168 2648 19174
rect 2594 19136 2596 19145
rect 2648 19136 2650 19145
rect 2594 19071 2650 19080
rect 2516 18720 2636 18748
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 1766 18456 1822 18465
rect 1766 18391 1822 18400
rect 1780 17882 1808 18391
rect 1860 18216 1912 18222
rect 1858 18184 1860 18193
rect 1912 18184 1914 18193
rect 1858 18119 1914 18128
rect 2608 18086 2636 18720
rect 2700 18290 2728 19246
rect 2884 18970 2912 19926
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2778 18864 2834 18873
rect 2778 18799 2834 18808
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 1952 18080 2004 18086
rect 2504 18080 2556 18086
rect 1952 18022 2004 18028
rect 2502 18048 2504 18057
rect 2596 18080 2648 18086
rect 2556 18048 2558 18057
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1596 17270 1624 17682
rect 1964 17513 1992 18022
rect 2596 18022 2648 18028
rect 2502 17983 2558 17992
rect 2044 17808 2096 17814
rect 2044 17750 2096 17756
rect 1950 17504 2006 17513
rect 1950 17439 2006 17448
rect 1584 17264 1636 17270
rect 1584 17206 1636 17212
rect 2056 17134 2084 17750
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 2044 17128 2096 17134
rect 1674 17096 1730 17105
rect 2044 17070 2096 17076
rect 1674 17031 1730 17040
rect 1688 16998 1716 17031
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 2148 16794 2176 17682
rect 2136 16788 2188 16794
rect 2136 16730 2188 16736
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 1674 16552 1730 16561
rect 1674 16487 1730 16496
rect 1688 16250 1716 16487
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1674 16144 1730 16153
rect 2240 16114 2268 16594
rect 1674 16079 1730 16088
rect 2228 16108 2280 16114
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 1596 15502 1624 15982
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1688 15162 1716 16079
rect 2228 16050 2280 16056
rect 2792 15706 2820 18799
rect 2976 17882 3004 21814
rect 3054 20360 3110 20369
rect 3054 20295 3110 20304
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 3068 16726 3096 20295
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 3160 18970 3188 20198
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 3160 16726 3188 17070
rect 3056 16720 3108 16726
rect 3056 16662 3108 16668
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 3252 15706 3280 22607
rect 3422 22200 3478 23000
rect 3882 22200 3938 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6182 22200 6238 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 3436 19224 3464 22200
rect 3700 19712 3752 19718
rect 3700 19654 3752 19660
rect 3606 19408 3662 19417
rect 3606 19343 3662 19352
rect 3436 19196 3556 19224
rect 3422 19136 3478 19145
rect 3422 19071 3478 19080
rect 3436 18902 3464 19071
rect 3424 18896 3476 18902
rect 3528 18873 3556 19196
rect 3424 18838 3476 18844
rect 3514 18864 3570 18873
rect 3514 18799 3570 18808
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3436 16046 3464 17478
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3238 15600 3294 15609
rect 1952 15564 2004 15570
rect 1952 15506 2004 15512
rect 2964 15564 3016 15570
rect 3238 15535 3294 15544
rect 2964 15506 3016 15512
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1964 15026 1992 15506
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 2228 14884 2280 14890
rect 2228 14826 2280 14832
rect 1858 14648 1914 14657
rect 1858 14583 1914 14592
rect 1492 14068 1544 14074
rect 1492 14010 1544 14016
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1504 13462 1532 13806
rect 1492 13456 1544 13462
rect 1492 13398 1544 13404
rect 1872 9654 1900 14583
rect 2240 13938 2268 14826
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2792 13870 2820 14214
rect 2780 13864 2832 13870
rect 1950 13832 2006 13841
rect 2780 13806 2832 13812
rect 1950 13767 2006 13776
rect 1964 12986 1992 13767
rect 2884 13530 2912 14418
rect 2976 13938 3004 15506
rect 3054 15192 3110 15201
rect 3054 15127 3110 15136
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 3068 12986 3096 15127
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3160 13394 3188 13670
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 2056 11762 2084 12718
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2148 11830 2176 12242
rect 2136 11824 2188 11830
rect 2136 11766 2188 11772
rect 2792 11762 2820 12718
rect 3160 12374 3188 12718
rect 3252 12646 3280 15535
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3344 14618 3372 15302
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3344 14278 3372 14554
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 3436 14090 3464 15982
rect 3344 14062 3464 14090
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3148 12368 3200 12374
rect 3148 12310 3200 12316
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1964 11354 1992 11630
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2332 10810 2360 11154
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2320 10668 2372 10674
rect 2424 10656 2452 11018
rect 2372 10628 2452 10656
rect 2320 10610 2372 10616
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2148 10266 2176 10406
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2332 10198 2360 10610
rect 2320 10192 2372 10198
rect 2320 10134 2372 10140
rect 2700 9926 2728 11086
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2792 10130 2820 10542
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1780 8022 1808 9454
rect 2700 9058 2728 9862
rect 2884 9722 2912 10406
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2608 9042 2728 9058
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2596 9036 2728 9042
rect 2648 9030 2728 9036
rect 2596 8978 2648 8984
rect 2240 8498 2268 8978
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 1768 8016 1820 8022
rect 1768 7958 1820 7964
rect 2792 7002 2820 9522
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2976 8090 3004 8366
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2792 2961 2820 6938
rect 3068 3913 3096 9318
rect 3148 9036 3200 9042
rect 3252 9024 3280 10066
rect 3344 9586 3372 14062
rect 3620 12986 3648 19343
rect 3712 18766 3740 19654
rect 3700 18760 3752 18766
rect 3700 18702 3752 18708
rect 3712 18154 3740 18702
rect 3896 18154 3924 22200
rect 3976 21956 4028 21962
rect 3976 21898 4028 21904
rect 3700 18148 3752 18154
rect 3700 18090 3752 18096
rect 3884 18148 3936 18154
rect 3884 18090 3936 18096
rect 3988 17610 4016 21898
rect 4160 20324 4212 20330
rect 4160 20266 4212 20272
rect 4172 20058 4200 20266
rect 4356 20074 4384 22200
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4160 20052 4212 20058
rect 4080 20012 4160 20040
rect 4080 19378 4108 20012
rect 4160 19994 4212 20000
rect 4264 20046 4384 20074
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4172 19310 4200 19654
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4172 17678 4200 18362
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 3976 17604 4028 17610
rect 3976 17546 4028 17552
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4080 16794 4108 17478
rect 4172 17134 4200 17614
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4172 16590 4200 16934
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 4172 14958 4200 16526
rect 4264 15162 4292 20046
rect 4344 19916 4396 19922
rect 4344 19858 4396 19864
rect 4356 19514 4384 19858
rect 4816 19802 4844 22200
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4908 20058 4936 20198
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4816 19774 4936 19802
rect 4804 19712 4856 19718
rect 4804 19654 4856 19660
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4356 18766 4384 19450
rect 4816 19310 4844 19654
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4540 18834 4568 19110
rect 4528 18828 4580 18834
rect 4528 18770 4580 18776
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4816 17354 4844 18090
rect 4908 17882 4936 19774
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 5000 18970 5028 19314
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 4816 17326 4936 17354
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4816 16590 4844 17206
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4816 15570 4844 16526
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 3804 14414 3832 14758
rect 4264 14618 4292 15098
rect 4816 15094 4844 15506
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 4068 14408 4120 14414
rect 4356 14362 4384 14962
rect 4120 14356 4384 14362
rect 4068 14350 4384 14356
rect 4080 14334 4384 14350
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 3792 13796 3844 13802
rect 3792 13738 3844 13744
rect 3804 13326 3832 13738
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 3896 13530 3924 13670
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3792 13320 3844 13326
rect 4724 13297 4752 13670
rect 3792 13262 3844 13268
rect 4710 13288 4766 13297
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3804 12782 3832 13262
rect 4710 13223 4766 13232
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3988 12889 4016 13126
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 3974 12880 4030 12889
rect 3974 12815 4030 12824
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3436 12238 3464 12718
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3528 11937 3556 12378
rect 3804 12238 3832 12718
rect 4066 12336 4122 12345
rect 4172 12306 4200 12922
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4066 12271 4122 12280
rect 4160 12300 4212 12306
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3514 11928 3570 11937
rect 3514 11863 3570 11872
rect 3422 11792 3478 11801
rect 3422 11727 3478 11736
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3436 9489 3464 11727
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3528 10062 3556 10474
rect 3804 10198 3832 12174
rect 4080 11898 4108 12271
rect 4160 12242 4212 12248
rect 4816 12102 4844 12650
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4816 11762 4844 12038
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 3974 11384 4030 11393
rect 4908 11354 4936 17326
rect 3974 11319 4030 11328
rect 4896 11348 4948 11354
rect 3988 11286 4016 11319
rect 4896 11290 4948 11296
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 3974 10976 4030 10985
rect 3974 10911 4030 10920
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3516 10056 3568 10062
rect 3896 10033 3924 10678
rect 3988 10538 4016 10911
rect 3976 10532 4028 10538
rect 3976 10474 4028 10480
rect 4080 10266 4108 11154
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4172 10810 4200 11018
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3516 9998 3568 10004
rect 3882 10024 3938 10033
rect 3528 9586 3556 9998
rect 3882 9959 3938 9968
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3976 9512 4028 9518
rect 3422 9480 3478 9489
rect 3976 9454 4028 9460
rect 3422 9415 3478 9424
rect 3200 8996 3280 9024
rect 3148 8978 3200 8984
rect 3160 8430 3188 8978
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3712 8430 3740 8774
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3804 8276 3832 8774
rect 3712 8248 3832 8276
rect 3054 3904 3110 3913
rect 3054 3839 3110 3848
rect 2778 2952 2834 2961
rect 2778 2887 2834 2896
rect 3712 2553 3740 8248
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3804 3505 3832 7142
rect 3790 3496 3846 3505
rect 3790 3431 3846 3440
rect 3698 2544 3754 2553
rect 3698 2479 3754 2488
rect 3516 2100 3568 2106
rect 3516 2042 3568 2048
rect 3528 2009 3556 2042
rect 3514 2000 3570 2009
rect 3514 1935 3570 1944
rect 3896 1601 3924 8910
rect 3988 8673 4016 9454
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4068 9104 4120 9110
rect 4066 9072 4068 9081
rect 4120 9072 4122 9081
rect 4066 9007 4122 9016
rect 3974 8664 4030 8673
rect 3974 8599 4030 8608
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 7886 4016 8230
rect 4264 8090 4292 9318
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 4172 7546 4200 7890
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4356 7426 4384 11154
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4540 10266 4568 10610
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4816 10062 4844 10950
rect 4908 10810 4936 11290
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 5000 10266 5028 18906
rect 5092 18222 5120 19246
rect 5276 19174 5304 22200
rect 5736 20074 5764 22200
rect 5736 20046 5856 20074
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5460 19514 5488 19790
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5736 18970 5764 19858
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5828 18902 5856 20046
rect 6092 19236 6144 19242
rect 6092 19178 6144 19184
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5092 17338 5120 18158
rect 5184 18154 5212 18770
rect 6104 18766 6132 19178
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 5172 18148 5224 18154
rect 5172 18090 5224 18096
rect 5552 17882 5580 18702
rect 6104 18358 6132 18702
rect 6092 18352 6144 18358
rect 6092 18294 6144 18300
rect 6196 18272 6224 22200
rect 6460 19916 6512 19922
rect 6460 19858 6512 19864
rect 6472 19514 6500 19858
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6472 18698 6500 19450
rect 6460 18692 6512 18698
rect 6460 18634 6512 18640
rect 6552 18352 6604 18358
rect 6552 18294 6604 18300
rect 6196 18244 6316 18272
rect 6184 18148 6236 18154
rect 6184 18090 6236 18096
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 6012 16998 6040 17682
rect 6196 17678 6224 18090
rect 6288 17882 6316 18244
rect 6564 18193 6592 18294
rect 6550 18184 6606 18193
rect 6550 18119 6606 18128
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 6196 16794 6224 17614
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5460 16114 5488 16594
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5368 15706 5396 15846
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5460 15366 5488 16050
rect 6656 15706 6684 22200
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6748 18970 6776 19110
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 5908 15428 5960 15434
rect 5908 15370 5960 15376
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5460 14618 5488 14758
rect 5736 14618 5764 14826
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5920 14074 5948 15370
rect 6288 15162 6316 15506
rect 6656 15162 6684 15642
rect 6276 15156 6328 15162
rect 6644 15156 6696 15162
rect 6328 15116 6500 15144
rect 6276 15098 6328 15104
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6288 14006 6316 14282
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 13530 5488 13738
rect 5736 13530 5764 13806
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5828 12986 5856 13398
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5920 12714 5948 13330
rect 5908 12708 5960 12714
rect 5908 12650 5960 12656
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5460 11762 5488 12242
rect 5920 12102 5948 12650
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 9178 4660 9318
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4816 8566 4844 9522
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 8634 4936 9318
rect 5000 9042 5028 10202
rect 5276 10130 5304 10542
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4804 8560 4856 8566
rect 4804 8502 4856 8508
rect 4434 8120 4490 8129
rect 4434 8055 4436 8064
rect 4488 8055 4490 8064
rect 4436 8026 4488 8032
rect 4816 8022 4844 8502
rect 5552 8362 5580 12038
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5644 11150 5672 11494
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5644 9450 5672 11086
rect 5736 10810 5764 11630
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 6012 11218 6040 11494
rect 6104 11218 6132 12038
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 6196 11082 6224 11630
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6104 9722 6132 10406
rect 6196 10198 6224 11018
rect 6472 10742 6500 15116
rect 6644 15098 6696 15104
rect 6748 15042 6776 18906
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6932 16658 6960 17138
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 15094 6868 15846
rect 6656 15014 6776 15042
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11830 6592 12038
rect 6552 11824 6604 11830
rect 6552 11766 6604 11772
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4816 7426 4844 7958
rect 4264 7398 4384 7426
rect 4724 7410 4844 7426
rect 4712 7404 4844 7410
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3988 6225 4016 6802
rect 3974 6216 4030 6225
rect 3974 6151 4030 6160
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5817 4108 6054
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 3976 5296 4028 5302
rect 4080 5273 4108 5306
rect 3976 5238 4028 5244
rect 4066 5264 4122 5273
rect 3988 4457 4016 5238
rect 4066 5199 4122 5208
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4865 4108 4966
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 3974 4448 4030 4457
rect 3974 4383 4030 4392
rect 3882 1592 3938 1601
rect 3882 1527 3938 1536
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 3344 649 3372 1294
rect 3330 640 3386 649
rect 3330 575 3386 584
rect 4264 241 4292 7398
rect 4764 7398 4844 7404
rect 4712 7346 4764 7352
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 5552 1358 5580 8298
rect 5644 6798 5672 9386
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5736 7886 5764 8230
rect 5828 8090 5856 8230
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 6288 7206 6316 8774
rect 6472 7410 6500 10678
rect 6656 10606 6684 15014
rect 6840 14414 6868 15030
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6840 13870 6868 14350
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6932 13530 6960 14418
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6932 12646 6960 13330
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 7024 12306 7052 18022
rect 7116 14362 7144 22200
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7288 18896 7340 18902
rect 7288 18838 7340 18844
rect 7300 18222 7328 18838
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7208 16794 7236 17614
rect 7392 17610 7420 19246
rect 7576 18086 7604 22200
rect 8036 20346 8064 22200
rect 7668 20318 8064 20346
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 7380 17604 7432 17610
rect 7380 17546 7432 17552
rect 7392 17338 7420 17546
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7668 15722 7696 20318
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7760 18766 7788 19110
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 8220 18970 8248 20198
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 8312 19718 8340 19858
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8312 18902 8340 19654
rect 8300 18896 8352 18902
rect 7930 18864 7986 18873
rect 7840 18828 7892 18834
rect 8300 18838 8352 18844
rect 7930 18799 7932 18808
rect 7840 18770 7892 18776
rect 7984 18799 7986 18808
rect 7932 18770 7984 18776
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7760 17134 7788 18702
rect 7852 18290 7880 18770
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7944 18154 7972 18566
rect 8312 18222 8340 18566
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 7932 18148 7984 18154
rect 7932 18090 7984 18096
rect 8404 18086 8432 18158
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 8220 16658 8248 16934
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8220 16114 8248 16594
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8312 16046 8340 17682
rect 8496 17338 8524 22200
rect 8956 20602 8984 22200
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8772 19990 8800 20402
rect 9416 20058 9444 22200
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 8760 19984 8812 19990
rect 8760 19926 8812 19932
rect 8772 19310 8800 19926
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 8760 19304 8812 19310
rect 8666 19272 8722 19281
rect 8760 19246 8812 19252
rect 8666 19207 8722 19216
rect 8680 18290 8708 19207
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8956 18970 8984 19110
rect 9048 18970 9076 19654
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 9692 18766 9720 19314
rect 9784 19174 9812 19858
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9784 18834 9812 19110
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 9692 17746 9720 18702
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 8668 17604 8720 17610
rect 8668 17546 8720 17552
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 7576 15694 7696 15722
rect 8312 15706 8340 15982
rect 8300 15700 8352 15706
rect 7116 14334 7328 14362
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7116 12782 7144 14214
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7208 13530 7236 14010
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7300 13258 7328 14334
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7392 13394 7420 13738
rect 7576 13462 7604 15694
rect 8300 15642 8352 15648
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7668 14618 7696 15506
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6840 11558 6868 12242
rect 7208 12238 7236 12582
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6932 11286 6960 11562
rect 6920 11280 6972 11286
rect 7012 11280 7064 11286
rect 6920 11222 6972 11228
rect 7010 11248 7012 11257
rect 7064 11248 7066 11257
rect 7010 11183 7066 11192
rect 7300 11150 7328 11562
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6656 10146 6684 10542
rect 6748 10266 6776 10610
rect 6828 10600 6880 10606
rect 6880 10560 6960 10588
rect 6828 10542 6880 10548
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6656 10118 6868 10146
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6380 7002 6408 7142
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 1352 5592 1358
rect 5540 1294 5592 1300
rect 6472 1057 6500 7346
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6748 6798 6776 7210
rect 6840 7177 6868 10118
rect 6932 9586 6960 10560
rect 7392 10554 7420 13330
rect 7668 12374 7696 14554
rect 8404 14482 8432 16390
rect 8496 15978 8524 17274
rect 8680 16114 8708 17546
rect 8956 17270 8984 17682
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 9048 17338 9076 17614
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 8944 17264 8996 17270
rect 8944 17206 8996 17212
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8864 16658 8892 17070
rect 9324 16794 9352 17478
rect 9876 17134 9904 22200
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10048 19780 10100 19786
rect 10048 19722 10100 19728
rect 10060 19242 10088 19722
rect 10152 19514 10180 19790
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10048 19236 10100 19242
rect 10048 19178 10100 19184
rect 10060 18970 10088 19178
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9968 17542 9996 18770
rect 10048 17808 10100 17814
rect 10048 17750 10100 17756
rect 10140 17808 10192 17814
rect 10140 17750 10192 17756
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 10060 17202 10088 17750
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9508 16658 9536 16934
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8680 14958 8708 16050
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8036 14074 8064 14214
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8220 13870 8248 14214
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 8220 13326 8248 13806
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7484 11218 7512 11494
rect 7564 11348 7616 11354
rect 7760 11336 7788 12650
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8496 11898 8524 12310
rect 8772 12306 8800 13806
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 7616 11308 7788 11336
rect 7564 11290 7616 11296
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 8024 11212 8076 11218
rect 8404 11200 8432 11494
rect 8496 11286 8524 11562
rect 8484 11280 8536 11286
rect 8576 11280 8628 11286
rect 8484 11222 8536 11228
rect 8574 11248 8576 11257
rect 8628 11248 8630 11257
rect 8076 11172 8432 11200
rect 8574 11183 8630 11192
rect 8024 11154 8076 11160
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 8128 10810 8156 11018
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 7300 10526 7420 10554
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7300 9382 7328 10526
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7392 10266 7420 10406
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7668 9518 7696 10542
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 8220 10062 8248 10406
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 7944 9586 7972 9998
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 8838 7328 9318
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7392 8430 7420 9454
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8404 9178 8432 11172
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8496 10606 8524 11018
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8864 10062 8892 16594
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9048 16250 9076 16526
rect 10060 16250 10088 17138
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8956 11354 8984 12582
rect 9048 12374 9076 12786
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 9232 11801 9260 15982
rect 9404 15972 9456 15978
rect 9404 15914 9456 15920
rect 9416 15502 9444 15914
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9416 15162 9444 15438
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9692 14618 9720 15370
rect 9956 14884 10008 14890
rect 9956 14826 10008 14832
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9968 14006 9996 14826
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 9324 12442 9352 13194
rect 9508 12850 9536 13330
rect 9600 13258 9628 13738
rect 9968 13326 9996 13942
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 10060 12782 10088 13330
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9218 11792 9274 11801
rect 9508 11762 9536 12242
rect 9218 11727 9274 11736
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9508 11354 9536 11698
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10810 9260 10950
rect 9416 10810 9444 11018
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9508 10674 9536 11290
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9586 10568 9642 10577
rect 8944 10532 8996 10538
rect 9586 10503 9642 10512
rect 8944 10474 8996 10480
rect 8956 10062 8984 10474
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7116 8090 7144 8298
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7392 7954 7420 8366
rect 7668 8294 7696 8910
rect 8036 8634 8064 8978
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 7954 7696 8230
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 6826 7168 6882 7177
rect 6826 7103 6882 7112
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6840 2106 6868 7103
rect 7116 7002 7144 7414
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 7668 6798 7696 7890
rect 8220 7546 8248 9114
rect 8404 8430 8432 9114
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8496 8090 8524 8774
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 7840 7336 7892 7342
rect 7838 7304 7840 7313
rect 7892 7304 7894 7313
rect 7838 7239 7894 7248
rect 7748 7200 7800 7206
rect 7746 7168 7748 7177
rect 7800 7168 7802 7177
rect 7746 7103 7802 7112
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 8496 6662 8524 7890
rect 8680 7818 8708 9386
rect 8864 8906 8892 9998
rect 8956 9722 8984 9998
rect 9600 9926 9628 10503
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 9784 9586 9812 11630
rect 10060 10266 10088 12718
rect 10152 11626 10180 17750
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10244 16182 10272 16730
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10336 15706 10364 22200
rect 10508 18896 10560 18902
rect 10508 18838 10560 18844
rect 10416 18352 10468 18358
rect 10416 18294 10468 18300
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10244 14958 10272 15438
rect 10336 15162 10364 15642
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 10244 14822 10272 14894
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10428 13734 10456 18294
rect 10520 14958 10548 18838
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10612 15978 10640 16594
rect 10600 15972 10652 15978
rect 10600 15914 10652 15920
rect 10508 14952 10560 14958
rect 10508 14894 10560 14900
rect 10520 14618 10548 14894
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10612 13190 10640 15914
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10704 15706 10732 15846
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10796 13530 10824 22200
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10888 14550 10916 18022
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10980 15570 11008 16594
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 11072 15450 11100 20198
rect 11256 19394 11284 22200
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11716 20074 11744 22200
rect 12176 20262 12204 22200
rect 12636 20482 12664 22200
rect 12636 20454 13032 20482
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 11716 20046 12204 20074
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11256 19366 11928 19394
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11164 16114 11192 16730
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11164 15638 11192 16050
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11072 15422 11192 15450
rect 10876 14544 10928 14550
rect 10876 14486 10928 14492
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10140 11620 10192 11626
rect 10140 11562 10192 11568
rect 10336 11354 10364 12242
rect 11072 12186 11100 12582
rect 11164 12374 11192 15422
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 10416 12164 10468 12170
rect 11072 12158 11192 12186
rect 10416 12106 10468 12112
rect 10428 11694 10456 12106
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11072 11694 11100 12038
rect 11164 11898 11192 12158
rect 11256 11898 11284 19246
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11900 17814 11928 19366
rect 11992 17882 12020 19858
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11716 16250 11744 17682
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11808 17338 11836 17614
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11900 15910 11928 17070
rect 11992 16658 12020 17274
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11900 14278 11928 15846
rect 12084 15094 12112 18158
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 11888 14272 11940 14278
rect 11940 14220 12020 14226
rect 11888 14214 12020 14220
rect 11900 14198 12020 14214
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11716 12986 11744 13670
rect 11900 13530 11928 13874
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11900 12646 11928 12718
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11900 12442 11928 12582
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11808 12186 11836 12310
rect 11992 12306 12020 14198
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11808 12158 11928 12186
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11808 11762 11836 12038
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10888 10713 10916 10746
rect 10874 10704 10930 10713
rect 10874 10639 10930 10648
rect 11072 10538 11100 11494
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11256 10810 11284 11154
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9876 9994 9904 10202
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 10060 9722 10088 10202
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10704 9586 10732 10066
rect 11256 9994 11284 10746
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 11244 9988 11296 9994
rect 11244 9930 11296 9936
rect 11164 9654 11192 9930
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11152 9648 11204 9654
rect 11150 9616 11152 9625
rect 11204 9616 11206 9625
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 10692 9580 10744 9586
rect 11150 9551 11206 9560
rect 10692 9522 10744 9528
rect 11164 9525 11192 9551
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 11164 8566 11192 9318
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11900 8634 11928 12158
rect 11992 10266 12020 12242
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8772 8022 8800 8434
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8772 7410 8800 7958
rect 8864 7857 8892 7958
rect 8850 7848 8906 7857
rect 8850 7783 8906 7792
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8574 6760 8630 6769
rect 8574 6695 8630 6704
rect 8588 6662 8616 6695
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 12084 4826 12112 14826
rect 12176 12458 12204 20046
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12268 17338 12296 18158
rect 12360 17814 12388 18226
rect 12452 17882 12480 18362
rect 12544 18222 12572 18770
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12348 17808 12400 17814
rect 12348 17750 12400 17756
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12268 12646 12296 17138
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12360 16794 12388 17070
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12452 15366 12480 17614
rect 12544 17202 12572 17750
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12544 16250 12572 17002
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12452 14550 12480 15302
rect 12544 15162 12572 15846
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12440 14544 12492 14550
rect 12440 14486 12492 14492
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12360 12986 12388 13806
rect 12452 13190 12480 13806
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12530 12472 12586 12481
rect 12176 12430 12296 12458
rect 12268 12356 12296 12430
rect 12530 12407 12586 12416
rect 12268 12328 12388 12356
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12176 10198 12204 11086
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 12268 10130 12296 10406
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12360 9659 12388 12328
rect 12544 11762 12572 12407
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12452 11286 12480 11494
rect 12636 11354 12664 19246
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12728 17202 12756 18566
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12728 16726 12756 17138
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12728 16114 12756 16662
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12820 14074 12848 20334
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12912 18358 12940 18702
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12912 14906 12940 17818
rect 13004 16674 13032 20454
rect 13096 19174 13124 22200
rect 13556 20058 13584 22200
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 14016 19786 14044 22200
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 14004 19780 14056 19786
rect 14004 19722 14056 19728
rect 14108 19446 14136 20334
rect 14476 20058 14504 22200
rect 14936 20602 14964 22200
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 14556 20324 14608 20330
rect 14556 20266 14608 20272
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14568 19922 14596 20266
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 15396 20058 15424 22200
rect 15856 20058 15884 22200
rect 16316 20058 16344 22200
rect 16776 20058 16804 22200
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14096 19440 14148 19446
rect 14096 19382 14148 19388
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 13174 18728 13230 18737
rect 13174 18663 13230 18672
rect 13188 17542 13216 18663
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13188 16998 13216 17478
rect 13176 16992 13228 16998
rect 13176 16934 13228 16940
rect 13372 16794 13400 19246
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13556 17882 13584 18770
rect 14200 18698 14228 19790
rect 14660 19242 14688 19858
rect 15396 19310 15424 19858
rect 16408 19378 16436 19858
rect 16960 19378 16988 19858
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 14648 19236 14700 19242
rect 14648 19178 14700 19184
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14280 18896 14332 18902
rect 14660 18850 14688 18906
rect 14280 18838 14332 18844
rect 14188 18692 14240 18698
rect 14188 18634 14240 18640
rect 14292 18426 14320 18838
rect 14568 18822 14688 18850
rect 14568 18630 14596 18822
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 13648 17082 13676 18362
rect 14568 17882 14596 18566
rect 14660 18426 14688 18702
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14556 17876 14608 17882
rect 14476 17836 14556 17864
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13556 17054 13676 17082
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13004 16646 13400 16674
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 12912 14878 13032 14906
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 12306 12756 13126
rect 12912 12782 12940 14758
rect 13004 13326 13032 14878
rect 13280 14618 13308 15506
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 13004 12850 13032 13126
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12820 12481 12848 12650
rect 12806 12472 12862 12481
rect 12806 12407 12862 12416
rect 13096 12374 13124 13466
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12728 11558 12756 12242
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12452 10606 12480 11222
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12452 10470 12480 10542
rect 12544 10538 12572 11154
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12728 10606 12756 11018
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12346 9650 12402 9659
rect 12346 9585 12402 9594
rect 13372 9382 13400 16646
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13464 15366 13492 15914
rect 13556 15910 13584 17054
rect 13636 16040 13688 16046
rect 13740 16028 13768 17138
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 14016 16794 14044 17002
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 13688 16000 13768 16028
rect 13636 15982 13688 15988
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13556 14618 13584 14962
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13648 14482 13676 15982
rect 13924 15162 13952 16662
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 14016 15706 14044 16594
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 14108 15434 14136 17070
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14200 16590 14228 16934
rect 14292 16658 14320 17478
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14292 16402 14320 16594
rect 14200 16374 14320 16402
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 14200 15042 14228 16374
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 13832 15014 14228 15042
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13464 13394 13492 13942
rect 13740 13870 13768 14554
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13464 12850 13492 13330
rect 13740 13326 13768 13806
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13556 12986 13584 13262
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13464 11218 13492 11494
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13464 10130 13492 11154
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13556 10062 13584 12922
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13648 11354 13676 12174
rect 13832 11898 13860 15014
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14200 14074 14228 14894
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13832 11354 13860 11834
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 14016 11014 14044 13126
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 14108 9926 14136 13194
rect 14292 12782 14320 15506
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14384 14958 14412 15438
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 13870 14412 14214
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14476 13530 14504 17836
rect 14556 17818 14608 17824
rect 14648 17060 14700 17066
rect 14648 17002 14700 17008
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14568 15638 14596 16390
rect 14660 16250 14688 17002
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14556 15632 14608 15638
rect 14556 15574 14608 15580
rect 14660 15502 14688 16186
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14660 15026 14688 15438
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14568 13734 14596 14214
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14476 12986 14504 13466
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14200 11762 14228 12106
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14292 11694 14320 12582
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14476 11354 14504 12242
rect 14568 12186 14596 13670
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14660 12306 14688 12718
rect 14752 12442 14780 19246
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 15304 18290 15332 18566
rect 15396 18426 15424 18634
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15488 18222 15516 18566
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15292 18148 15344 18154
rect 15292 18090 15344 18096
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15120 17066 15148 17682
rect 15304 17678 15332 18090
rect 15764 17814 15792 18702
rect 15752 17808 15804 17814
rect 15752 17750 15804 17756
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 15304 16658 15332 17614
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15212 15978 15240 16526
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15672 16114 15700 16390
rect 16040 16114 16068 16526
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15200 15972 15252 15978
rect 15200 15914 15252 15920
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15304 15706 15332 15846
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15396 15434 15424 15982
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15488 15450 15516 15914
rect 15488 15434 15608 15450
rect 15384 15428 15436 15434
rect 15384 15370 15436 15376
rect 15488 15428 15620 15434
rect 15488 15422 15568 15428
rect 15488 15162 15516 15422
rect 15568 15370 15620 15376
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15672 15094 15700 16050
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 15672 13938 15700 15030
rect 15856 14890 15884 15438
rect 16040 14958 16068 16050
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15948 14482 15976 14894
rect 15844 14476 15896 14482
rect 15844 14418 15896 14424
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15856 13938 15884 14418
rect 16040 14006 16068 14894
rect 16316 14074 16344 19246
rect 16580 19236 16632 19242
rect 16580 19178 16632 19184
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 15292 13728 15344 13734
rect 15212 13676 15292 13682
rect 15212 13670 15344 13676
rect 15212 13654 15332 13670
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 15212 13410 15240 13654
rect 15120 13382 15240 13410
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14936 12714 14964 13194
rect 15120 13190 15148 13382
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 15856 12374 15884 13262
rect 16408 12986 16436 13874
rect 16592 12986 16620 19178
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16684 18154 16712 18634
rect 16672 18148 16724 18154
rect 16672 18090 16724 18096
rect 16684 17882 16712 18090
rect 16672 17876 16724 17882
rect 16672 17818 16724 17824
rect 16672 17536 16724 17542
rect 16776 17524 16804 18702
rect 16724 17496 16804 17524
rect 16672 17478 16724 17484
rect 16684 15502 16712 17478
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16776 15502 16804 16662
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16776 15178 16804 15438
rect 16776 15162 16896 15178
rect 16776 15156 16908 15162
rect 16776 15150 16856 15156
rect 16856 15098 16908 15104
rect 16960 15042 16988 18770
rect 17052 17338 17080 19246
rect 17236 18970 17264 22200
rect 17696 19786 17724 22200
rect 18156 20482 18184 22200
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18064 20454 18184 20482
rect 17684 19780 17736 19786
rect 17684 19722 17736 19728
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17144 18714 17172 18906
rect 17144 18686 17264 18714
rect 17236 18086 17264 18686
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 16868 15014 16988 15042
rect 17236 15026 17264 18022
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17328 16114 17356 16934
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17224 15020 17276 15026
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16684 14618 16712 14826
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16684 13938 16712 14554
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16776 12442 16804 12650
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 15200 12232 15252 12238
rect 14568 12158 14688 12186
rect 15200 12174 15252 12180
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14384 10810 14412 11086
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14384 10606 14412 10746
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 14660 5302 14688 12158
rect 15212 11626 15240 12174
rect 15856 11898 15884 12310
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15488 10810 15516 11562
rect 16120 11280 16172 11286
rect 16120 11222 16172 11228
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 14752 8090 14780 10066
rect 16132 10062 16160 11222
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16316 10674 16344 11154
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16868 10266 16896 15014
rect 17224 14962 17276 14968
rect 17236 14822 17264 14962
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16960 13870 16988 14350
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17052 12782 17080 13262
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17144 12850 17172 13126
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 17052 10606 17080 10950
rect 17040 10600 17092 10606
rect 17092 10548 17172 10554
rect 17040 10542 17172 10548
rect 17052 10526 17172 10542
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 17144 10062 17172 10526
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 15120 9722 15148 9998
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 17328 9110 17356 15846
rect 17420 15706 17448 16934
rect 17788 16794 17816 17138
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17420 9518 17448 14758
rect 17972 14074 18000 19246
rect 18064 19174 18092 20454
rect 18616 20058 18644 22200
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18880 19984 18932 19990
rect 18880 19926 18932 19932
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18156 18290 18184 19858
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18236 19236 18288 19242
rect 18236 19178 18288 19184
rect 18248 18834 18276 19178
rect 18236 18828 18288 18834
rect 18236 18770 18288 18776
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18064 17882 18092 18158
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18064 16250 18092 17614
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18156 16658 18184 17070
rect 18604 17060 18656 17066
rect 18604 17002 18656 17008
rect 18616 16794 18644 17002
rect 18800 16998 18828 17614
rect 18788 16992 18840 16998
rect 18788 16934 18840 16940
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18144 16652 18196 16658
rect 18144 16594 18196 16600
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 18156 16182 18184 16594
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18144 16176 18196 16182
rect 18144 16118 18196 16124
rect 18156 15570 18184 16118
rect 18616 16114 18644 16730
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18144 15564 18196 15570
rect 18144 15506 18196 15512
rect 18524 15434 18552 15846
rect 18800 15638 18828 16934
rect 18788 15632 18840 15638
rect 18788 15574 18840 15580
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18512 15428 18564 15434
rect 18512 15370 18564 15376
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18616 14958 18644 15506
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18064 13938 18092 14758
rect 18616 14498 18644 14894
rect 18524 14482 18644 14498
rect 18512 14476 18644 14482
rect 18564 14470 18644 14476
rect 18512 14418 18564 14424
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18708 13938 18736 14214
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18708 13462 18736 13874
rect 18696 13456 18748 13462
rect 18696 13398 18748 13404
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17696 12850 17724 13194
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17788 12374 17816 13262
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18892 12986 18920 19926
rect 19076 18970 19104 22200
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19260 14006 19288 18158
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19352 14550 19380 14962
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 19168 12850 19196 13126
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17604 11830 17632 12310
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17512 8294 17540 11494
rect 17604 11218 17632 11766
rect 18064 11762 18092 12242
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 18156 11286 18184 12038
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18708 11762 18736 12786
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18800 12102 18828 12718
rect 19260 12646 19288 13942
rect 19352 13802 19380 14350
rect 19340 13796 19392 13802
rect 19340 13738 19392 13744
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19260 12442 19288 12582
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18892 11694 18920 12174
rect 19444 11898 19472 12582
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 17684 10736 17736 10742
rect 17682 10704 17684 10713
rect 17736 10704 17738 10713
rect 17682 10639 17738 10648
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18064 10266 18092 10406
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 19536 7478 19564 22200
rect 19996 17354 20024 22200
rect 19720 17326 20024 17354
rect 19720 7546 19748 17326
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19904 15026 19932 15302
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19524 7472 19576 7478
rect 19524 7414 19576 7420
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 18800 6662 18828 7278
rect 20456 6730 20484 22200
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20732 18970 20760 19246
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 20916 6458 20944 22200
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21192 18154 21220 19178
rect 21180 18148 21232 18154
rect 21180 18090 21232 18096
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20456 5574 20484 5714
rect 20444 5568 20496 5574
rect 20444 5510 20496 5516
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 20456 5370 20484 5510
rect 21008 5370 21036 18022
rect 21376 17354 21404 22200
rect 21836 18086 21864 22200
rect 22296 18970 22324 22200
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22756 18222 22784 22200
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21100 17326 21404 17354
rect 21100 5914 21128 17326
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 21376 14278 21404 14894
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21376 11529 21404 14214
rect 21362 11520 21418 11529
rect 21362 11455 21418 11464
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 20996 5364 21048 5370
rect 20996 5306 21048 5312
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 6828 2100 6880 2106
rect 6828 2042 6880 2048
rect 11716 1986 11744 4762
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 11532 1958 11744 1986
rect 6458 1048 6514 1057
rect 6458 983 6514 992
rect 11532 800 11560 1958
rect 4250 232 4306 241
rect 4250 167 4306 176
rect 11518 0 11574 800
<< via2 >>
rect 2870 22208 2926 22264
rect 202 19080 258 19136
rect 1950 21256 2006 21312
rect 1582 20712 1638 20768
rect 1490 19760 1546 19816
rect 1122 18672 1178 18728
rect 1398 14184 1454 14240
rect 3238 22616 3294 22672
rect 2778 21664 2834 21720
rect 2594 19116 2596 19136
rect 2596 19116 2648 19136
rect 2648 19116 2650 19136
rect 2594 19080 2650 19116
rect 1766 18400 1822 18456
rect 1858 18164 1860 18184
rect 1860 18164 1912 18184
rect 1912 18164 1914 18184
rect 1858 18128 1914 18164
rect 2778 18808 2834 18864
rect 2502 18028 2504 18048
rect 2504 18028 2556 18048
rect 2556 18028 2558 18048
rect 2502 17992 2558 18028
rect 1950 17448 2006 17504
rect 1674 17040 1730 17096
rect 1674 16496 1730 16552
rect 1674 16088 1730 16144
rect 3054 20304 3110 20360
rect 3606 19352 3662 19408
rect 3422 19080 3478 19136
rect 3514 18808 3570 18864
rect 3238 15544 3294 15600
rect 1858 14592 1914 14648
rect 1950 13776 2006 13832
rect 3054 15136 3110 15192
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4710 13232 4766 13288
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 3974 12824 4030 12880
rect 4066 12280 4122 12336
rect 3514 11872 3570 11928
rect 3422 11736 3478 11792
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 3974 11328 4030 11384
rect 3974 10920 4030 10976
rect 3882 9968 3938 10024
rect 3422 9424 3478 9480
rect 3054 3848 3110 3904
rect 2778 2896 2834 2952
rect 3790 3440 3846 3496
rect 3698 2488 3754 2544
rect 3514 1944 3570 2000
rect 4066 9052 4068 9072
rect 4068 9052 4120 9072
rect 4120 9052 4122 9072
rect 4066 9016 4122 9052
rect 3974 8608 4030 8664
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 6550 18128 6606 18184
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4434 8084 4490 8120
rect 4434 8064 4436 8084
rect 4436 8064 4488 8084
rect 4488 8064 4490 8084
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 3974 6160 4030 6216
rect 4066 5752 4122 5808
rect 4066 5208 4122 5264
rect 4066 4800 4122 4856
rect 3974 4392 4030 4448
rect 3882 1536 3938 1592
rect 3330 584 3386 640
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7930 18828 7986 18864
rect 7930 18808 7932 18828
rect 7932 18808 7984 18828
rect 7984 18808 7986 18828
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 8666 19216 8722 19272
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7010 11228 7012 11248
rect 7012 11228 7064 11248
rect 7064 11228 7066 11248
rect 7010 11192 7066 11228
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 8574 11228 8576 11248
rect 8576 11228 8628 11248
rect 8628 11228 8630 11248
rect 8574 11192 8630 11228
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 9218 11736 9274 11792
rect 9586 10512 9642 10568
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 6826 7112 6882 7168
rect 7838 7284 7840 7304
rect 7840 7284 7892 7304
rect 7892 7284 7894 7304
rect 7838 7248 7894 7284
rect 7746 7148 7748 7168
rect 7748 7148 7800 7168
rect 7800 7148 7802 7168
rect 7746 7112 7802 7148
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 10874 10648 10930 10704
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11150 9596 11152 9616
rect 11152 9596 11204 9616
rect 11204 9596 11206 9616
rect 11150 9560 11206 9596
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 8850 7792 8906 7848
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 8574 6704 8630 6760
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 12530 12416 12586 12472
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 13174 18672 13230 18728
rect 12806 12416 12862 12472
rect 12346 9594 12402 9650
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 17682 10684 17684 10704
rect 17684 10684 17736 10704
rect 17736 10684 17738 10704
rect 17682 10648 17738 10684
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 21362 11464 21418 11520
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 6458 992 6514 1048
rect 4250 176 4306 232
<< metal3 >>
rect 0 22674 800 22704
rect 3233 22674 3299 22677
rect 0 22672 3299 22674
rect 0 22616 3238 22672
rect 3294 22616 3299 22672
rect 0 22614 3299 22616
rect 0 22584 800 22614
rect 3233 22611 3299 22614
rect 0 22266 800 22296
rect 2865 22266 2931 22269
rect 0 22264 2931 22266
rect 0 22208 2870 22264
rect 2926 22208 2931 22264
rect 0 22206 2931 22208
rect 0 22176 800 22206
rect 2865 22203 2931 22206
rect 0 21722 800 21752
rect 2773 21722 2839 21725
rect 0 21720 2839 21722
rect 0 21664 2778 21720
rect 2834 21664 2839 21720
rect 0 21662 2839 21664
rect 0 21632 800 21662
rect 2773 21659 2839 21662
rect 0 21314 800 21344
rect 1945 21314 2011 21317
rect 0 21312 2011 21314
rect 0 21256 1950 21312
rect 2006 21256 2011 21312
rect 0 21254 2011 21256
rect 0 21224 800 21254
rect 1945 21251 2011 21254
rect 0 20770 800 20800
rect 1577 20770 1643 20773
rect 0 20768 1643 20770
rect 0 20712 1582 20768
rect 1638 20712 1643 20768
rect 0 20710 1643 20712
rect 0 20680 800 20710
rect 1577 20707 1643 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 0 20362 800 20392
rect 3049 20362 3115 20365
rect 0 20360 3115 20362
rect 0 20304 3054 20360
rect 3110 20304 3115 20360
rect 0 20302 3115 20304
rect 0 20272 800 20302
rect 3049 20299 3115 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 0 19818 800 19848
rect 1485 19818 1551 19821
rect 0 19816 1551 19818
rect 0 19760 1490 19816
rect 1546 19760 1551 19816
rect 0 19758 1551 19760
rect 0 19728 800 19758
rect 1485 19755 1551 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 0 19410 800 19440
rect 3601 19410 3667 19413
rect 0 19408 3667 19410
rect 0 19352 3606 19408
rect 3662 19352 3667 19408
rect 0 19350 3667 19352
rect 0 19320 800 19350
rect 3601 19347 3667 19350
rect 8661 19274 8727 19277
rect 982 19272 8727 19274
rect 982 19216 8666 19272
rect 8722 19216 8727 19272
rect 982 19214 8727 19216
rect 197 19138 263 19141
rect 982 19138 1042 19214
rect 8661 19211 8727 19214
rect 197 19136 1042 19138
rect 197 19080 202 19136
rect 258 19080 1042 19136
rect 197 19078 1042 19080
rect 2589 19138 2655 19141
rect 3417 19138 3483 19141
rect 2589 19136 3483 19138
rect 2589 19080 2594 19136
rect 2650 19080 3422 19136
rect 3478 19080 3483 19136
rect 2589 19078 3483 19080
rect 197 19075 263 19078
rect 2589 19075 2655 19078
rect 3417 19075 3483 19078
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 0 18866 800 18896
rect 2773 18866 2839 18869
rect 0 18864 2839 18866
rect 0 18808 2778 18864
rect 2834 18808 2839 18864
rect 0 18806 2839 18808
rect 0 18776 800 18806
rect 2773 18803 2839 18806
rect 3509 18866 3575 18869
rect 7925 18866 7991 18869
rect 3509 18864 7991 18866
rect 3509 18808 3514 18864
rect 3570 18808 7930 18864
rect 7986 18808 7991 18864
rect 3509 18806 7991 18808
rect 3509 18803 3575 18806
rect 7925 18803 7991 18806
rect 1117 18730 1183 18733
rect 13169 18730 13235 18733
rect 1117 18728 13235 18730
rect 1117 18672 1122 18728
rect 1178 18672 13174 18728
rect 13230 18672 13235 18728
rect 1117 18670 13235 18672
rect 1117 18667 1183 18670
rect 13169 18667 13235 18670
rect 4409 18528 4729 18529
rect 0 18458 800 18488
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 1761 18458 1827 18461
rect 0 18456 1827 18458
rect 0 18400 1766 18456
rect 1822 18400 1827 18456
rect 0 18398 1827 18400
rect 0 18368 800 18398
rect 1761 18395 1827 18398
rect 1853 18186 1919 18189
rect 6545 18186 6611 18189
rect 1853 18184 6611 18186
rect 1853 18128 1858 18184
rect 1914 18128 6550 18184
rect 6606 18128 6611 18184
rect 1853 18126 6611 18128
rect 1853 18123 1919 18126
rect 6545 18123 6611 18126
rect 0 18050 800 18080
rect 2497 18050 2563 18053
rect 0 18048 2563 18050
rect 0 17992 2502 18048
rect 2558 17992 2563 18048
rect 0 17990 2563 17992
rect 0 17960 800 17990
rect 2497 17987 2563 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 17919 15125 17920
rect 0 17506 800 17536
rect 1945 17506 2011 17509
rect 0 17504 2011 17506
rect 0 17448 1950 17504
rect 2006 17448 2011 17504
rect 0 17446 2011 17448
rect 0 17416 800 17446
rect 1945 17443 2011 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 0 17098 800 17128
rect 1669 17098 1735 17101
rect 0 17096 1735 17098
rect 0 17040 1674 17096
rect 1730 17040 1735 17096
rect 0 17038 1735 17040
rect 0 17008 800 17038
rect 1669 17035 1735 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 0 16554 800 16584
rect 1669 16554 1735 16557
rect 0 16552 1735 16554
rect 0 16496 1674 16552
rect 1730 16496 1735 16552
rect 0 16494 1735 16496
rect 0 16464 800 16494
rect 1669 16491 1735 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16146 800 16176
rect 1669 16146 1735 16149
rect 0 16144 1735 16146
rect 0 16088 1674 16144
rect 1730 16088 1735 16144
rect 0 16086 1735 16088
rect 0 16056 800 16086
rect 1669 16083 1735 16086
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 0 15602 800 15632
rect 3233 15602 3299 15605
rect 0 15600 3299 15602
rect 0 15544 3238 15600
rect 3294 15544 3299 15600
rect 0 15542 3299 15544
rect 0 15512 800 15542
rect 3233 15539 3299 15542
rect 4409 15264 4729 15265
rect 0 15194 800 15224
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 3049 15194 3115 15197
rect 0 15192 3115 15194
rect 0 15136 3054 15192
rect 3110 15136 3115 15192
rect 0 15134 3115 15136
rect 0 15104 800 15134
rect 3049 15131 3115 15134
rect 7874 14720 8194 14721
rect 0 14650 800 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 1853 14650 1919 14653
rect 0 14648 1919 14650
rect 0 14592 1858 14648
rect 1914 14592 1919 14648
rect 0 14590 1919 14592
rect 0 14560 800 14590
rect 1853 14587 1919 14590
rect 0 14242 800 14272
rect 1393 14242 1459 14245
rect 0 14240 1459 14242
rect 0 14184 1398 14240
rect 1454 14184 1459 14240
rect 0 14182 1459 14184
rect 0 14152 800 14182
rect 1393 14179 1459 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 0 13834 800 13864
rect 1945 13834 2011 13837
rect 0 13832 2011 13834
rect 0 13776 1950 13832
rect 2006 13776 2011 13832
rect 0 13774 2011 13776
rect 0 13744 800 13774
rect 1945 13771 2011 13774
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 0 13290 800 13320
rect 4705 13290 4771 13293
rect 0 13288 4771 13290
rect 0 13232 4710 13288
rect 4766 13232 4771 13288
rect 0 13230 4771 13232
rect 0 13200 800 13230
rect 4705 13227 4771 13230
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 0 12882 800 12912
rect 3969 12882 4035 12885
rect 0 12880 4035 12882
rect 0 12824 3974 12880
rect 4030 12824 4035 12880
rect 0 12822 4035 12824
rect 0 12792 800 12822
rect 3969 12819 4035 12822
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 12525 12474 12591 12477
rect 12801 12474 12867 12477
rect 12525 12472 12867 12474
rect 12525 12416 12530 12472
rect 12586 12416 12806 12472
rect 12862 12416 12867 12472
rect 12525 12414 12867 12416
rect 12525 12411 12591 12414
rect 12801 12411 12867 12414
rect 0 12338 800 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 800 12278
rect 4061 12275 4127 12278
rect 4409 12000 4729 12001
rect 0 11930 800 11960
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 3509 11930 3575 11933
rect 0 11928 3575 11930
rect 0 11872 3514 11928
rect 3570 11872 3575 11928
rect 0 11870 3575 11872
rect 0 11840 800 11870
rect 3509 11867 3575 11870
rect 3417 11794 3483 11797
rect 9213 11794 9279 11797
rect 3417 11792 9279 11794
rect 3417 11736 3422 11792
rect 3478 11736 9218 11792
rect 9274 11736 9279 11792
rect 3417 11734 9279 11736
rect 3417 11731 3483 11734
rect 9213 11731 9279 11734
rect 21357 11522 21423 11525
rect 22200 11522 23000 11552
rect 21357 11520 23000 11522
rect 21357 11464 21362 11520
rect 21418 11464 23000 11520
rect 21357 11462 23000 11464
rect 21357 11459 21423 11462
rect 7874 11456 8194 11457
rect 0 11386 800 11416
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 22200 11432 23000 11462
rect 14805 11391 15125 11392
rect 3969 11386 4035 11389
rect 0 11384 4035 11386
rect 0 11328 3974 11384
rect 4030 11328 4035 11384
rect 0 11326 4035 11328
rect 0 11296 800 11326
rect 3969 11323 4035 11326
rect 7005 11250 7071 11253
rect 8569 11250 8635 11253
rect 7005 11248 8635 11250
rect 7005 11192 7010 11248
rect 7066 11192 8574 11248
rect 8630 11192 8635 11248
rect 7005 11190 8635 11192
rect 7005 11187 7071 11190
rect 8569 11187 8635 11190
rect 0 10978 800 11008
rect 3969 10978 4035 10981
rect 0 10976 4035 10978
rect 0 10920 3974 10976
rect 4030 10920 4035 10976
rect 0 10918 4035 10920
rect 0 10888 800 10918
rect 3969 10915 4035 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 10869 10706 10935 10709
rect 17677 10706 17743 10709
rect 10869 10704 17743 10706
rect 10869 10648 10874 10704
rect 10930 10648 17682 10704
rect 17738 10648 17743 10704
rect 10869 10646 17743 10648
rect 10869 10643 10935 10646
rect 17677 10643 17743 10646
rect 9581 10570 9647 10573
rect 4846 10568 9647 10570
rect 4846 10512 9586 10568
rect 9642 10512 9647 10568
rect 4846 10510 9647 10512
rect 0 10434 800 10464
rect 4846 10434 4906 10510
rect 9581 10507 9647 10510
rect 0 10374 4906 10434
rect 0 10344 800 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 0 10026 800 10056
rect 3877 10026 3943 10029
rect 0 10024 3943 10026
rect 0 9968 3882 10024
rect 3938 9968 3943 10024
rect 0 9966 3943 9968
rect 0 9936 800 9966
rect 3877 9963 3943 9966
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 12341 9652 12407 9655
rect 12206 9650 12407 9652
rect 11145 9618 11211 9621
rect 12206 9618 12346 9650
rect 11145 9616 12346 9618
rect 11145 9560 11150 9616
rect 11206 9594 12346 9616
rect 12402 9594 12407 9650
rect 11206 9592 12407 9594
rect 11206 9560 12266 9592
rect 12341 9589 12407 9592
rect 11145 9558 12266 9560
rect 11145 9555 11211 9558
rect 0 9482 800 9512
rect 3417 9482 3483 9485
rect 0 9480 3483 9482
rect 0 9424 3422 9480
rect 3478 9424 3483 9480
rect 0 9422 3483 9424
rect 0 9392 800 9422
rect 3417 9419 3483 9422
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 0 9074 800 9104
rect 4061 9074 4127 9077
rect 0 9072 4127 9074
rect 0 9016 4066 9072
rect 4122 9016 4127 9072
rect 0 9014 4127 9016
rect 0 8984 800 9014
rect 4061 9011 4127 9014
rect 4409 8736 4729 8737
rect 0 8666 800 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 3969 8666 4035 8669
rect 0 8664 4035 8666
rect 0 8608 3974 8664
rect 4030 8608 4035 8664
rect 0 8606 4035 8608
rect 0 8576 800 8606
rect 3969 8603 4035 8606
rect 7874 8192 8194 8193
rect 0 8122 800 8152
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 4429 8122 4495 8125
rect 0 8120 4495 8122
rect 0 8064 4434 8120
rect 4490 8064 4495 8120
rect 0 8062 4495 8064
rect 0 8032 800 8062
rect 4429 8059 4495 8062
rect 8845 7850 8911 7853
rect 4248 7848 8911 7850
rect 4248 7792 8850 7848
rect 8906 7792 8911 7848
rect 4248 7790 8911 7792
rect 0 7714 800 7744
rect 4248 7714 4308 7790
rect 8845 7787 8911 7790
rect 0 7654 4308 7714
rect 0 7624 800 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 7833 7306 7899 7309
rect 4846 7304 7899 7306
rect 4846 7248 7838 7304
rect 7894 7248 7899 7304
rect 4846 7246 7899 7248
rect 0 7170 800 7200
rect 4846 7170 4906 7246
rect 7833 7243 7899 7246
rect 0 7110 4906 7170
rect 6821 7170 6887 7173
rect 7741 7170 7807 7173
rect 6821 7168 7807 7170
rect 6821 7112 6826 7168
rect 6882 7112 7746 7168
rect 7802 7112 7807 7168
rect 6821 7110 7807 7112
rect 0 7080 800 7110
rect 6821 7107 6887 7110
rect 7741 7107 7807 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 0 6762 800 6792
rect 8569 6762 8635 6765
rect 0 6760 8635 6762
rect 0 6704 8574 6760
rect 8630 6704 8635 6760
rect 0 6702 8635 6704
rect 0 6672 800 6702
rect 8569 6699 8635 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 0 6218 800 6248
rect 3969 6218 4035 6221
rect 0 6216 4035 6218
rect 0 6160 3974 6216
rect 4030 6160 4035 6216
rect 0 6158 4035 6160
rect 0 6128 800 6158
rect 3969 6155 4035 6158
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 0 5810 800 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 800 5750
rect 4061 5747 4127 5750
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 0 5266 800 5296
rect 4061 5266 4127 5269
rect 0 5264 4127 5266
rect 0 5208 4066 5264
rect 4122 5208 4127 5264
rect 0 5206 4127 5208
rect 0 5176 800 5206
rect 4061 5203 4127 5206
rect 7874 4928 8194 4929
rect 0 4858 800 4888
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 4061 4858 4127 4861
rect 0 4856 4127 4858
rect 0 4800 4066 4856
rect 4122 4800 4127 4856
rect 0 4798 4127 4800
rect 0 4768 800 4798
rect 4061 4795 4127 4798
rect 0 4450 800 4480
rect 3969 4450 4035 4453
rect 0 4448 4035 4450
rect 0 4392 3974 4448
rect 4030 4392 4035 4448
rect 0 4390 4035 4392
rect 0 4360 800 4390
rect 3969 4387 4035 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 0 3906 800 3936
rect 3049 3906 3115 3909
rect 0 3904 3115 3906
rect 0 3848 3054 3904
rect 3110 3848 3115 3904
rect 0 3846 3115 3848
rect 0 3816 800 3846
rect 3049 3843 3115 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 3775 15125 3776
rect 0 3498 800 3528
rect 3785 3498 3851 3501
rect 0 3496 3851 3498
rect 0 3440 3790 3496
rect 3846 3440 3851 3496
rect 0 3438 3851 3440
rect 0 3408 800 3438
rect 3785 3435 3851 3438
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 0 2954 800 2984
rect 2773 2954 2839 2957
rect 0 2952 2839 2954
rect 0 2896 2778 2952
rect 2834 2896 2839 2952
rect 0 2894 2839 2896
rect 0 2864 800 2894
rect 2773 2891 2839 2894
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 0 2546 800 2576
rect 3693 2546 3759 2549
rect 0 2544 3759 2546
rect 0 2488 3698 2544
rect 3754 2488 3759 2544
rect 0 2486 3759 2488
rect 0 2456 800 2486
rect 3693 2483 3759 2486
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 0 2002 800 2032
rect 3509 2002 3575 2005
rect 0 2000 3575 2002
rect 0 1944 3514 2000
rect 3570 1944 3575 2000
rect 0 1942 3575 1944
rect 0 1912 800 1942
rect 3509 1939 3575 1942
rect 0 1594 800 1624
rect 3877 1594 3943 1597
rect 0 1592 3943 1594
rect 0 1536 3882 1592
rect 3938 1536 3943 1592
rect 0 1534 3943 1536
rect 0 1504 800 1534
rect 3877 1531 3943 1534
rect 0 1050 800 1080
rect 6453 1050 6519 1053
rect 0 1048 6519 1050
rect 0 992 6458 1048
rect 6514 992 6519 1048
rect 0 990 6519 992
rect 0 960 800 990
rect 6453 987 6519 990
rect 0 642 800 672
rect 3325 642 3391 645
rect 0 640 3391 642
rect 0 584 3330 640
rect 3386 584 3391 640
rect 0 582 3391 584
rect 0 552 800 582
rect 3325 579 3391 582
rect 0 234 800 264
rect 4245 234 4311 237
rect 0 232 4311 234
rect 0 176 4250 232
rect 4306 176 4311 232
rect 0 174 4311 176
rect 0 144 800 174
rect 4245 171 4311 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__decap_12  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608910539
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1608910539
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608910539
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608910539
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1608910539
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1608910539
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1608910539
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1608910539
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608910539
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1608910539
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1608910539
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1608910539
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1608910539
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1608910539
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1608910539
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1608910539
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1608910539
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1608910539
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1608910539
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1608910539
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1608910539
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1608910539
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1608910539
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1608910539
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1608910539
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_220
timestamp 1608910539
transform 1 0 21344 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1608910539
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1608910539
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608910539
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608910539
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1608910539
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608910539
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1608910539
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1608910539
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1608910539
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1608910539
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1608910539
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1608910539
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1608910539
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1608910539
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1608910539
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1608910539
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1608910539
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608910539
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1608910539
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608910539
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608910539
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1608910539
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1608910539
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1608910539
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1608910539
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1608910539
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1608910539
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1608910539
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1608910539
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1608910539
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1608910539
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1608910539
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1608910539
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp 1608910539
transform 1 0 21344 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608910539
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608910539
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1608910539
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1608910539
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1608910539
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1608910539
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1608910539
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1608910539
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1608910539
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1608910539
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1608910539
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1608910539
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1608910539
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1608910539
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1608910539
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608910539
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1608910539
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608910539
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608910539
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1608910539
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1608910539
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1608910539
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1608910539
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1608910539
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1608910539
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1608910539
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1608910539
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1608910539
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1608910539
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_208
timestamp 1608910539
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1608910539
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1608910539
transform 1 0 21528 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1608910539
transform 1 0 21160 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_212
timestamp 1608910539
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _107_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 20792 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608910539
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608910539
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1608910539
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1608910539
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608910539
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608910539
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1608910539
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1608910539
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1608910539
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1608910539
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1608910539
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1608910539
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1608910539
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1608910539
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1608910539
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1608910539
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1608910539
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1608910539
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1608910539
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1608910539
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1608910539
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1608910539
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1608910539
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1608910539
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1608910539
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1608910539
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_204
timestamp 1608910539
transform 1 0 19872 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_196
timestamp 1608910539
transform 1 0 19136 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_202
timestamp 1608910539
transform 1 0 19688 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1608910539
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608910539
transform 1 0 19964 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_213
timestamp 1608910539
transform 1 0 20700 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_209
timestamp 1608910539
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1608910539
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1608910539
transform 1 0 20516 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1608910539
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608910539
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1608910539
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1608910539
transform 1 0 21252 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608910539
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608910539
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_60
timestamp 1608910539
transform 1 0 6624 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_56
timestamp 1608910539
transform 1 0 6256 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1608910539
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1608910539
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_75
timestamp 1608910539
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_63
timestamp 1608910539
transform 1 0 6900 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7176 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _039_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 8188 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1608910539
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1608910539
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1608910539
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1608910539
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1608910539
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1608910539
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1608910539
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_198
timestamp 1608910539
transform 1 0 19320 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_190
timestamp 1608910539
transform 1 0 18584 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1608910539
transform 1 0 20148 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608910539
transform 1 0 19596 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1608910539
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1608910539
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1608910539
transform 1 0 20332 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1608910539
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_31
timestamp 1608910539
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27
timestamp 1608910539
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4140 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_62
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608910539
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_55
timestamp 1608910539
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1608910539
transform 1 0 5428 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_42
timestamp 1608910539
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1608910539
transform 1 0 5152 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_74
timestamp 1608910539
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1608910539
transform 1 0 7084 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8096 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1608910539
transform 1 0 9660 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_89
timestamp 1608910539
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_85
timestamp 1608910539
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1608910539
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_117
timestamp 1608910539
transform 1 0 11868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_105
timestamp 1608910539
transform 1 0 10764 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1608910539
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1608910539
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1608910539
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_184
timestamp 1608910539
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1608910539
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1608910539
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1608910539
transform 1 0 19964 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_201
timestamp 1608910539
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_195
timestamp 1608910539
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_189
timestamp 1608910539
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1608910539
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608910539
transform 1 0 19228 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608910539
transform 1 0 18676 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1608910539
transform 1 0 21068 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_19
timestamp 1608910539
transform 1 0 2852 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp 1608910539
transform 1 0 2484 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1932 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1608910539
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_48
timestamp 1608910539
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5704 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_66
timestamp 1608910539
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 7360 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_102
timestamp 1608910539
transform 1 0 10488 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1608910539
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_114
timestamp 1608910539
transform 1 0 11592 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_138
timestamp 1608910539
transform 1 0 13800 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_126
timestamp 1608910539
transform 1 0 12696 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1608910539
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1608910539
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1608910539
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1608910539
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1608910539
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1608910539
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_16
timestamp 1608910539
transform 1 0 2576 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1608910539
transform 1 0 1932 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_38
timestamp 1608910539
transform 1 0 4600 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4876 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3128 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_58
timestamp 1608910539
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1608910539
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_50
timestamp 1608910539
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1608910539
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8464 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1608910539
transform 1 0 9660 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_89
timestamp 1608910539
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1608910539
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1608910539
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_105
timestamp 1608910539
transform 1 0 10764 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1608910539
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1608910539
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1608910539
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1608910539
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1608910539
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1608910539
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1608910539
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_220
timestamp 1608910539
transform 1 0 21344 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1608910539
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2300 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608910539
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_36
timestamp 1608910539
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1608910539
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 4600 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_62
timestamp 1608910539
transform 1 0 6808 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_59
timestamp 1608910539
transform 1 0 6532 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_51
timestamp 1608910539
transform 1 0 5796 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_47
timestamp 1608910539
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_83
timestamp 1608910539
transform 1 0 8740 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 1608910539
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1608910539
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7544 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1608910539
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1608910539
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1608910539
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1608910539
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1608910539
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1608910539
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1608910539
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1608910539
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1608910539
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1608910539
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608910539
transform 1 0 1748 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_17
timestamp 1608910539
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_11
timestamp 1608910539
transform 1 0 2116 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1608910539
transform 1 0 2852 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_14_28
timestamp 1608910539
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1608910539
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_28
timestamp 1608910539
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1608910539
transform 1 0 3404 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_32
timestamp 1608910539
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4232 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1608910539
transform 1 0 4876 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_62
timestamp 1608910539
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_45
timestamp 1608910539
transform 1 0 5244 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608910539
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1608910539
transform 1 0 6164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_43
timestamp 1608910539
transform 1 0 5060 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5336 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1608910539
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_77
timestamp 1608910539
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_66
timestamp 1608910539
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_71
timestamp 1608910539
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7360 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8372 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8004 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_102
timestamp 1608910539
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1608910539
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_103
timestamp 1608910539
transform 1 0 10580 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_95
timestamp 1608910539
transform 1 0 9844 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_91
timestamp 1608910539
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_106
timestamp 1608910539
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10856 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_119
timestamp 1608910539
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_115
timestamp 1608910539
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1608910539
transform 1 0 12420 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1608910539
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_135
timestamp 1608910539
transform 1 0 13524 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1608910539
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1608910539
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_147
timestamp 1608910539
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_151
timestamp 1608910539
transform 1 0 14996 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_147
timestamp 1608910539
transform 1 0 14628 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15456 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_165
timestamp 1608910539
transform 1 0 16284 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_166
timestamp 1608910539
transform 1 0 16376 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_154
timestamp 1608910539
transform 1 0 15272 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1608910539
transform 1 0 17388 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1608910539
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1608910539
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1608910539
transform 1 0 17480 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16560 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1608910539
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_189
timestamp 1608910539
transform 1 0 18492 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1608910539
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1608910539
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1608910539
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1608910539
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_220
timestamp 1608910539
transform 1 0 21344 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_16
timestamp 1608910539
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 1748 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 2760 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_38
timestamp 1608910539
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_34
timestamp 1608910539
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608910539
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_46
timestamp 1608910539
transform 1 0 5336 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_42
timestamp 1608910539
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1608910539
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8464 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_96
timestamp 1608910539
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10120 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1608910539
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_114
timestamp 1608910539
transform 1 0 11592 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608910539
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_139
timestamp 1608910539
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14076 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_157
timestamp 1608910539
transform 1 0 15548 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16284 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_187
timestamp 1608910539
transform 1 0 18308 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608910539
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608910539
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_199
timestamp 1608910539
transform 1 0 19412 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_211
timestamp 1608910539
transform 1 0 20516 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 1608910539
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 1932 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2944 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1608910539
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1608910539
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_58
timestamp 1608910539
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_53
timestamp 1608910539
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_49
timestamp 1608910539
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_45
timestamp 1608910539
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_left_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6164 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1608910539
transform 1 0 6624 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_80
timestamp 1608910539
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_69
timestamp 1608910539
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7636 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608910539
transform 1 0 8648 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_103
timestamp 1608910539
transform 1 0 10580 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_99
timestamp 1608910539
transform 1 0 10212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_93
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608910539
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1608910539
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608910539
transform 1 0 10304 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_123
timestamp 1608910539
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12604 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10948 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1608910539
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_134
timestamp 1608910539
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1608910539
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15640 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608910539
transform 1 0 14628 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_174
timestamp 1608910539
transform 1 0 17112 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 17480 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1608910539
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_194
timestamp 1608910539
transform 1 0 18952 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1608910539
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_13
timestamp 1608910539
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2484 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1748 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1608910539
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_29
timestamp 1608910539
transform 1 0 3772 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_21
timestamp 1608910539
transform 1 0 3036 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1608910539
transform 1 0 3864 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1608910539
transform 1 0 4876 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608910539
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_55
timestamp 1608910539
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_50
timestamp 1608910539
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1608910539
transform 1 0 5888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1608910539
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7084 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_89
timestamp 1608910539
transform 1 0 9292 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_85
timestamp 1608910539
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_123
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1608910539
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_109
timestamp 1608910539
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11316 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608910539
transform 1 0 12512 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_140
timestamp 1608910539
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_136
timestamp 1608910539
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1608910539
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_127
timestamp 1608910539
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 12972 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 14168 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_166
timestamp 1608910539
transform 1 0 16376 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_162
timestamp 1608910539
transform 1 0 16008 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_158
timestamp 1608910539
transform 1 0 15640 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 16100 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1608910539
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_178
timestamp 1608910539
transform 1 0 17480 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608910539
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1608910539
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1608910539
transform 1 0 19964 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1608910539
transform 1 0 18860 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1608910539
transform 1 0 21068 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_17
timestamp 1608910539
transform 1 0 2668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2852 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2116 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_25
timestamp 1608910539
transform 1 0 3404 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_57
timestamp 1608910539
transform 1 0 6348 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1608910539
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1608910539
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 6072 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6532 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_72
timestamp 1608910539
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1608910539
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7912 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_95
timestamp 1608910539
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1608910539
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10028 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_118
timestamp 1608910539
transform 1 0 11960 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_106
timestamp 1608910539
transform 1 0 10856 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11132 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12144 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_140
timestamp 1608910539
transform 1 0 13984 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1608910539
transform 1 0 13616 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14076 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1608910539
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_174
timestamp 1608910539
transform 1 0 17112 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_170
timestamp 1608910539
transform 1 0 16744 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 17204 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_200
timestamp 1608910539
transform 1 0 19504 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_196
timestamp 1608910539
transform 1 0 19136 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_191
timestamp 1608910539
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608910539
transform 1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1608910539
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1608910539
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608910539
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1608910539
transform 1 0 1932 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1608910539
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608910539
transform 1 0 2300 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608910539
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_16
timestamp 1608910539
transform 1 0 2576 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1608910539
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608910539
transform 1 0 2852 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608910539
transform 1 0 2944 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1608910539
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_23
timestamp 1608910539
transform 1 0 3220 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_29
timestamp 1608910539
transform 1 0 3772 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1608910539
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608910539
transform 1 0 3404 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1608910539
transform 1 0 3496 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_35
timestamp 1608910539
transform 1 0 4324 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4416 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_20_59
timestamp 1608910539
transform 1 0 6532 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_48
timestamp 1608910539
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608910539
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_56
timestamp 1608910539
transform 1 0 6256 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_52
timestamp 1608910539
transform 1 0 5888 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5704 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_20_77
timestamp 1608910539
transform 1 0 8188 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_73
timestamp 1608910539
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_63
timestamp 1608910539
transform 1 0 6900 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1608910539
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8464 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6992 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8556 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1608910539
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_89
timestamp 1608910539
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1608910539
transform 1 0 9476 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1608910539
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_102
timestamp 1608910539
transform 1 0 10488 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1608910539
transform 1 0 10120 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_94
timestamp 1608910539
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_111
timestamp 1608910539
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_106
timestamp 1608910539
transform 1 0 10856 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_109
timestamp 1608910539
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_105
timestamp 1608910539
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1608910539
transform 1 0 11316 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_123
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1608910539
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12512 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11500 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_129
timestamp 1608910539
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_133
timestamp 1608910539
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13156 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_144
timestamp 1608910539
transform 1 0 14352 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_140
timestamp 1608910539
transform 1 0 13984 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_141
timestamp 1608910539
transform 1 0 14076 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_137
timestamp 1608910539
transform 1 0 13708 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 14168 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_145
timestamp 1608910539
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1608910539
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_147
timestamp 1608910539
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_149
timestamp 1608910539
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1608910539
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608910539
transform 1 0 16284 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 14996 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_20_176
timestamp 1608910539
transform 1 0 17296 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_168
timestamp 1608910539
transform 1 0 16560 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_167
timestamp 1608910539
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 17388 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16652 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp 1608910539
transform 1 0 17572 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1608910539
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1608910539
transform 1 0 17480 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608910539
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 17756 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1608910539
transform 1 0 19228 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_204
timestamp 1608910539
transform 1 0 19872 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1608910539
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1608910539
transform 1 0 19044 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1608910539
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1608910539
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1608910539
transform 1 0 20332 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_222
timestamp 1608910539
transform 1 0 21528 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_216
timestamp 1608910539
transform 1 0 20976 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608910539
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_16
timestamp 1608910539
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_8
timestamp 1608910539
transform 1 0 1840 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2760 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608910539
transform 1 0 1472 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_35
timestamp 1608910539
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_24
timestamp 1608910539
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1608910539
transform 1 0 3496 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4508 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1608910539
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_53
timestamp 1608910539
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_82
timestamp 1608910539
transform 1 0 8648 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_78
timestamp 1608910539
transform 1 0 8280 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8740 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_99
timestamp 1608910539
transform 1 0 10212 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1608910539
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11316 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_21_139
timestamp 1608910539
transform 1 0 13892 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 14168 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1608910539
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_151
timestamp 1608910539
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16192 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15180 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_21_177
timestamp 1608910539
transform 1 0 17388 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_173
timestamp 1608910539
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608910539
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1608910539
transform 1 0 19964 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1608910539
transform 1 0 18860 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1608910539
transform 1 0 21068 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_18
timestamp 1608910539
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1608910539
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1608910539
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1608910539
transform 1 0 1932 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1608910539
transform 1 0 2944 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1608910539
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_22_59
timestamp 1608910539
transform 1 0 6532 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_48
timestamp 1608910539
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5704 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_83
timestamp 1608910539
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_78
timestamp 1608910539
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1608910539
transform 1 0 8464 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_104
timestamp 1608910539
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_101
timestamp 1608910539
transform 1 0 10396 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_95
timestamp 1608910539
transform 1 0 9844 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1608910539
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 8924 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608910539
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_left_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 10856 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_22_144
timestamp 1608910539
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_126
timestamp 1608910539
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12880 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1608910539
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_148
timestamp 1608910539
transform 1 0 14720 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 14536 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608910539
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15272 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_22_179
timestamp 1608910539
transform 1 0 17572 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1608910539
transform 1 0 17204 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_170
timestamp 1608910539
transform 1 0 16744 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 17664 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608910539
transform 1 0 16928 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1608910539
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_196
timestamp 1608910539
transform 1 0 19136 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608910539
transform 1 0 19320 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1608910539
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1608910539
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_213
timestamp 1608910539
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608910539
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_16
timestamp 1608910539
transform 1 0 2576 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_8
timestamp 1608910539
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1608910539
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2852 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608910539
transform 1 0 1472 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1608910539
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_35
timestamp 1608910539
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1608910539
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1608910539
transform 1 0 6348 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1608910539
transform 1 0 5796 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608910539
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_74
timestamp 1608910539
transform 1 0 7912 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_68
timestamp 1608910539
transform 1 0 7360 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8004 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_91
timestamp 1608910539
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9660 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_23_125
timestamp 1608910539
transform 1 0 12604 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1608910539
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_117
timestamp 1608910539
transform 1 0 11868 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1608910539
transform 1 0 11500 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_109
timestamp 1608910539
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608910539
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_137
timestamp 1608910539
transform 1 0 13708 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12880 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13984 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_157
timestamp 1608910539
transform 1 0 15548 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_153
timestamp 1608910539
transform 1 0 15180 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_149
timestamp 1608910539
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15916 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1608910539
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_177
timestamp 1608910539
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608910539
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_197
timestamp 1608910539
transform 1 0 19228 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_193
timestamp 1608910539
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 19964 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1608910539
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_16
timestamp 1608910539
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_8
timestamp 1608910539
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608910539
transform 1 0 2760 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608910539
transform 1 0 1472 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_38
timestamp 1608910539
transform 1 0 4600 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_32
timestamp 1608910539
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1608910539
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_26
timestamp 1608910539
transform 1 0 3496 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_22
timestamp 1608910539
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608910539
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4692 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_55
timestamp 1608910539
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6348 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_79
timestamp 1608910539
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_75
timestamp 1608910539
transform 1 0 8004 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_71
timestamp 1608910539
transform 1 0 7636 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_66
timestamp 1608910539
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 7360 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8556 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1608910539
transform 1 0 8096 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_102
timestamp 1608910539
transform 1 0 10488 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1608910539
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608910539
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_122
timestamp 1608910539
transform 1 0 12328 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10856 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608910539
transform 1 0 12512 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1608910539
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1608910539
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_127
timestamp 1608910539
transform 1 0 12788 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 13064 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13984 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608910539
transform 1 0 13524 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_163
timestamp 1608910539
transform 1 0 16100 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1608910539
transform 1 0 15732 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1608910539
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1608910539
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 15456 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608910539
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16192 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_185
timestamp 1608910539
transform 1 0 18124 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_181
timestamp 1608910539
transform 1 0 17756 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_177
timestamp 1608910539
transform 1 0 17388 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_173
timestamp 1608910539
transform 1 0 17020 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 17940 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 17572 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17204 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_205
timestamp 1608910539
transform 1 0 19964 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18492 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1608910539
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1608910539
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608910539
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_16
timestamp 1608910539
transform 1 0 2576 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_8
timestamp 1608910539
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1608910539
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608910539
transform 1 0 1472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_40
timestamp 1608910539
transform 1 0 4784 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_28
timestamp 1608910539
transform 1 0 3680 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4876 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1608910539
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_55
timestamp 1608910539
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_50
timestamp 1608910539
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608910539
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1608910539
transform 1 0 5888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_81
timestamp 1608910539
transform 1 0 8556 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_77
timestamp 1608910539
transform 1 0 8188 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_65
timestamp 1608910539
transform 1 0 7084 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7360 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8648 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_98
timestamp 1608910539
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10304 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1608910539
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_109
timestamp 1608910539
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608910539
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 11316 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_132
timestamp 1608910539
transform 1 0 13248 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13616 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 1608910539
transform 1 0 16100 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_152
timestamp 1608910539
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 15272 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1608910539
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_176
timestamp 1608910539
transform 1 0 17296 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_171
timestamp 1608910539
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1608910539
transform 1 0 16468 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 16560 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608910539
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1608910539
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608910539
transform 1 0 17020 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1608910539
transform 1 0 19964 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1608910539
transform 1 0 18860 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1608910539
transform 1 0 21068 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_8
timestamp 1608910539
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1608910539
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1608910539
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608910539
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608910539
transform 1 0 1472 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1608910539
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_19
timestamp 1608910539
transform 1 0 2852 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_11
timestamp 1608910539
transform 1 0 2116 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2760 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2944 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_24
timestamp 1608910539
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_35
timestamp 1608910539
transform 1 0 4324 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1608910539
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608910539
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3496 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4876 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608910539
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_62
timestamp 1608910539
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_49
timestamp 1608910539
transform 1 0 5612 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_46
timestamp 1608910539
transform 1 0 5336 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_42
timestamp 1608910539
transform 1 0 4968 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_57
timestamp 1608910539
transform 1 0 6348 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608910539
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_81
timestamp 1608910539
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_79
timestamp 1608910539
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8556 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6900 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7084 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1608910539
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1608910539
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608910539
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9108 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_101
timestamp 1608910539
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_96
timestamp 1608910539
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1608910539
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_95
timestamp 1608910539
transform 1 0 9844 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1608910539
transform 1 0 10120 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_109
timestamp 1608910539
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_105
timestamp 1608910539
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1608910539
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11316 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1608910539
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_123
timestamp 1608910539
transform 1 0 12420 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608910539
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10948 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 1608910539
transform 1 0 14076 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_137
timestamp 1608910539
transform 1 0 13708 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1608910539
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_137
timestamp 1608910539
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_127
timestamp 1608910539
transform 1 0 12788 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 13432 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 12880 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13892 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 14168 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_158
timestamp 1608910539
transform 1 0 15640 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_160
timestamp 1608910539
transform 1 0 15824 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_156
timestamp 1608910539
transform 1 0 15456 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1608910539
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1608910539
transform 1 0 14720 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 15640 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608910539
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16376 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_27_184
timestamp 1608910539
transform 1 0 18032 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1608910539
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_170
timestamp 1608910539
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_182
timestamp 1608910539
transform 1 0 17848 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608910539
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16928 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 18124 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 18032 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_201
timestamp 1608910539
transform 1 0 19596 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_200
timestamp 1608910539
transform 1 0 19504 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1608910539
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_213
timestamp 1608910539
transform 1 0 20700 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1608910539
transform 1 0 20884 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1608910539
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608910539
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_17
timestamp 1608910539
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_9
timestamp 1608910539
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1608910539
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608910539
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2116 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608910539
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608910539
transform 1 0 1564 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1608910539
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1608910539
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1608910539
transform 1 0 3220 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608910539
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_62
timestamp 1608910539
transform 1 0 6808 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_58
timestamp 1608910539
transform 1 0 6440 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_45
timestamp 1608910539
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6624 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5612 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_79
timestamp 1608910539
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_75
timestamp 1608910539
transform 1 0 8004 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_69
timestamp 1608910539
transform 1 0 7452 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_left_track_1.prog_clk
timestamp 1608910539
transform 1 0 8096 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8556 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1608910539
transform 1 0 7176 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1608910539
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608910539
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_124
timestamp 1608910539
transform 1 0 12512 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_120
timestamp 1608910539
transform 1 0 12144 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1608910539
transform 1 0 11132 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12328 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11316 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_28_142
timestamp 1608910539
transform 1 0 14168 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1608910539
transform 1 0 13800 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_134
timestamp 1608910539
transform 1 0 13432 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_128
timestamp 1608910539
transform 1 0 12880 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608910539
transform 1 0 13524 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1608910539
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_147
timestamp 1608910539
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608910539
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15272 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_28_182
timestamp 1608910539
transform 1 0 17848 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_174
timestamp 1608910539
transform 1 0 17112 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_170
timestamp 1608910539
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 16928 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1608910539
transform 1 0 18124 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_199
timestamp 1608910539
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1608910539
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608910539
transform 1 0 19136 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_215
timestamp 1608910539
transform 1 0 20884 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1608910539
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608910539
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608910539
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_17
timestamp 1608910539
transform 1 0 2668 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1608910539
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1608910539
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608910539
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2944 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608910539
transform 1 0 2300 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608910539
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_41
timestamp 1608910539
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp 1608910539
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1608910539
transform 1 0 4600 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1608910539
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1608910539
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608910539
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5060 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_76
timestamp 1608910539
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_70
timestamp 1608910539
transform 1 0 7544 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 6992 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 8280 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1608910539
transform 1 0 7820 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_96
timestamp 1608910539
transform 1 0 9936 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_84
timestamp 1608910539
transform 1 0 8832 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_123
timestamp 1608910539
transform 1 0 12420 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1608910539
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_108
timestamp 1608910539
transform 1 0 11040 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 12512 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608910539
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_144
timestamp 1608910539
transform 1 0 14352 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_126
timestamp 1608910539
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 12880 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_158
timestamp 1608910539
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_148
timestamp 1608910539
transform 1 0 14720 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14812 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15824 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_29_180
timestamp 1608910539
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_176
timestamp 1608910539
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 17480 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608910539
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_202
timestamp 1608910539
transform 1 0 19688 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_190
timestamp 1608910539
transform 1 0 18584 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_222
timestamp 1608910539
transform 1 0 21528 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_214
timestamp 1608910539
transform 1 0 20792 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608910539
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_15
timestamp 1608910539
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1608910539
transform 1 0 1380 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608910539
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2852 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1932 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_41
timestamp 1608910539
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_28
timestamp 1608910539
transform 1 0 3680 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608910539
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_52
timestamp 1608910539
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6072 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5060 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_30_78
timestamp 1608910539
transform 1 0 8280 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_67
timestamp 1608910539
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_63
timestamp 1608910539
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7452 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8556 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1608910539
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608910539
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9660 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_109
timestamp 1608910539
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11316 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_140
timestamp 1608910539
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_127
timestamp 1608910539
transform 1 0 12788 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13156 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_163
timestamp 1608910539
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1608910539
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608910539
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1608910539
transform 1 0 16284 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_184
timestamp 1608910539
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_174
timestamp 1608910539
transform 1 0 17112 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 17480 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608910539
transform 1 0 18216 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_208
timestamp 1608910539
transform 1 0 20240 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_196
timestamp 1608910539
transform 1 0 19136 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1608910539
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608910539
transform 1 0 18768 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1608910539
transform 1 0 21436 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1608910539
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 21252 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608910539
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608910539
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_15
timestamp 1608910539
transform 1 0 2484 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1608910539
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608910539
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1932 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608910539
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_41
timestamp 1608910539
transform 1 0 4876 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_37
timestamp 1608910539
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4692 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 3036 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1608910539
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608910539
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5060 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_64
timestamp 1608910539
transform 1 0 6992 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7360 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_92
timestamp 1608910539
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_88
timestamp 1608910539
transform 1 0 9200 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_84
timestamp 1608910539
transform 1 0 8832 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9752 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1608910539
transform 1 0 9292 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_123
timestamp 1608910539
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1608910539
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_110
timestamp 1608910539
transform 1 0 11224 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608910539
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 11500 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12512 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_145
timestamp 1608910539
transform 1 0 14444 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1608910539
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_130
timestamp 1608910539
transform 1 0 13064 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13340 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608910539
transform 1 0 14076 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_163
timestamp 1608910539
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_154
timestamp 1608910539
transform 1 0 15272 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16284 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 15548 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14720 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1608910539
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1608910539
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608910539
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 17020 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_208
timestamp 1608910539
transform 1 0 20240 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1608910539
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_190
timestamp 1608910539
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608910539
transform 1 0 18768 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1608910539
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608910539
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 20332 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1608910539
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1608910539
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608910539
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1564 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 2300 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_32_34
timestamp 1608910539
transform 1 0 4232 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1608910539
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608910539
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4508 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_32_46
timestamp 1608910539
transform 1 0 5336 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5612 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_79
timestamp 1608910539
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1608910539
transform 1 0 7084 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8188 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8556 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_32_95
timestamp 1608910539
transform 1 0 9844 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1608910539
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608910539
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10120 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_124
timestamp 1608910539
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1608910539
transform 1 0 11592 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1608910539
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1608910539
transform 1 0 13800 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_130
timestamp 1608910539
transform 1 0 13064 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13248 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608910539
transform 1 0 12696 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608910539
transform 1 0 13984 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_164
timestamp 1608910539
transform 1 0 16192 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_158
timestamp 1608910539
transform 1 0 15640 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_150
timestamp 1608910539
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608910539
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608910539
transform 1 0 16376 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608910539
transform 1 0 15824 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608910539
transform 1 0 15272 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608910539
transform 1 0 14536 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_186
timestamp 1608910539
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_176
timestamp 1608910539
transform 1 0 17296 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_170
timestamp 1608910539
transform 1 0 16744 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608910539
transform 1 0 16928 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_198
timestamp 1608910539
transform 1 0 19320 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_192
timestamp 1608910539
transform 1 0 18768 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608910539
transform 1 0 18952 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608910539
transform 1 0 18400 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1608910539
transform 1 0 20884 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_210
timestamp 1608910539
transform 1 0 20424 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608910539
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608910539
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_17
timestamp 1608910539
transform 1 0 2668 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1608910539
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1608910539
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608910539
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608910539
transform 1 0 2300 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608910539
transform 1 0 1748 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_40
timestamp 1608910539
transform 1 0 4784 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_32
timestamp 1608910539
transform 1 0 4048 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_25
timestamp 1608910539
transform 1 0 3404 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_21
timestamp 1608910539
transform 1 0 3036 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608910539
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608910539
transform 1 0 3128 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608910539
transform 1 0 4876 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_56
timestamp 1608910539
transform 1 0 6256 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1608910539
transform 1 0 5152 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608910539
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_74
timestamp 1608910539
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_71
timestamp 1608910539
transform 1 0 7636 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_63
timestamp 1608910539
transform 1 0 6900 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7728 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8096 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1608910539
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_89
timestamp 1608910539
transform 1 0 9292 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_85
timestamp 1608910539
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608910539
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_125
timestamp 1608910539
transform 1 0 12604 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_118
timestamp 1608910539
transform 1 0 11960 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_106
timestamp 1608910539
transform 1 0 10856 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608910539
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_145
timestamp 1608910539
transform 1 0 14444 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_133
timestamp 1608910539
transform 1 0 13340 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12788 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608910539
transform 1 0 14076 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1608910539
transform 1 0 15456 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_153
timestamp 1608910539
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608910539
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_187
timestamp 1608910539
transform 1 0 18308 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_180
timestamp 1608910539
transform 1 0 17664 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1608910539
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608910539
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_199
timestamp 1608910539
transform 1 0 19412 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1608910539
transform 1 0 21528 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1608910539
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_211
timestamp 1608910539
transform 1 0 20516 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608910539
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608910539
transform -1 0 21896 0 1 20128
box -38 -48 314 592
<< labels >>
rlabel metal3 s 22200 11432 23000 11552 6 ccff_head
port 0 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 ccff_tail
port 1 nsew signal tristate
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[0]
port 2 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[10]
port 3 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[11]
port 4 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[12]
port 5 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[13]
port 6 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[14]
port 7 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[15]
port 8 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[16]
port 9 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 10 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[18]
port 11 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_in[19]
port 12 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[1]
port 13 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[2]
port 14 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[3]
port 15 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[4]
port 16 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[5]
port 17 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[6]
port 18 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[7]
port 19 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[8]
port 20 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[9]
port 21 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[0]
port 22 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[10]
port 23 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[11]
port 24 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[12]
port 25 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[13]
port 26 nsew signal tristate
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[14]
port 27 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[15]
port 28 nsew signal tristate
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[16]
port 29 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[17]
port 30 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[18]
port 31 nsew signal tristate
rlabel metal3 s 0 22584 800 22704 6 chanx_left_out[19]
port 32 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[1]
port 33 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[2]
port 34 nsew signal tristate
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[3]
port 35 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[4]
port 36 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[5]
port 37 nsew signal tristate
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[6]
port 38 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[7]
port 39 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[8]
port 40 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[9]
port 41 nsew signal tristate
rlabel metal2 s 3882 22200 3938 23000 6 chany_top_in[0]
port 42 nsew signal input
rlabel metal2 s 8482 22200 8538 23000 6 chany_top_in[10]
port 43 nsew signal input
rlabel metal2 s 8942 22200 8998 23000 6 chany_top_in[11]
port 44 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[12]
port 45 nsew signal input
rlabel metal2 s 9862 22200 9918 23000 6 chany_top_in[13]
port 46 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[14]
port 47 nsew signal input
rlabel metal2 s 10782 22200 10838 23000 6 chany_top_in[15]
port 48 nsew signal input
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_in[16]
port 49 nsew signal input
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_in[17]
port 50 nsew signal input
rlabel metal2 s 12162 22200 12218 23000 6 chany_top_in[18]
port 51 nsew signal input
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_in[19]
port 52 nsew signal input
rlabel metal2 s 4342 22200 4398 23000 6 chany_top_in[1]
port 53 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[2]
port 54 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[3]
port 55 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 chany_top_in[4]
port 56 nsew signal input
rlabel metal2 s 6182 22200 6238 23000 6 chany_top_in[5]
port 57 nsew signal input
rlabel metal2 s 6642 22200 6698 23000 6 chany_top_in[6]
port 58 nsew signal input
rlabel metal2 s 7102 22200 7158 23000 6 chany_top_in[7]
port 59 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[8]
port 60 nsew signal input
rlabel metal2 s 8022 22200 8078 23000 6 chany_top_in[9]
port 61 nsew signal input
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_out[0]
port 62 nsew signal tristate
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 63 nsew signal tristate
rlabel metal2 s 18142 22200 18198 23000 6 chany_top_out[11]
port 64 nsew signal tristate
rlabel metal2 s 18602 22200 18658 23000 6 chany_top_out[12]
port 65 nsew signal tristate
rlabel metal2 s 19062 22200 19118 23000 6 chany_top_out[13]
port 66 nsew signal tristate
rlabel metal2 s 19522 22200 19578 23000 6 chany_top_out[14]
port 67 nsew signal tristate
rlabel metal2 s 19982 22200 20038 23000 6 chany_top_out[15]
port 68 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[16]
port 69 nsew signal tristate
rlabel metal2 s 20902 22200 20958 23000 6 chany_top_out[17]
port 70 nsew signal tristate
rlabel metal2 s 21362 22200 21418 23000 6 chany_top_out[18]
port 71 nsew signal tristate
rlabel metal2 s 21822 22200 21878 23000 6 chany_top_out[19]
port 72 nsew signal tristate
rlabel metal2 s 13542 22200 13598 23000 6 chany_top_out[1]
port 73 nsew signal tristate
rlabel metal2 s 14002 22200 14058 23000 6 chany_top_out[2]
port 74 nsew signal tristate
rlabel metal2 s 14462 22200 14518 23000 6 chany_top_out[3]
port 75 nsew signal tristate
rlabel metal2 s 14922 22200 14978 23000 6 chany_top_out[4]
port 76 nsew signal tristate
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[5]
port 77 nsew signal tristate
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[6]
port 78 nsew signal tristate
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[7]
port 79 nsew signal tristate
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[8]
port 80 nsew signal tristate
rlabel metal2 s 17222 22200 17278 23000 6 chany_top_out[9]
port 81 nsew signal tristate
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_11_
port 82 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_13_
port 83 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_15_
port 84 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 left_bottom_grid_pin_17_
port 85 nsew signal input
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_1_
port 86 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_3_
port 87 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_5_
port 88 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_7_
port 89 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_9_
port 90 nsew signal input
rlabel metal2 s 22282 22200 22338 23000 6 prog_clk_0_N_in
port 91 nsew signal input
rlabel metal2 s 202 22200 258 23000 6 top_left_grid_pin_42_
port 92 nsew signal input
rlabel metal2 s 662 22200 718 23000 6 top_left_grid_pin_43_
port 93 nsew signal input
rlabel metal2 s 1122 22200 1178 23000 6 top_left_grid_pin_44_
port 94 nsew signal input
rlabel metal2 s 1582 22200 1638 23000 6 top_left_grid_pin_45_
port 95 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_46_
port 96 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 top_left_grid_pin_47_
port 97 nsew signal input
rlabel metal2 s 2962 22200 3018 23000 6 top_left_grid_pin_48_
port 98 nsew signal input
rlabel metal2 s 3422 22200 3478 23000 6 top_left_grid_pin_49_
port 99 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 top_right_grid_pin_1_
port 100 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 101 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 102 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 103 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 104 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 105 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
