VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__1_
  CLASS BLOCK ;
  FOREIGN sb_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 120.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 2.760 120.000 3.360 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 117.600 4.970 120.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 2.400 2.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 2.400 5.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 2.400 9.480 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 117.600 14.170 120.000 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.400 13.560 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 8.200 120.000 8.800 ;
    END
  END bottom_right_grid_pin_11_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 117.600 23.370 120.000 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 2.400 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 117.600 32.570 120.000 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 13.640 120.000 14.240 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 2.400 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 2.400 29.880 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 2.400 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 2.400 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.400 37.360 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 2.400 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.490 117.600 41.770 120.000 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 2.400 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.400 41.440 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 19.080 120.000 19.680 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 2.400 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 117.600 50.970 120.000 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 2.400 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 2.400 45.520 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.400 49.600 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 24.520 120.000 25.120 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 2.400 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 29.960 120.000 30.560 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 2.400 53.680 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 35.400 120.000 36.000 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 2.400 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 2.400 57.760 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 2.400 61.840 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 117.600 60.170 120.000 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 2.400 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 2.400 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 117.600 69.370 120.000 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 2.400 65.240 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 2.400 69.320 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 40.840 120.000 41.440 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 46.280 120.000 46.880 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 51.720 120.000 52.320 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 57.160 120.000 57.760 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.290 117.600 78.570 120.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 117.600 87.770 120.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 62.600 120.000 63.200 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 2.400 81.560 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 68.040 120.000 68.640 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 117.600 96.970 120.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 2.400 89.720 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 73.480 120.000 74.080 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 2.400 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 78.920 120.000 79.520 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 84.360 120.000 84.960 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.400 93.120 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 2.400 97.200 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 2.400 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 89.800 120.000 90.400 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 95.240 120.000 95.840 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 2.400 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.400 101.280 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 2.400 105.360 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 100.680 120.000 101.280 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 2.400 109.440 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 117.600 106.170 120.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 117.600 106.120 120.000 106.720 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 2.400 113.520 ;
    END
  END left_bottom_grid_pin_12_
  PIN left_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 111.560 120.000 112.160 ;
    END
  END left_top_grid_pin_10_
  PIN right_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 117.600 115.370 120.000 ;
    END
  END right_bottom_grid_pin_12_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 2.400 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 2.400 117.600 ;
    END
  END top_left_grid_pin_13_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 117.600 117.000 120.000 117.600 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 24.720 10.640 26.320 109.040 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 44.720 10.640 46.320 109.040 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 0.145 0.425 114.080 117.895 ;
      LAYER met1 ;
        RECT 0.070 0.040 118.150 117.940 ;
      LAYER met2 ;
        RECT 0.090 117.320 4.410 118.050 ;
        RECT 5.250 117.320 13.610 118.050 ;
        RECT 14.450 117.320 22.810 118.050 ;
        RECT 23.650 117.320 32.010 118.050 ;
        RECT 32.850 117.320 41.210 118.050 ;
        RECT 42.050 117.320 50.410 118.050 ;
        RECT 51.250 117.320 59.610 118.050 ;
        RECT 60.450 117.320 68.810 118.050 ;
        RECT 69.650 117.320 78.010 118.050 ;
        RECT 78.850 117.320 87.210 118.050 ;
        RECT 88.050 117.320 96.410 118.050 ;
        RECT 97.250 117.320 105.610 118.050 ;
        RECT 106.450 117.320 114.810 118.050 ;
        RECT 115.650 117.320 118.130 118.050 ;
        RECT 0.090 2.680 118.130 117.320 ;
        RECT 0.090 0.010 2.110 2.680 ;
        RECT 2.950 0.010 6.710 2.680 ;
        RECT 7.550 0.010 11.770 2.680 ;
        RECT 12.610 0.010 16.830 2.680 ;
        RECT 17.670 0.010 21.890 2.680 ;
        RECT 22.730 0.010 26.950 2.680 ;
        RECT 27.790 0.010 32.010 2.680 ;
        RECT 32.850 0.010 37.070 2.680 ;
        RECT 37.910 0.010 42.130 2.680 ;
        RECT 42.970 0.010 46.730 2.680 ;
        RECT 47.570 0.010 51.790 2.680 ;
        RECT 52.630 0.010 56.850 2.680 ;
        RECT 57.690 0.010 61.910 2.680 ;
        RECT 62.750 0.010 66.970 2.680 ;
        RECT 67.810 0.010 72.030 2.680 ;
        RECT 72.870 0.010 77.090 2.680 ;
        RECT 77.930 0.010 82.150 2.680 ;
        RECT 82.990 0.010 86.750 2.680 ;
        RECT 87.590 0.010 91.810 2.680 ;
        RECT 92.650 0.010 96.870 2.680 ;
        RECT 97.710 0.010 101.930 2.680 ;
        RECT 102.770 0.010 106.990 2.680 ;
        RECT 107.830 0.010 112.050 2.680 ;
        RECT 112.890 0.010 117.110 2.680 ;
        RECT 117.950 0.010 118.130 2.680 ;
      LAYER met3 ;
        RECT 2.800 116.600 117.200 117.000 ;
        RECT 0.065 113.920 118.410 116.600 ;
        RECT 2.800 112.560 118.410 113.920 ;
        RECT 2.800 112.520 117.200 112.560 ;
        RECT 0.065 111.160 117.200 112.520 ;
        RECT 0.065 109.840 118.410 111.160 ;
        RECT 2.800 108.440 118.410 109.840 ;
        RECT 0.065 107.120 118.410 108.440 ;
        RECT 0.065 105.760 117.200 107.120 ;
        RECT 2.800 105.720 117.200 105.760 ;
        RECT 2.800 104.360 118.410 105.720 ;
        RECT 0.065 101.680 118.410 104.360 ;
        RECT 2.800 100.280 117.200 101.680 ;
        RECT 0.065 97.600 118.410 100.280 ;
        RECT 2.800 96.240 118.410 97.600 ;
        RECT 2.800 96.200 117.200 96.240 ;
        RECT 0.065 94.840 117.200 96.200 ;
        RECT 0.065 93.520 118.410 94.840 ;
        RECT 2.800 92.120 118.410 93.520 ;
        RECT 0.065 90.800 118.410 92.120 ;
        RECT 0.065 90.120 117.200 90.800 ;
        RECT 2.800 89.400 117.200 90.120 ;
        RECT 2.800 88.720 118.410 89.400 ;
        RECT 0.065 86.040 118.410 88.720 ;
        RECT 2.800 85.360 118.410 86.040 ;
        RECT 2.800 84.640 117.200 85.360 ;
        RECT 0.065 83.960 117.200 84.640 ;
        RECT 0.065 81.960 118.410 83.960 ;
        RECT 2.800 80.560 118.410 81.960 ;
        RECT 0.065 79.920 118.410 80.560 ;
        RECT 0.065 78.520 117.200 79.920 ;
        RECT 0.065 77.880 118.410 78.520 ;
        RECT 2.800 76.480 118.410 77.880 ;
        RECT 0.065 74.480 118.410 76.480 ;
        RECT 0.065 73.800 117.200 74.480 ;
        RECT 2.800 73.080 117.200 73.800 ;
        RECT 2.800 72.400 118.410 73.080 ;
        RECT 0.065 69.720 118.410 72.400 ;
        RECT 2.800 69.040 118.410 69.720 ;
        RECT 2.800 68.320 117.200 69.040 ;
        RECT 0.065 67.640 117.200 68.320 ;
        RECT 0.065 65.640 118.410 67.640 ;
        RECT 2.800 64.240 118.410 65.640 ;
        RECT 0.065 63.600 118.410 64.240 ;
        RECT 0.065 62.240 117.200 63.600 ;
        RECT 2.800 62.200 117.200 62.240 ;
        RECT 2.800 60.840 118.410 62.200 ;
        RECT 0.065 58.160 118.410 60.840 ;
        RECT 2.800 56.760 117.200 58.160 ;
        RECT 0.065 54.080 118.410 56.760 ;
        RECT 2.800 52.720 118.410 54.080 ;
        RECT 2.800 52.680 117.200 52.720 ;
        RECT 0.065 51.320 117.200 52.680 ;
        RECT 0.065 50.000 118.410 51.320 ;
        RECT 2.800 48.600 118.410 50.000 ;
        RECT 0.065 47.280 118.410 48.600 ;
        RECT 0.065 45.920 117.200 47.280 ;
        RECT 2.800 45.880 117.200 45.920 ;
        RECT 2.800 44.520 118.410 45.880 ;
        RECT 0.065 41.840 118.410 44.520 ;
        RECT 2.800 40.440 117.200 41.840 ;
        RECT 0.065 37.760 118.410 40.440 ;
        RECT 2.800 36.400 118.410 37.760 ;
        RECT 2.800 36.360 117.200 36.400 ;
        RECT 0.065 35.000 117.200 36.360 ;
        RECT 0.065 33.680 118.410 35.000 ;
        RECT 2.800 32.280 118.410 33.680 ;
        RECT 0.065 30.960 118.410 32.280 ;
        RECT 0.065 30.280 117.200 30.960 ;
        RECT 2.800 29.560 117.200 30.280 ;
        RECT 2.800 28.880 118.410 29.560 ;
        RECT 0.065 26.200 118.410 28.880 ;
        RECT 2.800 25.520 118.410 26.200 ;
        RECT 2.800 24.800 117.200 25.520 ;
        RECT 0.065 24.120 117.200 24.800 ;
        RECT 0.065 22.120 118.410 24.120 ;
        RECT 2.800 20.720 118.410 22.120 ;
        RECT 0.065 20.080 118.410 20.720 ;
        RECT 0.065 18.680 117.200 20.080 ;
        RECT 0.065 18.040 118.410 18.680 ;
        RECT 2.800 16.640 118.410 18.040 ;
        RECT 0.065 14.640 118.410 16.640 ;
        RECT 0.065 13.960 117.200 14.640 ;
        RECT 2.800 13.240 117.200 13.960 ;
        RECT 2.800 12.560 118.410 13.240 ;
        RECT 0.065 9.880 118.410 12.560 ;
        RECT 2.800 9.200 118.410 9.880 ;
        RECT 2.800 8.480 117.200 9.200 ;
        RECT 0.065 7.800 117.200 8.480 ;
        RECT 0.065 5.800 118.410 7.800 ;
        RECT 2.800 4.400 118.410 5.800 ;
        RECT 0.065 3.760 118.410 4.400 ;
        RECT 0.065 2.400 117.200 3.760 ;
        RECT 2.800 2.360 117.200 2.400 ;
        RECT 2.800 1.000 118.410 2.360 ;
        RECT 0.065 0.175 118.410 1.000 ;
      LAYER met4 ;
        RECT 0.295 109.440 118.385 115.425 ;
        RECT 0.295 10.240 24.320 109.440 ;
        RECT 26.720 10.240 44.320 109.440 ;
        RECT 46.720 10.240 118.385 109.440 ;
        RECT 0.295 0.175 118.385 10.240 ;
      LAYER met5 ;
        RECT 1.500 4.300 110.740 101.100 ;
  END
END sb_1__1_
END LIBRARY

