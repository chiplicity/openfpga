magic
tech EFS8A
magscale 1 2
timestamp 1603801254
<< locali >>
rect 9965 16983 9999 17085
rect 15669 16031 15703 16201
rect 12633 15351 12667 15657
rect 1961 14875 1995 15113
rect 17693 14807 17727 15045
rect 14841 13855 14875 13957
rect 24317 12767 24351 12937
rect 18061 8415 18095 8517
rect 10057 5559 10091 5729
rect 2881 5083 2915 5185
rect 10241 5015 10275 5185
rect 7665 3927 7699 4233
rect 7113 3383 7147 3485
rect 16037 2839 16071 3145
<< viali >>
rect 17141 24361 17175 24395
rect 18245 24361 18279 24395
rect 10676 24225 10710 24259
rect 11656 24225 11690 24259
rect 16957 24225 16991 24259
rect 18061 24225 18095 24259
rect 10747 24021 10781 24055
rect 11759 24021 11793 24055
rect 1593 23817 1627 23851
rect 10701 23817 10735 23851
rect 14565 23817 14599 23851
rect 16221 23817 16255 23851
rect 18245 23817 18279 23851
rect 20361 23817 20395 23851
rect 21465 23817 21499 23851
rect 22569 23817 22603 23851
rect 24777 23817 24811 23851
rect 1409 23613 1443 23647
rect 8953 23613 8987 23647
rect 9413 23613 9447 23647
rect 11136 23613 11170 23647
rect 12484 23613 12518 23647
rect 12909 23613 12943 23647
rect 14381 23613 14415 23647
rect 14933 23613 14967 23647
rect 16037 23613 16071 23647
rect 16589 23613 16623 23647
rect 17877 23613 17911 23647
rect 18061 23613 18095 23647
rect 20177 23613 20211 23647
rect 21281 23613 21315 23647
rect 21833 23613 21867 23647
rect 22385 23613 22419 23647
rect 22937 23613 22971 23647
rect 24593 23613 24627 23647
rect 25145 23613 25179 23647
rect 2053 23477 2087 23511
rect 9137 23477 9171 23511
rect 9965 23477 9999 23511
rect 11207 23477 11241 23511
rect 11621 23477 11655 23511
rect 12587 23477 12621 23511
rect 17049 23477 17083 23511
rect 18705 23477 18739 23511
rect 20821 23477 20855 23511
rect 1593 23273 1627 23307
rect 11161 23273 11195 23307
rect 13691 23273 13725 23307
rect 18245 23273 18279 23307
rect 24777 23273 24811 23307
rect 9873 23205 9907 23239
rect 1409 23137 1443 23171
rect 7332 23137 7366 23171
rect 8620 23137 8654 23171
rect 11320 23137 11354 23171
rect 12300 23137 12334 23171
rect 13588 23137 13622 23171
rect 15552 23137 15586 23171
rect 16808 23137 16842 23171
rect 18061 23137 18095 23171
rect 24593 23137 24627 23171
rect 7757 23069 7791 23103
rect 9781 23069 9815 23103
rect 10149 23069 10183 23103
rect 7435 22933 7469 22967
rect 8723 22933 8757 22967
rect 11391 22933 11425 22967
rect 12403 22933 12437 22967
rect 15623 22933 15657 22967
rect 16911 22933 16945 22967
rect 1593 22729 1627 22763
rect 6285 22729 6319 22763
rect 8585 22729 8619 22763
rect 10609 22729 10643 22763
rect 14289 22729 14323 22763
rect 15577 22729 15611 22763
rect 16773 22729 16807 22763
rect 7205 22661 7239 22695
rect 14611 22661 14645 22695
rect 17095 22661 17129 22695
rect 18245 22661 18279 22695
rect 7389 22593 7423 22627
rect 7665 22593 7699 22627
rect 9965 22593 9999 22627
rect 12909 22593 12943 22627
rect 1409 22525 1443 22559
rect 5784 22525 5818 22559
rect 6653 22525 6687 22559
rect 10828 22525 10862 22559
rect 11621 22525 11655 22559
rect 12449 22525 12483 22559
rect 13277 22525 13311 22559
rect 13512 22525 13546 22559
rect 14524 22525 14558 22559
rect 14933 22525 14967 22559
rect 17024 22525 17058 22559
rect 17417 22525 17451 22559
rect 5871 22457 5905 22491
rect 7481 22457 7515 22491
rect 9321 22457 9355 22491
rect 9413 22457 9447 22491
rect 13599 22457 13633 22491
rect 14013 22457 14047 22491
rect 2053 22389 2087 22423
rect 9045 22389 9079 22423
rect 10241 22389 10275 22423
rect 10931 22389 10965 22423
rect 11345 22389 11379 22423
rect 12633 22389 12667 22423
rect 15669 22389 15703 22423
rect 24593 22389 24627 22423
rect 8769 22185 8803 22219
rect 11069 22185 11103 22219
rect 12357 22185 12391 22219
rect 5181 22117 5215 22151
rect 7389 22117 7423 22151
rect 10149 22117 10183 22151
rect 13185 22117 13219 22151
rect 13277 22117 13311 22151
rect 16129 22117 16163 22151
rect 6228 22049 6262 22083
rect 11564 22049 11598 22083
rect 1685 21981 1719 22015
rect 6331 21981 6365 22015
rect 7297 21981 7331 22015
rect 7573 21981 7607 22015
rect 10057 21981 10091 22015
rect 13461 21981 13495 22015
rect 14289 21981 14323 22015
rect 16037 21981 16071 22015
rect 10609 21913 10643 21947
rect 16589 21913 16623 21947
rect 9321 21845 9355 21879
rect 11667 21845 11701 21879
rect 12817 21845 12851 21879
rect 1593 21641 1627 21675
rect 5641 21641 5675 21675
rect 8309 21641 8343 21675
rect 11529 21641 11563 21675
rect 13829 21641 13863 21675
rect 24777 21641 24811 21675
rect 10977 21573 11011 21607
rect 15301 21573 15335 21607
rect 16497 21573 16531 21607
rect 7573 21505 7607 21539
rect 8861 21505 8895 21539
rect 9137 21505 9171 21539
rect 10425 21505 10459 21539
rect 12265 21505 12299 21539
rect 12817 21505 12851 21539
rect 13461 21505 13495 21539
rect 14381 21505 14415 21539
rect 15945 21505 15979 21539
rect 17233 21505 17267 21539
rect 1409 21437 1443 21471
rect 2053 21437 2087 21471
rect 4604 21437 4638 21471
rect 5800 21437 5834 21471
rect 18128 21437 18162 21471
rect 24593 21437 24627 21471
rect 6285 21369 6319 21403
rect 7297 21369 7331 21403
rect 7389 21369 7423 21403
rect 8953 21369 8987 21403
rect 10517 21369 10551 21403
rect 12909 21369 12943 21403
rect 14473 21369 14507 21403
rect 15025 21369 15059 21403
rect 16037 21369 16071 21403
rect 16957 21369 16991 21403
rect 4675 21301 4709 21335
rect 5089 21301 5123 21335
rect 5871 21301 5905 21335
rect 6653 21301 6687 21335
rect 7113 21301 7147 21335
rect 8677 21301 8711 21335
rect 9873 21301 9907 21335
rect 10149 21301 10183 21335
rect 14197 21301 14231 21335
rect 15761 21301 15795 21335
rect 18199 21301 18233 21335
rect 18613 21301 18647 21335
rect 25145 21301 25179 21335
rect 5273 21097 5307 21131
rect 7389 21097 7423 21131
rect 8033 21097 8067 21131
rect 8723 21097 8757 21131
rect 6790 21029 6824 21063
rect 9505 21029 9539 21063
rect 10609 21029 10643 21063
rect 13829 21029 13863 21063
rect 14381 21029 14415 21063
rect 15945 21029 15979 21063
rect 16037 21029 16071 21063
rect 17509 21029 17543 21063
rect 17601 21029 17635 21063
rect 4445 20961 4479 20995
rect 5524 20961 5558 20995
rect 8652 20961 8686 20995
rect 11161 20961 11195 20995
rect 12081 20961 12115 20995
rect 12633 20961 12667 20995
rect 6285 20893 6319 20927
rect 6469 20893 6503 20927
rect 10517 20893 10551 20927
rect 12817 20893 12851 20927
rect 13277 20893 13311 20927
rect 13737 20893 13771 20927
rect 16221 20893 16255 20927
rect 17785 20893 17819 20927
rect 4629 20757 4663 20791
rect 5595 20757 5629 20791
rect 7665 20757 7699 20791
rect 9045 20757 9079 20791
rect 10149 20757 10183 20791
rect 15761 20757 15795 20791
rect 16865 20757 16899 20791
rect 3341 20553 3375 20587
rect 7757 20553 7791 20587
rect 8493 20553 8527 20587
rect 9965 20553 9999 20587
rect 11161 20553 11195 20587
rect 12081 20553 12115 20587
rect 12633 20553 12667 20587
rect 14197 20553 14231 20587
rect 15853 20553 15887 20587
rect 17417 20553 17451 20587
rect 17785 20553 17819 20587
rect 18199 20553 18233 20587
rect 1823 20485 1857 20519
rect 6285 20485 6319 20519
rect 8677 20417 8711 20451
rect 9137 20417 9171 20451
rect 10241 20417 10275 20451
rect 10517 20417 10551 20451
rect 13277 20417 13311 20451
rect 15577 20417 15611 20451
rect 16681 20417 16715 20451
rect 1752 20349 1786 20383
rect 2856 20349 2890 20383
rect 3836 20349 3870 20383
rect 4261 20349 4295 20383
rect 5089 20349 5123 20383
rect 5181 20349 5215 20383
rect 5641 20349 5675 20383
rect 6837 20349 6871 20383
rect 15092 20349 15126 20383
rect 18128 20349 18162 20383
rect 19108 20349 19142 20383
rect 19533 20349 19567 20383
rect 5917 20281 5951 20315
rect 7158 20281 7192 20315
rect 8033 20281 8067 20315
rect 8769 20281 8803 20315
rect 10333 20281 10367 20315
rect 13598 20281 13632 20315
rect 16221 20281 16255 20315
rect 16313 20281 16347 20315
rect 2145 20213 2179 20247
rect 2927 20213 2961 20247
rect 3939 20213 3973 20247
rect 4721 20213 4755 20247
rect 6653 20213 6687 20247
rect 9689 20213 9723 20247
rect 13185 20213 13219 20247
rect 14473 20213 14507 20247
rect 15163 20213 15197 20247
rect 18521 20213 18555 20247
rect 19211 20213 19245 20247
rect 7297 20009 7331 20043
rect 8723 20009 8757 20043
rect 11575 20009 11609 20043
rect 14105 20009 14139 20043
rect 15853 20009 15887 20043
rect 5549 19941 5583 19975
rect 6698 19941 6732 19975
rect 10010 19941 10044 19975
rect 13271 19941 13305 19975
rect 16221 19941 16255 19975
rect 17785 19941 17819 19975
rect 1476 19873 1510 19907
rect 2973 19873 3007 19907
rect 5089 19873 5123 19907
rect 5273 19873 5307 19907
rect 5825 19873 5859 19907
rect 8652 19873 8686 19907
rect 9689 19873 9723 19907
rect 10609 19873 10643 19907
rect 11504 19873 11538 19907
rect 13829 19873 13863 19907
rect 19232 19873 19266 19907
rect 6377 19805 6411 19839
rect 9137 19805 9171 19839
rect 12909 19805 12943 19839
rect 16129 19805 16163 19839
rect 17693 19805 17727 19839
rect 17969 19805 18003 19839
rect 16681 19737 16715 19771
rect 1547 19669 1581 19703
rect 3157 19669 3191 19703
rect 7757 19669 7791 19703
rect 12541 19669 12575 19703
rect 19303 19669 19337 19703
rect 2513 19465 2547 19499
rect 4721 19465 4755 19499
rect 10425 19465 10459 19499
rect 15853 19465 15887 19499
rect 16221 19465 16255 19499
rect 17693 19465 17727 19499
rect 24777 19465 24811 19499
rect 10701 19397 10735 19431
rect 2743 19329 2777 19363
rect 5917 19329 5951 19363
rect 9045 19329 9079 19363
rect 16497 19329 16531 19363
rect 1409 19261 1443 19295
rect 2656 19261 2690 19295
rect 3525 19261 3559 19295
rect 3617 19261 3651 19295
rect 4169 19261 4203 19295
rect 5089 19261 5123 19295
rect 5181 19261 5215 19295
rect 5641 19261 5675 19295
rect 7021 19261 7055 19295
rect 7757 19261 7791 19295
rect 8677 19261 8711 19295
rect 9505 19261 9539 19295
rect 11345 19261 11379 19295
rect 12541 19261 12575 19295
rect 13461 19261 13495 19295
rect 14105 19261 14139 19295
rect 14933 19261 14967 19295
rect 16716 19261 16750 19295
rect 18096 19261 18130 19295
rect 18521 19261 18555 19295
rect 19073 19261 19107 19295
rect 19533 19261 19567 19295
rect 19901 19261 19935 19295
rect 24593 19261 24627 19295
rect 25145 19261 25179 19295
rect 8078 19193 8112 19227
rect 9867 19193 9901 19227
rect 12903 19193 12937 19227
rect 15254 19193 15288 19227
rect 16819 19193 16853 19227
rect 20085 19193 20119 19227
rect 1593 19125 1627 19159
rect 2053 19125 2087 19159
rect 3065 19125 3099 19159
rect 3893 19125 3927 19159
rect 6377 19125 6411 19159
rect 7573 19125 7607 19159
rect 9321 19125 9355 19159
rect 11161 19125 11195 19159
rect 11529 19125 11563 19159
rect 11897 19125 11931 19159
rect 12265 19125 12299 19159
rect 13737 19125 13771 19159
rect 14749 19125 14783 19159
rect 17233 19125 17267 19159
rect 18199 19125 18233 19159
rect 19257 19125 19291 19159
rect 3709 18921 3743 18955
rect 4905 18921 4939 18955
rect 9505 18921 9539 18955
rect 11253 18921 11287 18955
rect 12541 18921 12575 18955
rect 14013 18921 14047 18955
rect 16221 18921 16255 18955
rect 17141 18921 17175 18955
rect 18061 18921 18095 18955
rect 24777 18921 24811 18955
rect 6101 18853 6135 18887
rect 9965 18853 9999 18887
rect 10241 18853 10275 18887
rect 10333 18853 10367 18887
rect 10885 18853 10919 18887
rect 13179 18853 13213 18887
rect 15622 18853 15656 18887
rect 16589 18853 16623 18887
rect 2028 18785 2062 18819
rect 3040 18785 3074 18819
rect 5457 18785 5491 18819
rect 5825 18785 5859 18819
rect 7021 18785 7055 18819
rect 7481 18785 7515 18819
rect 8652 18785 8686 18819
rect 11780 18785 11814 18819
rect 13737 18785 13771 18819
rect 17049 18785 17083 18819
rect 17601 18785 17635 18819
rect 18680 18785 18714 18819
rect 19660 18785 19694 18819
rect 24593 18785 24627 18819
rect 4077 18717 4111 18751
rect 7665 18717 7699 18751
rect 12817 18717 12851 18751
rect 15301 18717 15335 18751
rect 20913 18717 20947 18751
rect 1685 18581 1719 18615
rect 2099 18581 2133 18615
rect 3111 18581 3145 18615
rect 5273 18581 5307 18615
rect 8033 18581 8067 18615
rect 8723 18581 8757 18615
rect 11851 18581 11885 18615
rect 14933 18581 14967 18615
rect 18751 18581 18785 18615
rect 19763 18581 19797 18615
rect 2513 18377 2547 18411
rect 7021 18377 7055 18411
rect 9045 18377 9079 18411
rect 11805 18377 11839 18411
rect 15853 18377 15887 18411
rect 20085 18377 20119 18411
rect 6653 18309 6687 18343
rect 16589 18309 16623 18343
rect 24593 18309 24627 18343
rect 8033 18241 8067 18275
rect 10333 18241 10367 18275
rect 11529 18241 11563 18275
rect 14749 18241 14783 18275
rect 16037 18241 16071 18275
rect 18751 18241 18785 18275
rect 20453 18241 20487 18275
rect 1660 18173 1694 18207
rect 3525 18173 3559 18207
rect 3893 18173 3927 18207
rect 4169 18173 4203 18207
rect 5089 18173 5123 18207
rect 5365 18173 5399 18207
rect 5733 18173 5767 18207
rect 8677 18173 8711 18207
rect 9229 18173 9263 18207
rect 9781 18173 9815 18207
rect 10977 18173 11011 18207
rect 11253 18173 11287 18207
rect 12449 18173 12483 18207
rect 12909 18173 12943 18207
rect 14013 18173 14047 18207
rect 14473 18173 14507 18207
rect 18648 18173 18682 18207
rect 19441 18173 19475 18207
rect 19660 18173 19694 18207
rect 2145 18105 2179 18139
rect 5917 18105 5951 18139
rect 7389 18105 7423 18139
rect 7481 18105 7515 18139
rect 9965 18105 9999 18139
rect 13185 18105 13219 18139
rect 16129 18105 16163 18139
rect 1731 18037 1765 18071
rect 2605 18037 2639 18071
rect 3157 18037 3191 18071
rect 3893 18037 3927 18071
rect 6285 18037 6319 18071
rect 10701 18037 10735 18071
rect 12265 18037 12299 18071
rect 13461 18037 13495 18071
rect 13829 18037 13863 18071
rect 15301 18037 15335 18071
rect 17049 18037 17083 18071
rect 17509 18037 17543 18071
rect 19165 18037 19199 18071
rect 19763 18037 19797 18071
rect 20637 18037 20671 18071
rect 21649 18037 21683 18071
rect 3709 17833 3743 17867
rect 5549 17833 5583 17867
rect 6929 17833 6963 17867
rect 7389 17833 7423 17867
rect 9321 17833 9355 17867
rect 10149 17833 10183 17867
rect 13093 17833 13127 17867
rect 16497 17833 16531 17867
rect 18429 17833 18463 17867
rect 6330 17765 6364 17799
rect 7941 17765 7975 17799
rect 8493 17765 8527 17799
rect 10609 17765 10643 17799
rect 14289 17765 14323 17799
rect 16037 17765 16071 17799
rect 16951 17765 16985 17799
rect 1961 17697 1995 17731
rect 4721 17697 4755 17731
rect 4997 17697 5031 17731
rect 11989 17697 12023 17731
rect 12449 17697 12483 17731
rect 13553 17697 13587 17731
rect 14013 17697 14047 17731
rect 15644 17697 15678 17731
rect 16589 17697 16623 17731
rect 18613 17697 18647 17731
rect 18797 17697 18831 17731
rect 20948 17697 20982 17731
rect 22268 17697 22302 17731
rect 23280 17697 23314 17731
rect 2973 17629 3007 17663
rect 5181 17629 5215 17663
rect 6009 17629 6043 17663
rect 7849 17629 7883 17663
rect 10517 17629 10551 17663
rect 12541 17629 12575 17663
rect 11069 17561 11103 17595
rect 2145 17493 2179 17527
rect 4353 17493 4387 17527
rect 14565 17493 14599 17527
rect 15715 17493 15749 17527
rect 17509 17493 17543 17527
rect 18153 17493 18187 17527
rect 21051 17493 21085 17527
rect 22339 17493 22373 17527
rect 23351 17493 23385 17527
rect 1593 17289 1627 17323
rect 4537 17289 4571 17323
rect 5733 17289 5767 17323
rect 7757 17289 7791 17323
rect 8033 17289 8067 17323
rect 21097 17289 21131 17323
rect 24777 17289 24811 17323
rect 10977 17221 11011 17255
rect 11713 17221 11747 17255
rect 17049 17221 17083 17255
rect 3157 17153 3191 17187
rect 4721 17153 4755 17187
rect 6837 17153 6871 17187
rect 8585 17153 8619 17187
rect 10425 17153 10459 17187
rect 13553 17153 13587 17187
rect 14381 17153 14415 17187
rect 16129 17153 16163 17187
rect 18429 17153 18463 17187
rect 1409 17085 1443 17119
rect 2605 17085 2639 17119
rect 3684 17085 3718 17119
rect 4077 17085 4111 17119
rect 9965 17085 9999 17119
rect 12817 17085 12851 17119
rect 13277 17085 13311 17119
rect 17785 17085 17819 17119
rect 19692 17085 19726 17119
rect 20704 17085 20738 17119
rect 21465 17085 21499 17119
rect 21716 17085 21750 17119
rect 22109 17085 22143 17119
rect 24593 17085 24627 17119
rect 25145 17085 25179 17119
rect 4813 17017 4847 17051
rect 5365 17017 5399 17051
rect 7158 17017 7192 17051
rect 8906 17017 8940 17051
rect 9873 17017 9907 17051
rect 10241 17017 10275 17051
rect 10517 17017 10551 17051
rect 14197 17017 14231 17051
rect 14702 17017 14736 17051
rect 15945 17017 15979 17051
rect 16450 17017 16484 17051
rect 17325 17017 17359 17051
rect 18153 17017 18187 17051
rect 18245 17017 18279 17051
rect 20177 17017 20211 17051
rect 2053 16949 2087 16983
rect 2421 16949 2455 16983
rect 2789 16949 2823 16983
rect 3755 16949 3789 16983
rect 6101 16949 6135 16983
rect 6561 16949 6595 16983
rect 8401 16949 8435 16983
rect 9505 16949 9539 16983
rect 9965 16949 9999 16983
rect 11989 16949 12023 16983
rect 12633 16949 12667 16983
rect 13829 16949 13863 16983
rect 15301 16949 15335 16983
rect 15669 16949 15703 16983
rect 19073 16949 19107 16983
rect 19763 16949 19797 16983
rect 20775 16949 20809 16983
rect 21787 16949 21821 16983
rect 22569 16949 22603 16983
rect 23305 16949 23339 16983
rect 3111 16745 3145 16779
rect 4997 16745 5031 16779
rect 6837 16745 6871 16779
rect 7573 16745 7607 16779
rect 8677 16745 8711 16779
rect 11069 16745 11103 16779
rect 14381 16745 14415 16779
rect 16681 16745 16715 16779
rect 18613 16745 18647 16779
rect 21051 16745 21085 16779
rect 4398 16677 4432 16711
rect 5273 16677 5307 16711
rect 6009 16677 6043 16711
rect 7849 16677 7883 16711
rect 9781 16677 9815 16711
rect 9873 16677 9907 16711
rect 10793 16677 10827 16711
rect 11437 16677 11471 16711
rect 12817 16677 12851 16711
rect 13506 16677 13540 16711
rect 15761 16677 15795 16711
rect 17785 16677 17819 16711
rect 19349 16677 19383 16711
rect 19901 16677 19935 16711
rect 25099 16677 25133 16711
rect 1961 16609 1995 16643
rect 3040 16609 3074 16643
rect 4077 16609 4111 16643
rect 15117 16609 15151 16643
rect 20980 16609 21014 16643
rect 21992 16609 22026 16643
rect 22972 16609 23006 16643
rect 23075 16609 23109 16643
rect 23949 16609 23983 16643
rect 25012 16609 25046 16643
rect 5917 16541 5951 16575
rect 6561 16541 6595 16575
rect 7757 16541 7791 16575
rect 8033 16541 8067 16575
rect 10057 16541 10091 16575
rect 11345 16541 11379 16575
rect 11713 16541 11747 16575
rect 13185 16541 13219 16575
rect 15669 16541 15703 16575
rect 17509 16541 17543 16575
rect 17693 16541 17727 16575
rect 17969 16541 18003 16575
rect 19257 16541 19291 16575
rect 14105 16473 14139 16507
rect 16221 16473 16255 16507
rect 2145 16405 2179 16439
rect 22063 16405 22097 16439
rect 1593 16201 1627 16235
rect 5089 16201 5123 16235
rect 5917 16201 5951 16235
rect 6193 16201 6227 16235
rect 6653 16201 6687 16235
rect 7205 16201 7239 16235
rect 7573 16201 7607 16235
rect 9045 16201 9079 16235
rect 10793 16201 10827 16235
rect 11345 16201 11379 16235
rect 14013 16201 14047 16235
rect 15669 16201 15703 16235
rect 15853 16201 15887 16235
rect 17509 16201 17543 16235
rect 20729 16201 20763 16235
rect 24777 16201 24811 16235
rect 15485 16133 15519 16167
rect 2053 16065 2087 16099
rect 4077 16065 4111 16099
rect 7757 16065 7791 16099
rect 8401 16065 8435 16099
rect 14657 16065 14691 16099
rect 14933 16065 14967 16099
rect 16497 16065 16531 16099
rect 16773 16065 16807 16099
rect 18153 16065 18187 16099
rect 19717 16065 19751 16099
rect 19993 16065 20027 16099
rect 21097 16065 21131 16099
rect 1409 15997 1443 16031
rect 2513 15997 2547 16031
rect 2881 15997 2915 16031
rect 3157 15997 3191 16031
rect 4169 15997 4203 16031
rect 9873 15997 9907 16031
rect 13093 15997 13127 16031
rect 14289 15997 14323 16031
rect 15669 15997 15703 16031
rect 16221 15997 16255 16031
rect 21240 15997 21274 16031
rect 22236 15997 22270 16031
rect 23029 15997 23063 16031
rect 24593 15997 24627 16031
rect 25145 15997 25179 16031
rect 3341 15929 3375 15963
rect 3709 15929 3743 15963
rect 4531 15929 4565 15963
rect 7849 15929 7883 15963
rect 10194 15929 10228 15963
rect 13414 15929 13448 15963
rect 15025 15929 15059 15963
rect 16589 15929 16623 15963
rect 18245 15929 18279 15963
rect 18797 15929 18831 15963
rect 19809 15929 19843 15963
rect 21327 15929 21361 15963
rect 22109 15929 22143 15963
rect 5365 15861 5399 15895
rect 9321 15861 9355 15895
rect 9781 15861 9815 15895
rect 11621 15861 11655 15895
rect 12265 15861 12299 15895
rect 13001 15861 13035 15895
rect 17785 15861 17819 15895
rect 19073 15861 19107 15895
rect 19441 15861 19475 15895
rect 21741 15861 21775 15895
rect 22339 15861 22373 15895
rect 25513 15861 25547 15895
rect 1593 15657 1627 15691
rect 4261 15657 4295 15691
rect 5273 15657 5307 15691
rect 7481 15657 7515 15691
rect 8125 15657 8159 15691
rect 9505 15657 9539 15691
rect 12541 15657 12575 15691
rect 12633 15657 12667 15691
rect 14841 15657 14875 15691
rect 16497 15657 16531 15691
rect 18245 15657 18279 15691
rect 18613 15657 18647 15691
rect 19717 15657 19751 15691
rect 6882 15589 6916 15623
rect 12173 15589 12207 15623
rect 1409 15521 1443 15555
rect 2973 15521 3007 15555
rect 5181 15521 5215 15555
rect 5457 15521 5491 15555
rect 6561 15521 6595 15555
rect 8620 15521 8654 15555
rect 8723 15521 8757 15555
rect 9873 15521 9907 15555
rect 10333 15521 10367 15555
rect 11437 15521 11471 15555
rect 11989 15521 12023 15555
rect 10609 15453 10643 15487
rect 2697 15385 2731 15419
rect 3157 15385 3191 15419
rect 13322 15589 13356 15623
rect 15485 15589 15519 15623
rect 17325 15589 17359 15623
rect 17877 15589 17911 15623
rect 18889 15589 18923 15623
rect 19441 15589 19475 15623
rect 21189 15589 21223 15623
rect 21281 15589 21315 15623
rect 22728 15521 22762 15555
rect 23740 15521 23774 15555
rect 24752 15521 24786 15555
rect 12909 15453 12943 15487
rect 13001 15453 13035 15487
rect 15393 15453 15427 15487
rect 15669 15453 15703 15487
rect 17233 15453 17267 15487
rect 18797 15453 18831 15487
rect 22109 15453 22143 15487
rect 21741 15385 21775 15419
rect 1961 15317 1995 15351
rect 3617 15317 3651 15351
rect 4629 15317 4663 15351
rect 6377 15317 6411 15351
rect 7849 15317 7883 15351
rect 12633 15317 12667 15351
rect 13921 15317 13955 15351
rect 22799 15317 22833 15351
rect 23811 15317 23845 15351
rect 24823 15317 24857 15351
rect 1961 15113 1995 15147
rect 2421 15113 2455 15147
rect 4629 15113 4663 15147
rect 8033 15113 8067 15147
rect 9873 15113 9907 15147
rect 10609 15113 10643 15147
rect 12173 15113 12207 15147
rect 12587 15113 12621 15147
rect 12909 15113 12943 15147
rect 14749 15113 14783 15147
rect 16773 15113 16807 15147
rect 19073 15113 19107 15147
rect 21741 15113 21775 15147
rect 22845 15113 22879 15147
rect 1777 15045 1811 15079
rect 1593 14909 1627 14943
rect 10241 15045 10275 15079
rect 15945 15045 15979 15079
rect 17693 15045 17727 15079
rect 17785 15045 17819 15079
rect 4353 14977 4387 15011
rect 5917 14977 5951 15011
rect 6837 14977 6871 15011
rect 8953 14977 8987 15011
rect 11529 14977 11563 15011
rect 13829 14977 13863 15011
rect 14105 14977 14139 15011
rect 15393 14977 15427 15011
rect 16405 14977 16439 15011
rect 17417 14977 17451 15011
rect 2672 14909 2706 14943
rect 3157 14909 3191 14943
rect 3893 14909 3927 14943
rect 4169 14909 4203 14943
rect 5181 14909 5215 14943
rect 5641 14909 5675 14943
rect 10793 14909 10827 14943
rect 11345 14909 11379 14943
rect 12516 14909 12550 14943
rect 17008 14909 17042 14943
rect 1961 14841 1995 14875
rect 2053 14841 2087 14875
rect 3525 14841 3559 14875
rect 7158 14841 7192 14875
rect 8677 14841 8711 14875
rect 8769 14841 8803 14875
rect 11805 14841 11839 14875
rect 13921 14841 13955 14875
rect 15209 14841 15243 14875
rect 15485 14841 15519 14875
rect 17095 14841 17129 14875
rect 18153 14977 18187 15011
rect 18797 14977 18831 15011
rect 22109 14977 22143 15011
rect 20545 14909 20579 14943
rect 21465 14909 21499 14943
rect 22344 14909 22378 14943
rect 23121 14909 23155 14943
rect 23740 14909 23774 14943
rect 24133 14909 24167 14943
rect 18245 14841 18279 14875
rect 20866 14841 20900 14875
rect 24685 14841 24719 14875
rect 2743 14773 2777 14807
rect 5089 14773 5123 14807
rect 6285 14773 6319 14807
rect 6561 14773 6595 14807
rect 7757 14773 7791 14807
rect 8493 14773 8527 14807
rect 13277 14773 13311 14807
rect 17693 14773 17727 14807
rect 19441 14773 19475 14807
rect 20361 14773 20395 14807
rect 22431 14773 22465 14807
rect 23811 14773 23845 14807
rect 24501 14773 24535 14807
rect 25145 14773 25179 14807
rect 1593 14569 1627 14603
rect 3111 14569 3145 14603
rect 4169 14569 4203 14603
rect 5181 14569 5215 14603
rect 5549 14569 5583 14603
rect 8953 14569 8987 14603
rect 9965 14569 9999 14603
rect 10885 14569 10919 14603
rect 13829 14569 13863 14603
rect 17233 14569 17267 14603
rect 20637 14569 20671 14603
rect 22569 14569 22603 14603
rect 24777 14569 24811 14603
rect 3709 14501 3743 14535
rect 7757 14501 7791 14535
rect 8585 14501 8619 14535
rect 11989 14501 12023 14535
rect 13001 14501 13035 14535
rect 13553 14501 13587 14535
rect 15485 14501 15519 14535
rect 17601 14501 17635 14535
rect 17693 14501 17727 14535
rect 19394 14501 19428 14535
rect 21097 14501 21131 14535
rect 1409 14433 1443 14467
rect 3040 14433 3074 14467
rect 4169 14433 4203 14467
rect 4629 14433 4663 14467
rect 6101 14433 6135 14467
rect 6285 14433 6319 14467
rect 9781 14433 9815 14467
rect 10149 14433 10183 14467
rect 11253 14433 11287 14467
rect 11713 14433 11747 14467
rect 19993 14433 20027 14467
rect 22753 14433 22787 14467
rect 22937 14433 22971 14467
rect 24593 14433 24627 14467
rect 6377 14365 6411 14399
rect 7665 14365 7699 14399
rect 8033 14365 8067 14399
rect 12909 14365 12943 14399
rect 14197 14365 14231 14399
rect 15393 14365 15427 14399
rect 16037 14365 16071 14399
rect 18245 14365 18279 14399
rect 19073 14365 19107 14399
rect 21005 14365 21039 14399
rect 21465 14365 21499 14399
rect 15025 14297 15059 14331
rect 7205 14229 7239 14263
rect 9505 14229 9539 14263
rect 21925 14229 21959 14263
rect 22293 14229 22327 14263
rect 23765 14229 23799 14263
rect 1685 14025 1719 14059
rect 2053 14025 2087 14059
rect 5641 14025 5675 14059
rect 6101 14025 6135 14059
rect 6377 14025 6411 14059
rect 8125 14025 8159 14059
rect 8815 14025 8849 14059
rect 9781 14025 9815 14059
rect 11253 14025 11287 14059
rect 11713 14025 11747 14059
rect 14013 14025 14047 14059
rect 19073 14025 19107 14059
rect 21005 14025 21039 14059
rect 24685 14025 24719 14059
rect 25375 14025 25409 14059
rect 3801 13957 3835 13991
rect 13369 13957 13403 13991
rect 13645 13957 13679 13991
rect 14841 13957 14875 13991
rect 14933 13957 14967 13991
rect 16129 13957 16163 13991
rect 16865 13957 16899 13991
rect 17877 13957 17911 13991
rect 20453 13957 20487 13991
rect 2789 13889 2823 13923
rect 4169 13889 4203 13923
rect 7205 13889 7239 13923
rect 10057 13889 10091 13923
rect 12449 13889 12483 13923
rect 14657 13889 14691 13923
rect 15209 13889 15243 13923
rect 15853 13889 15887 13923
rect 17095 13889 17129 13923
rect 18153 13889 18187 13923
rect 19901 13889 19935 13923
rect 21465 13889 21499 13923
rect 21741 13889 21775 13923
rect 1869 13821 1903 13855
rect 2881 13821 2915 13855
rect 4537 13821 4571 13855
rect 4721 13821 4755 13855
rect 5181 13821 5215 13855
rect 7849 13821 7883 13855
rect 8744 13821 8778 13855
rect 10701 13821 10735 13855
rect 14841 13821 14875 13855
rect 16992 13821 17026 13855
rect 17417 13821 17451 13855
rect 22569 13821 22603 13855
rect 23765 13821 23799 13855
rect 24133 13821 24167 13855
rect 25304 13821 25338 13855
rect 25697 13821 25731 13855
rect 2421 13753 2455 13787
rect 3243 13753 3277 13787
rect 5365 13753 5399 13787
rect 7297 13753 7331 13787
rect 10149 13753 10183 13787
rect 12770 13753 12804 13787
rect 15301 13753 15335 13787
rect 18245 13753 18279 13787
rect 18797 13753 18831 13787
rect 19717 13753 19751 13787
rect 19993 13753 20027 13787
rect 21557 13753 21591 13787
rect 22937 13753 22971 13787
rect 23397 13753 23431 13787
rect 9229 13685 9263 13719
rect 12173 13685 12207 13719
rect 23765 13685 23799 13719
rect 3341 13481 3375 13515
rect 3893 13481 3927 13515
rect 6193 13481 6227 13515
rect 7205 13481 7239 13515
rect 7481 13481 7515 13515
rect 9137 13481 9171 13515
rect 9505 13481 9539 13515
rect 10609 13481 10643 13515
rect 11621 13481 11655 13515
rect 12449 13481 12483 13515
rect 13553 13481 13587 13515
rect 15025 13481 15059 13515
rect 17969 13481 18003 13515
rect 18245 13481 18279 13515
rect 19901 13481 19935 13515
rect 20729 13481 20763 13515
rect 2421 13413 2455 13447
rect 4439 13413 4473 13447
rect 6606 13413 6640 13447
rect 8217 13413 8251 13447
rect 10010 13413 10044 13447
rect 12954 13413 12988 13447
rect 15485 13413 15519 13447
rect 16037 13413 16071 13447
rect 17049 13413 17083 13447
rect 18613 13413 18647 13447
rect 19533 13413 19567 13447
rect 21557 13413 21591 13447
rect 23121 13413 23155 13447
rect 6285 13345 6319 13379
rect 11437 13345 11471 13379
rect 12633 13345 12667 13379
rect 24536 13345 24570 13379
rect 2329 13277 2363 13311
rect 4077 13277 4111 13311
rect 8125 13277 8159 13311
rect 8401 13277 8435 13311
rect 9689 13277 9723 13311
rect 15393 13277 15427 13311
rect 16957 13277 16991 13311
rect 17325 13277 17359 13311
rect 18521 13277 18555 13311
rect 18797 13277 18831 13311
rect 21465 13277 21499 13311
rect 23029 13277 23063 13311
rect 24639 13277 24673 13311
rect 2881 13209 2915 13243
rect 22017 13209 22051 13243
rect 23581 13209 23615 13243
rect 1685 13141 1719 13175
rect 4997 13141 5031 13175
rect 7941 13141 7975 13175
rect 13829 13141 13863 13175
rect 21097 13141 21131 13175
rect 1685 12937 1719 12971
rect 2697 12937 2731 12971
rect 5181 12937 5215 12971
rect 8401 12937 8435 12971
rect 8769 12937 8803 12971
rect 10793 12937 10827 12971
rect 12173 12937 12207 12971
rect 12679 12937 12713 12971
rect 15393 12937 15427 12971
rect 22017 12937 22051 12971
rect 22477 12937 22511 12971
rect 23397 12937 23431 12971
rect 24317 12937 24351 12971
rect 24869 12937 24903 12971
rect 25605 12937 25639 12971
rect 1961 12869 1995 12903
rect 5917 12869 5951 12903
rect 7757 12869 7791 12903
rect 11161 12869 11195 12903
rect 13369 12869 13403 12903
rect 18889 12869 18923 12903
rect 3341 12801 3375 12835
rect 4537 12801 4571 12835
rect 8125 12801 8159 12835
rect 9873 12801 9907 12835
rect 11483 12801 11517 12835
rect 13645 12801 13679 12835
rect 14105 12801 14139 12835
rect 16129 12801 16163 12835
rect 18337 12801 18371 12835
rect 20821 12801 20855 12835
rect 23121 12801 23155 12835
rect 24501 12869 24535 12903
rect 1777 12733 1811 12767
rect 2329 12733 2363 12767
rect 2789 12733 2823 12767
rect 5733 12733 5767 12767
rect 6837 12733 6871 12767
rect 8585 12733 8619 12767
rect 9045 12733 9079 12767
rect 11380 12733 11414 12767
rect 11805 12733 11839 12767
rect 12608 12733 12642 12767
rect 13001 12733 13035 12767
rect 19844 12733 19878 12767
rect 20269 12733 20303 12767
rect 22636 12733 22670 12767
rect 24108 12733 24142 12767
rect 24317 12733 24351 12767
rect 25104 12733 25138 12767
rect 3709 12665 3743 12699
rect 3893 12665 3927 12699
rect 3985 12665 4019 12699
rect 5641 12665 5675 12699
rect 6377 12665 6411 12699
rect 7158 12665 7192 12699
rect 9689 12665 9723 12699
rect 9965 12665 9999 12699
rect 10517 12665 10551 12699
rect 13737 12665 13771 12699
rect 14933 12665 14967 12699
rect 15853 12665 15887 12699
rect 15945 12665 15979 12699
rect 16865 12665 16899 12699
rect 17877 12665 17911 12699
rect 18429 12665 18463 12699
rect 19257 12665 19291 12699
rect 20729 12665 20763 12699
rect 21142 12665 21176 12699
rect 25191 12665 25225 12699
rect 2973 12597 3007 12631
rect 4905 12597 4939 12631
rect 14565 12597 14599 12631
rect 17233 12597 17267 12631
rect 19947 12597 19981 12631
rect 21741 12597 21775 12631
rect 22707 12597 22741 12631
rect 24179 12597 24213 12631
rect 3893 12393 3927 12427
rect 4169 12393 4203 12427
rect 9965 12393 9999 12427
rect 10241 12393 10275 12427
rect 12449 12393 12483 12427
rect 13461 12393 13495 12427
rect 13737 12393 13771 12427
rect 16405 12393 16439 12427
rect 18153 12393 18187 12427
rect 18521 12393 18555 12427
rect 21833 12393 21867 12427
rect 24317 12393 24351 12427
rect 3157 12325 3191 12359
rect 8769 12325 8803 12359
rect 10609 12325 10643 12359
rect 10701 12325 10735 12359
rect 12903 12325 12937 12359
rect 15485 12325 15519 12359
rect 16037 12325 16071 12359
rect 17595 12325 17629 12359
rect 19441 12325 19475 12359
rect 19993 12325 20027 12359
rect 21234 12325 21268 12359
rect 22845 12325 22879 12359
rect 1409 12257 1443 12291
rect 2421 12257 2455 12291
rect 2881 12257 2915 12291
rect 4077 12257 4111 12291
rect 4629 12257 4663 12291
rect 5917 12257 5951 12291
rect 6101 12257 6135 12291
rect 8309 12257 8343 12291
rect 8585 12257 8619 12291
rect 18797 12257 18831 12291
rect 22109 12257 22143 12291
rect 24501 12257 24535 12291
rect 24777 12257 24811 12291
rect 6377 12189 6411 12223
rect 7205 12189 7239 12223
rect 12541 12189 12575 12223
rect 15393 12189 15427 12223
rect 17233 12189 17267 12223
rect 19349 12189 19383 12223
rect 20913 12189 20947 12223
rect 22753 12189 22787 12223
rect 23029 12189 23063 12223
rect 1593 12121 1627 12155
rect 11161 12121 11195 12155
rect 1961 12053 1995 12087
rect 2329 12053 2363 12087
rect 5089 12053 5123 12087
rect 6929 12053 6963 12087
rect 7941 12053 7975 12087
rect 14105 12053 14139 12087
rect 20729 12053 20763 12087
rect 23673 12053 23707 12087
rect 1685 11849 1719 11883
rect 3249 11849 3283 11883
rect 3893 11849 3927 11883
rect 5733 11849 5767 11883
rect 7757 11849 7791 11883
rect 11161 11849 11195 11883
rect 16957 11849 16991 11883
rect 18797 11849 18831 11883
rect 21649 11849 21683 11883
rect 22615 11849 22649 11883
rect 25421 11849 25455 11883
rect 2513 11781 2547 11815
rect 6101 11781 6135 11815
rect 8953 11781 8987 11815
rect 18429 11781 18463 11815
rect 19809 11781 19843 11815
rect 22385 11781 22419 11815
rect 4261 11713 4295 11747
rect 4445 11713 4479 11747
rect 7941 11713 7975 11747
rect 8585 11713 8619 11747
rect 9597 11713 9631 11747
rect 15945 11713 15979 11747
rect 16221 11713 16255 11747
rect 17325 11713 17359 11747
rect 20729 11713 20763 11747
rect 21925 11713 21959 11747
rect 2329 11645 2363 11679
rect 3341 11645 3375 11679
rect 4353 11645 4387 11679
rect 4629 11645 4663 11679
rect 6837 11645 6871 11679
rect 7297 11645 7331 11679
rect 11345 11645 11379 11679
rect 11805 11645 11839 11679
rect 12541 11645 12575 11679
rect 13001 11645 13035 11679
rect 13553 11645 13587 11679
rect 14105 11645 14139 11679
rect 15025 11645 15059 11679
rect 15669 11645 15703 11679
rect 18889 11645 18923 11679
rect 22512 11645 22546 11679
rect 22937 11645 22971 11679
rect 23765 11645 23799 11679
rect 24133 11645 24167 11679
rect 25237 11645 25271 11679
rect 25789 11645 25823 11679
rect 5089 11577 5123 11611
rect 8033 11577 8067 11611
rect 9918 11577 9952 11611
rect 12173 11577 12207 11611
rect 13277 11577 13311 11611
rect 14426 11577 14460 11611
rect 16037 11577 16071 11611
rect 19210 11577 19244 11611
rect 20177 11577 20211 11611
rect 20545 11577 20579 11611
rect 21050 11577 21084 11611
rect 24685 11577 24719 11611
rect 2237 11509 2271 11543
rect 2881 11509 2915 11543
rect 3525 11509 3559 11543
rect 7021 11509 7055 11543
rect 9413 11509 9447 11543
rect 10517 11509 10551 11543
rect 10885 11509 10919 11543
rect 11529 11509 11563 11543
rect 13921 11509 13955 11543
rect 15301 11509 15335 11543
rect 17693 11509 17727 11543
rect 23397 11509 23431 11543
rect 23765 11509 23799 11543
rect 25145 11509 25179 11543
rect 1593 11305 1627 11339
rect 2329 11305 2363 11339
rect 4905 11305 4939 11339
rect 7389 11305 7423 11339
rect 8493 11305 8527 11339
rect 12449 11305 12483 11339
rect 12725 11305 12759 11339
rect 13093 11305 13127 11339
rect 14289 11305 14323 11339
rect 18245 11305 18279 11339
rect 18889 11305 18923 11339
rect 21005 11305 21039 11339
rect 22753 11305 22787 11339
rect 24961 11305 24995 11339
rect 3801 11237 3835 11271
rect 4261 11237 4295 11271
rect 7935 11237 7969 11271
rect 10885 11237 10919 11271
rect 13731 11237 13765 11271
rect 15577 11237 15611 11271
rect 15669 11237 15703 11271
rect 17646 11237 17680 11271
rect 18613 11237 18647 11271
rect 19993 11237 20027 11271
rect 23397 11237 23431 11271
rect 23489 11237 23523 11271
rect 1409 11169 1443 11203
rect 2421 11169 2455 11203
rect 2697 11169 2731 11203
rect 4445 11169 4479 11203
rect 4721 11169 4755 11203
rect 6009 11169 6043 11203
rect 6469 11169 6503 11203
rect 9689 11169 9723 11203
rect 12265 11169 12299 11203
rect 13369 11169 13403 11203
rect 15025 11169 15059 11203
rect 17325 11169 17359 11203
rect 19441 11169 19475 11203
rect 19717 11169 19751 11203
rect 20913 11169 20947 11203
rect 21327 11169 21361 11203
rect 24869 11169 24903 11203
rect 25329 11169 25363 11203
rect 2513 11101 2547 11135
rect 2881 11101 2915 11135
rect 6745 11101 6779 11135
rect 7573 11101 7607 11135
rect 10793 11101 10827 11135
rect 11069 11101 11103 11135
rect 12173 11101 12207 11135
rect 16037 11101 16071 11135
rect 23673 11101 23707 11135
rect 1869 11033 1903 11067
rect 4537 11033 4571 11067
rect 9873 11033 9907 11067
rect 3525 10965 3559 10999
rect 20545 10965 20579 10999
rect 22109 10965 22143 10999
rect 24317 10965 24351 10999
rect 1685 10761 1719 10795
rect 3249 10761 3283 10795
rect 4813 10761 4847 10795
rect 5549 10761 5583 10795
rect 6561 10761 6595 10795
rect 7205 10761 7239 10795
rect 7665 10761 7699 10795
rect 10885 10761 10919 10795
rect 11253 10761 11287 10795
rect 13553 10761 13587 10795
rect 14105 10761 14139 10795
rect 15485 10761 15519 10795
rect 15853 10761 15887 10795
rect 17785 10761 17819 10795
rect 21557 10761 21591 10795
rect 25375 10761 25409 10795
rect 2329 10693 2363 10727
rect 17417 10693 17451 10727
rect 21833 10693 21867 10727
rect 2973 10625 3007 10659
rect 6193 10625 6227 10659
rect 7849 10625 7883 10659
rect 8769 10625 8803 10659
rect 10517 10625 10551 10659
rect 12541 10625 12575 10659
rect 2237 10557 2271 10591
rect 2513 10557 2547 10591
rect 3617 10557 3651 10591
rect 4445 10557 4479 10591
rect 5733 10557 5767 10591
rect 8493 10557 8527 10591
rect 9321 10557 9355 10591
rect 11069 10557 11103 10591
rect 11529 10557 11563 10591
rect 14289 10557 14323 10591
rect 16037 10557 16071 10591
rect 16497 10557 16531 10591
rect 18061 10557 18095 10591
rect 18521 10557 18555 10591
rect 20453 10557 20487 10591
rect 21005 10557 21039 10591
rect 22293 10557 22327 10591
rect 22477 10557 22511 10591
rect 25304 10557 25338 10591
rect 26065 10557 26099 10591
rect 2145 10489 2179 10523
rect 7941 10489 7975 10523
rect 9229 10489 9263 10523
rect 9642 10489 9676 10523
rect 12633 10489 12667 10523
rect 13185 10489 13219 10523
rect 14610 10489 14644 10523
rect 19717 10489 19751 10523
rect 21189 10489 21223 10523
rect 23765 10489 23799 10523
rect 23857 10489 23891 10523
rect 24409 10489 24443 10523
rect 4261 10421 4295 10455
rect 5181 10421 5215 10455
rect 5917 10421 5951 10455
rect 10241 10421 10275 10455
rect 12173 10421 12207 10455
rect 15209 10421 15243 10455
rect 16129 10421 16163 10455
rect 18153 10421 18187 10455
rect 19349 10421 19383 10455
rect 20361 10421 20395 10455
rect 22109 10421 22143 10455
rect 23029 10421 23063 10455
rect 23397 10421 23431 10455
rect 24961 10421 24995 10455
rect 25697 10421 25731 10455
rect 5273 10217 5307 10251
rect 7849 10217 7883 10251
rect 11253 10217 11287 10251
rect 12127 10217 12161 10251
rect 12541 10217 12575 10251
rect 12909 10217 12943 10251
rect 14381 10217 14415 10251
rect 15025 10217 15059 10251
rect 16313 10217 16347 10251
rect 17233 10217 17267 10251
rect 18337 10217 18371 10251
rect 21051 10217 21085 10251
rect 21741 10217 21775 10251
rect 22845 10217 22879 10251
rect 23397 10217 23431 10251
rect 2237 10149 2271 10183
rect 3157 10149 3191 10183
rect 4353 10149 4387 10183
rect 8769 10149 8803 10183
rect 9321 10149 9355 10183
rect 10425 10149 10459 10183
rect 10977 10149 11011 10183
rect 13185 10149 13219 10183
rect 17509 10149 17543 10183
rect 22246 10149 22280 10183
rect 23857 10149 23891 10183
rect 24409 10149 24443 10183
rect 1409 10081 1443 10115
rect 2421 10081 2455 10115
rect 2697 10081 2731 10115
rect 3525 10081 3559 10115
rect 4813 10081 4847 10115
rect 5089 10081 5123 10115
rect 6382 10081 6416 10115
rect 6653 10081 6687 10115
rect 8033 10081 8067 10115
rect 8493 10081 8527 10115
rect 12024 10081 12058 10115
rect 15577 10081 15611 10115
rect 15761 10081 15795 10115
rect 18889 10081 18923 10115
rect 19349 10081 19383 10115
rect 20980 10081 21014 10115
rect 25237 10081 25271 10115
rect 6929 10013 6963 10047
rect 10333 10013 10367 10047
rect 13093 10013 13127 10047
rect 13369 10013 13403 10047
rect 15853 10013 15887 10047
rect 17417 10013 17451 10047
rect 18061 10013 18095 10047
rect 19441 10013 19475 10047
rect 21925 10013 21959 10047
rect 23765 10013 23799 10047
rect 2513 9945 2547 9979
rect 4721 9945 4755 9979
rect 4905 9945 4939 9979
rect 6285 9945 6319 9979
rect 6469 9945 6503 9979
rect 1593 9877 1627 9911
rect 1961 9877 1995 9911
rect 3893 9877 3927 9911
rect 16681 9877 16715 9911
rect 19901 9877 19935 9911
rect 20545 9877 20579 9911
rect 25421 9877 25455 9911
rect 6377 9673 6411 9707
rect 8033 9673 8067 9707
rect 8401 9673 8435 9707
rect 9689 9673 9723 9707
rect 10057 9673 10091 9707
rect 11989 9673 12023 9707
rect 12909 9673 12943 9707
rect 17417 9673 17451 9707
rect 20269 9673 20303 9707
rect 22753 9673 22787 9707
rect 24777 9673 24811 9707
rect 26065 9673 26099 9707
rect 1758 9605 1792 9639
rect 1869 9605 1903 9639
rect 2237 9605 2271 9639
rect 2973 9605 3007 9639
rect 10793 9605 10827 9639
rect 14933 9605 14967 9639
rect 18245 9605 18279 9639
rect 1961 9537 1995 9571
rect 2605 9537 2639 9571
rect 5273 9537 5307 9571
rect 11161 9537 11195 9571
rect 13369 9537 13403 9571
rect 19257 9537 19291 9571
rect 21833 9537 21867 9571
rect 23765 9537 23799 9571
rect 24225 9537 24259 9571
rect 1593 9469 1627 9503
rect 3157 9469 3191 9503
rect 3617 9469 3651 9503
rect 4813 9469 4847 9503
rect 4905 9469 4939 9503
rect 5089 9469 5123 9503
rect 6009 9469 6043 9503
rect 7113 9469 7147 9503
rect 7481 9469 7515 9503
rect 15025 9469 15059 9503
rect 15485 9469 15519 9503
rect 18061 9469 18095 9503
rect 18521 9469 18555 9503
rect 20796 9469 20830 9503
rect 25272 9469 25306 9503
rect 25697 9469 25731 9503
rect 4629 9401 4663 9435
rect 8677 9401 8711 9435
rect 8769 9401 8803 9435
rect 9321 9401 9355 9435
rect 10241 9401 10275 9435
rect 10333 9401 10367 9435
rect 13093 9401 13127 9435
rect 13185 9401 13219 9435
rect 16129 9401 16163 9435
rect 16221 9401 16255 9435
rect 16773 9401 16807 9435
rect 19349 9401 19383 9435
rect 19901 9401 19935 9435
rect 21281 9401 21315 9435
rect 22195 9401 22229 9435
rect 23029 9401 23063 9435
rect 23397 9401 23431 9435
rect 23857 9401 23891 9435
rect 25053 9401 25087 9435
rect 3249 9333 3283 9367
rect 4353 9333 4387 9367
rect 7021 9333 7055 9367
rect 14105 9333 14139 9367
rect 15209 9333 15243 9367
rect 15853 9333 15887 9367
rect 17693 9333 17727 9367
rect 18889 9333 18923 9367
rect 20867 9333 20901 9367
rect 21557 9333 21591 9367
rect 25375 9333 25409 9367
rect 1961 9129 1995 9163
rect 5825 9129 5859 9163
rect 10701 9129 10735 9163
rect 22569 9129 22603 9163
rect 2329 9061 2363 9095
rect 3157 9061 3191 9095
rect 3893 9061 3927 9095
rect 4077 9061 4111 9095
rect 7935 9061 7969 9095
rect 9873 9061 9907 9095
rect 12443 9061 12477 9095
rect 13737 9061 13771 9095
rect 15577 9061 15611 9095
rect 17141 9061 17175 9095
rect 17693 9061 17727 9095
rect 18975 9061 19009 9095
rect 22011 9061 22045 9095
rect 22937 9061 22971 9095
rect 24409 9061 24443 9095
rect 25099 9061 25133 9095
rect 1409 8993 1443 9027
rect 2881 8993 2915 9027
rect 4353 8993 4387 9027
rect 5089 8993 5123 9027
rect 6101 8993 6135 9027
rect 6561 8993 6595 9027
rect 14264 8993 14298 9027
rect 18613 8993 18647 9027
rect 23673 8993 23707 9027
rect 23857 8993 23891 9027
rect 25007 8993 25041 9027
rect 6745 8925 6779 8959
rect 7573 8925 7607 8959
rect 9781 8925 9815 8959
rect 10057 8925 10091 8959
rect 12081 8925 12115 8959
rect 15485 8925 15519 8959
rect 16129 8925 16163 8959
rect 17049 8925 17083 8959
rect 21649 8925 21683 8959
rect 23949 8925 23983 8959
rect 1593 8857 1627 8891
rect 8493 8857 8527 8891
rect 9229 8857 9263 8891
rect 13001 8857 13035 8891
rect 13369 8857 13403 8891
rect 14335 8857 14369 8891
rect 15025 8857 15059 8891
rect 21557 8857 21591 8891
rect 3525 8789 3559 8823
rect 5457 8789 5491 8823
rect 7113 8789 7147 8823
rect 7481 8789 7515 8823
rect 8769 8789 8803 8823
rect 16405 8789 16439 8823
rect 19533 8789 19567 8823
rect 19809 8789 19843 8823
rect 21189 8789 21223 8823
rect 23213 8789 23247 8823
rect 4813 8585 4847 8619
rect 6101 8585 6135 8619
rect 6469 8585 6503 8619
rect 7021 8585 7055 8619
rect 8493 8585 8527 8619
rect 8769 8585 8803 8619
rect 9137 8585 9171 8619
rect 11805 8585 11839 8619
rect 13369 8585 13403 8619
rect 14289 8585 14323 8619
rect 14611 8585 14645 8619
rect 17049 8585 17083 8619
rect 17877 8585 17911 8619
rect 18291 8585 18325 8619
rect 20269 8585 20303 8619
rect 20867 8585 20901 8619
rect 23029 8585 23063 8619
rect 25375 8585 25409 8619
rect 11483 8517 11517 8551
rect 18061 8517 18095 8551
rect 18613 8517 18647 8551
rect 19809 8517 19843 8551
rect 23489 8517 23523 8551
rect 2697 8449 2731 8483
rect 5549 8449 5583 8483
rect 7573 8449 7607 8483
rect 9689 8449 9723 8483
rect 15485 8449 15519 8483
rect 18981 8449 19015 8483
rect 19257 8449 19291 8483
rect 21833 8449 21867 8483
rect 23765 8449 23799 8483
rect 24225 8449 24259 8483
rect 1777 8381 1811 8415
rect 3157 8381 3191 8415
rect 4997 8381 5031 8415
rect 5457 8381 5491 8415
rect 11412 8381 11446 8415
rect 12449 8381 12483 8415
rect 14508 8381 14542 8415
rect 14933 8381 14967 8415
rect 15393 8381 15427 8415
rect 18061 8381 18095 8415
rect 18188 8381 18222 8415
rect 20764 8381 20798 8415
rect 21281 8381 21315 8415
rect 22753 8381 22787 8415
rect 25272 8381 25306 8415
rect 25697 8381 25731 8415
rect 1593 8313 1627 8347
rect 3478 8313 3512 8347
rect 7481 8313 7515 8347
rect 7935 8313 7969 8347
rect 9413 8313 9447 8347
rect 9505 8313 9539 8347
rect 10701 8313 10735 8347
rect 11253 8313 11287 8347
rect 12770 8313 12804 8347
rect 13645 8313 13679 8347
rect 15847 8313 15881 8347
rect 17325 8313 17359 8347
rect 19349 8313 19383 8347
rect 22154 8313 22188 8347
rect 23857 8313 23891 8347
rect 3065 8245 3099 8279
rect 4077 8245 4111 8279
rect 4353 8245 4387 8279
rect 10333 8245 10367 8279
rect 12173 8245 12207 8279
rect 16405 8245 16439 8279
rect 21741 8245 21775 8279
rect 25053 8245 25087 8279
rect 2053 8041 2087 8075
rect 3249 8041 3283 8075
rect 5181 8041 5215 8075
rect 5825 8041 5859 8075
rect 7665 8041 7699 8075
rect 12357 8041 12391 8075
rect 13001 8041 13035 8075
rect 15117 8041 15151 8075
rect 16129 8041 16163 8075
rect 17509 8041 17543 8075
rect 18429 8041 18463 8075
rect 19349 8041 19383 8075
rect 22753 8041 22787 8075
rect 23489 8041 23523 8075
rect 2329 7973 2363 8007
rect 4261 7973 4295 8007
rect 6653 7973 6687 8007
rect 8769 7973 8803 8007
rect 10051 7973 10085 8007
rect 11758 7973 11792 8007
rect 13553 7973 13587 8007
rect 13737 7973 13771 8007
rect 13829 7973 13863 8007
rect 15715 7973 15749 8007
rect 16910 7973 16944 8007
rect 22154 7973 22188 8007
rect 23765 7973 23799 8007
rect 8033 7905 8067 7939
rect 8585 7905 8619 7939
rect 15612 7905 15646 7939
rect 16589 7905 16623 7939
rect 18337 7905 18371 7939
rect 18797 7905 18831 7939
rect 25196 7905 25230 7939
rect 2237 7837 2271 7871
rect 2605 7837 2639 7871
rect 4169 7837 4203 7871
rect 4445 7837 4479 7871
rect 6377 7837 6411 7871
rect 6561 7837 6595 7871
rect 9689 7837 9723 7871
rect 11437 7837 11471 7871
rect 14013 7837 14047 7871
rect 21833 7837 21867 7871
rect 23673 7837 23707 7871
rect 25283 7837 25317 7871
rect 7113 7769 7147 7803
rect 21373 7769 21407 7803
rect 24225 7769 24259 7803
rect 1685 7701 1719 7735
rect 3617 7701 3651 7735
rect 5457 7701 5491 7735
rect 9413 7701 9447 7735
rect 10609 7701 10643 7735
rect 12633 7701 12667 7735
rect 21649 7701 21683 7735
rect 1731 7497 1765 7531
rect 2237 7497 2271 7531
rect 3985 7497 4019 7531
rect 4353 7497 4387 7531
rect 5917 7497 5951 7531
rect 6285 7497 6319 7531
rect 8539 7497 8573 7531
rect 8861 7497 8895 7531
rect 11345 7497 11379 7531
rect 13461 7497 13495 7531
rect 16221 7497 16255 7531
rect 17095 7497 17129 7531
rect 18337 7497 18371 7531
rect 22845 7497 22879 7531
rect 25053 7497 25087 7531
rect 25375 7497 25409 7531
rect 25789 7497 25823 7531
rect 3709 7429 3743 7463
rect 10149 7429 10183 7463
rect 17785 7429 17819 7463
rect 19257 7429 19291 7463
rect 4997 7361 5031 7395
rect 8033 7361 8067 7395
rect 10885 7361 10919 7395
rect 13737 7361 13771 7395
rect 14013 7361 14047 7395
rect 18705 7361 18739 7395
rect 19625 7361 19659 7395
rect 21649 7361 21683 7395
rect 1660 7293 1694 7327
rect 2789 7293 2823 7327
rect 6653 7293 6687 7327
rect 7113 7293 7147 7327
rect 7297 7293 7331 7327
rect 8468 7293 8502 7327
rect 11161 7293 11195 7327
rect 11989 7293 12023 7327
rect 12516 7293 12550 7327
rect 15209 7293 15243 7327
rect 15761 7293 15795 7327
rect 16992 7293 17026 7327
rect 17417 7293 17451 7327
rect 20177 7293 20211 7327
rect 20637 7293 20671 7327
rect 21741 7293 21775 7327
rect 22293 7293 22327 7327
rect 23673 7293 23707 7327
rect 24133 7293 24167 7327
rect 24685 7293 24719 7327
rect 25272 7293 25306 7327
rect 26065 7293 26099 7327
rect 2697 7225 2731 7259
rect 3151 7225 3185 7259
rect 4905 7225 4939 7259
rect 5359 7225 5393 7259
rect 9597 7225 9631 7259
rect 9689 7225 9723 7259
rect 13829 7225 13863 7259
rect 14749 7225 14783 7259
rect 18797 7225 18831 7259
rect 19993 7225 20027 7259
rect 6929 7157 6963 7191
rect 9413 7157 9447 7191
rect 10609 7157 10643 7191
rect 11713 7157 11747 7191
rect 12587 7157 12621 7191
rect 13001 7157 13035 7191
rect 15025 7157 15059 7191
rect 15485 7157 15519 7191
rect 16681 7157 16715 7191
rect 20269 7157 20303 7191
rect 21189 7157 21223 7191
rect 21833 7157 21867 7191
rect 23397 7157 23431 7191
rect 23765 7157 23799 7191
rect 1869 6953 1903 6987
rect 5549 6953 5583 6987
rect 9781 6953 9815 6987
rect 13737 6953 13771 6987
rect 17417 6953 17451 6987
rect 18797 6953 18831 6987
rect 19073 6953 19107 6987
rect 19763 6953 19797 6987
rect 20269 6953 20303 6987
rect 24317 6953 24351 6987
rect 25145 6953 25179 6987
rect 4905 6885 4939 6919
rect 6095 6885 6129 6919
rect 7665 6885 7699 6919
rect 12725 6885 12759 6919
rect 18198 6885 18232 6919
rect 21878 6885 21912 6919
rect 23489 6885 23523 6919
rect 1476 6817 1510 6851
rect 2421 6817 2455 6851
rect 2568 6817 2602 6851
rect 3525 6817 3559 6851
rect 4445 6817 4479 6851
rect 4721 6817 4755 6851
rect 5733 6817 5767 6851
rect 9689 6817 9723 6851
rect 10149 6817 10183 6851
rect 10701 6817 10735 6851
rect 11304 6817 11338 6851
rect 14264 6817 14298 6851
rect 15336 6817 15370 6851
rect 15439 6817 15473 6851
rect 16497 6817 16531 6851
rect 16773 6817 16807 6851
rect 19660 6817 19694 6851
rect 24041 6817 24075 6851
rect 24685 6817 24719 6851
rect 24869 6817 24903 6851
rect 25421 6817 25455 6851
rect 2789 6749 2823 6783
rect 2973 6749 3007 6783
rect 6929 6749 6963 6783
rect 7573 6749 7607 6783
rect 8033 6749 8067 6783
rect 8861 6749 8895 6783
rect 9505 6749 9539 6783
rect 11391 6749 11425 6783
rect 12633 6749 12667 6783
rect 17049 6749 17083 6783
rect 17877 6749 17911 6783
rect 21557 6749 21591 6783
rect 23397 6749 23431 6783
rect 3801 6681 3835 6715
rect 6653 6681 6687 6715
rect 13185 6681 13219 6715
rect 22477 6681 22511 6715
rect 23121 6681 23155 6715
rect 1547 6613 1581 6647
rect 2329 6613 2363 6647
rect 2697 6613 2731 6647
rect 5181 6613 5215 6647
rect 7297 6613 7331 6647
rect 8585 6613 8619 6647
rect 11713 6613 11747 6647
rect 14105 6613 14139 6647
rect 14335 6613 14369 6647
rect 15761 6613 15795 6647
rect 16221 6613 16255 6647
rect 17785 6613 17819 6647
rect 21465 6613 21499 6647
rect 22845 6613 22879 6647
rect 2789 6409 2823 6443
rect 3065 6409 3099 6443
rect 4721 6409 4755 6443
rect 6193 6409 6227 6443
rect 7389 6409 7423 6443
rect 8493 6409 8527 6443
rect 9045 6409 9079 6443
rect 9413 6409 9447 6443
rect 11621 6409 11655 6443
rect 12265 6409 12299 6443
rect 14749 6409 14783 6443
rect 15209 6409 15243 6443
rect 16405 6409 16439 6443
rect 17003 6409 17037 6443
rect 19625 6409 19659 6443
rect 23029 6409 23063 6443
rect 13277 6341 13311 6375
rect 23489 6341 23523 6375
rect 2421 6273 2455 6307
rect 3801 6273 3835 6307
rect 4905 6273 4939 6307
rect 5549 6273 5583 6307
rect 7573 6273 7607 6307
rect 8033 6273 8067 6307
rect 11253 6273 11287 6307
rect 13829 6273 13863 6307
rect 14197 6273 14231 6307
rect 15393 6273 15427 6307
rect 16773 6273 16807 6307
rect 2329 6205 2363 6239
rect 3525 6205 3559 6239
rect 3709 6205 3743 6239
rect 4353 6205 4387 6239
rect 9505 6205 9539 6239
rect 9965 6205 9999 6239
rect 10517 6205 10551 6239
rect 10977 6205 11011 6239
rect 12776 6205 12810 6239
rect 16932 6205 16966 6239
rect 18153 6205 18187 6239
rect 20177 6205 20211 6239
rect 20453 6205 20487 6239
rect 21557 6205 21591 6239
rect 23673 6205 23707 6239
rect 24133 6205 24167 6239
rect 25237 6205 25271 6239
rect 25789 6205 25823 6239
rect 4997 6137 5031 6171
rect 6653 6137 6687 6171
rect 7665 6137 7699 6171
rect 13921 6137 13955 6171
rect 15485 6137 15519 6171
rect 16037 6137 16071 6171
rect 18474 6137 18508 6171
rect 21878 6137 21912 6171
rect 5917 6069 5951 6103
rect 9689 6069 9723 6103
rect 10333 6069 10367 6103
rect 12863 6069 12897 6103
rect 13645 6069 13679 6103
rect 17417 6069 17451 6103
rect 17877 6069 17911 6103
rect 19073 6069 19107 6103
rect 19993 6069 20027 6103
rect 21097 6069 21131 6103
rect 21373 6069 21407 6103
rect 22477 6069 22511 6103
rect 23765 6069 23799 6103
rect 24869 6069 24903 6103
rect 25421 6069 25455 6103
rect 1547 5865 1581 5899
rect 1961 5865 1995 5899
rect 5273 5865 5307 5899
rect 6285 5865 6319 5899
rect 6929 5865 6963 5899
rect 7941 5865 7975 5899
rect 10977 5865 11011 5899
rect 13461 5865 13495 5899
rect 16221 5865 16255 5899
rect 18429 5865 18463 5899
rect 19993 5865 20027 5899
rect 21005 5865 21039 5899
rect 24225 5865 24259 5899
rect 25237 5865 25271 5899
rect 3157 5797 3191 5831
rect 4715 5797 4749 5831
rect 7383 5797 7417 5831
rect 8217 5797 8251 5831
rect 13093 5797 13127 5831
rect 13737 5797 13771 5831
rect 13829 5797 13863 5831
rect 15622 5797 15656 5831
rect 17233 5797 17267 5831
rect 18981 5797 19015 5831
rect 19073 5797 19107 5831
rect 20361 5797 20395 5831
rect 22753 5797 22787 5831
rect 23305 5797 23339 5831
rect 1444 5729 1478 5763
rect 2421 5729 2455 5763
rect 10057 5729 10091 5763
rect 10333 5729 10367 5763
rect 12081 5729 12115 5763
rect 12633 5729 12667 5763
rect 14749 5729 14783 5763
rect 20913 5729 20947 5763
rect 21373 5729 21407 5763
rect 24133 5729 24167 5763
rect 24593 5729 24627 5763
rect 2789 5661 2823 5695
rect 3801 5661 3835 5695
rect 4353 5661 4387 5695
rect 5549 5661 5583 5695
rect 5917 5661 5951 5695
rect 7021 5661 7055 5695
rect 2559 5593 2593 5627
rect 10701 5661 10735 5695
rect 12817 5661 12851 5695
rect 15301 5661 15335 5695
rect 17141 5661 17175 5695
rect 22661 5661 22695 5695
rect 10609 5593 10643 5627
rect 14289 5593 14323 5627
rect 17693 5593 17727 5627
rect 19533 5593 19567 5627
rect 2237 5525 2271 5559
rect 2697 5525 2731 5559
rect 3433 5525 3467 5559
rect 10057 5525 10091 5559
rect 10149 5525 10183 5559
rect 10471 5525 10505 5559
rect 11345 5525 11379 5559
rect 18061 5525 18095 5559
rect 21925 5525 21959 5559
rect 22385 5525 22419 5559
rect 23765 5525 23799 5559
rect 1850 5321 1884 5355
rect 2329 5321 2363 5355
rect 4445 5321 4479 5355
rect 6285 5321 6319 5355
rect 8401 5321 8435 5355
rect 10793 5321 10827 5355
rect 11161 5321 11195 5355
rect 12081 5321 12115 5355
rect 12725 5321 12759 5355
rect 13093 5321 13127 5355
rect 14841 5321 14875 5355
rect 17233 5321 17267 5355
rect 19625 5321 19659 5355
rect 20729 5321 20763 5355
rect 22753 5321 22787 5355
rect 23397 5321 23431 5355
rect 24685 5321 24719 5355
rect 1961 5253 1995 5287
rect 3065 5253 3099 5287
rect 10655 5253 10689 5287
rect 19349 5253 19383 5287
rect 2053 5185 2087 5219
rect 2881 5185 2915 5219
rect 3985 5185 4019 5219
rect 4905 5185 4939 5219
rect 6837 5185 6871 5219
rect 10241 5185 10275 5219
rect 10885 5185 10919 5219
rect 13921 5185 13955 5219
rect 15669 5185 15703 5219
rect 16865 5185 16899 5219
rect 21189 5185 21223 5219
rect 3525 5117 3559 5151
rect 3801 5117 3835 5151
rect 6653 5117 6687 5151
rect 8585 5117 8619 5151
rect 9045 5117 9079 5151
rect 1685 5049 1719 5083
rect 2789 5049 2823 5083
rect 2881 5049 2915 5083
rect 4997 5049 5031 5083
rect 5549 5049 5583 5083
rect 7199 5049 7233 5083
rect 8033 5049 8067 5083
rect 12909 5117 12943 5151
rect 13369 5117 13403 5151
rect 18981 5117 19015 5151
rect 20085 5117 20119 5151
rect 23673 5117 23707 5151
rect 24225 5117 24259 5151
rect 25237 5117 25271 5151
rect 25789 5117 25823 5151
rect 10517 5049 10551 5083
rect 14283 5049 14317 5083
rect 15990 5049 16024 5083
rect 18337 5049 18371 5083
rect 18438 5049 18472 5083
rect 21510 5049 21544 5083
rect 22385 5049 22419 5083
rect 5825 4981 5859 5015
rect 7757 4981 7791 5015
rect 8677 4981 8711 5015
rect 9689 4981 9723 5015
rect 9965 4981 9999 5015
rect 10241 4981 10275 5015
rect 10333 4981 10367 5015
rect 11529 4981 11563 5015
rect 13829 4981 13863 5015
rect 15301 4981 15335 5015
rect 16589 4981 16623 5015
rect 17785 4981 17819 5015
rect 20269 4981 20303 5015
rect 21097 4981 21131 5015
rect 22109 4981 22143 5015
rect 23765 4981 23799 5015
rect 25421 4981 25455 5015
rect 1547 4777 1581 4811
rect 2329 4777 2363 4811
rect 3433 4777 3467 4811
rect 3893 4777 3927 4811
rect 4261 4777 4295 4811
rect 4721 4777 4755 4811
rect 6929 4777 6963 4811
rect 8217 4777 8251 4811
rect 8585 4777 8619 4811
rect 9045 4777 9079 4811
rect 10793 4777 10827 4811
rect 11069 4777 11103 4811
rect 11345 4777 11379 4811
rect 14473 4777 14507 4811
rect 15025 4777 15059 4811
rect 17509 4777 17543 4811
rect 18153 4777 18187 4811
rect 19349 4777 19383 4811
rect 22569 4777 22603 4811
rect 1961 4709 1995 4743
rect 3157 4709 3191 4743
rect 5089 4709 5123 4743
rect 5641 4709 5675 4743
rect 7297 4709 7331 4743
rect 7389 4709 7423 4743
rect 9689 4709 9723 4743
rect 10425 4709 10459 4743
rect 13645 4709 13679 4743
rect 14197 4709 14231 4743
rect 16221 4709 16255 4743
rect 16773 4709 16807 4743
rect 18429 4709 18463 4743
rect 21418 4709 21452 4743
rect 23029 4709 23063 4743
rect 23581 4709 23615 4743
rect 1476 4641 1510 4675
rect 2421 4641 2455 4675
rect 6561 4641 6595 4675
rect 9413 4641 9447 4675
rect 11529 4641 11563 4675
rect 11805 4641 11839 4675
rect 19876 4641 19910 4675
rect 24685 4641 24719 4675
rect 24869 4641 24903 4675
rect 2789 4573 2823 4607
rect 4997 4573 5031 4607
rect 5917 4573 5951 4607
rect 7573 4573 7607 4607
rect 10057 4573 10091 4607
rect 13553 4573 13587 4607
rect 16129 4573 16163 4607
rect 18337 4573 18371 4607
rect 18981 4573 19015 4607
rect 21097 4573 21131 4607
rect 22937 4573 22971 4607
rect 24961 4573 24995 4607
rect 2697 4505 2731 4539
rect 9854 4505 9888 4539
rect 20729 4505 20763 4539
rect 2586 4437 2620 4471
rect 9965 4437 9999 4471
rect 12265 4437 12299 4471
rect 13277 4437 13311 4471
rect 15669 4437 15703 4471
rect 17049 4437 17083 4471
rect 19947 4437 19981 4471
rect 22017 4437 22051 4471
rect 24225 4437 24259 4471
rect 1961 4233 1995 4267
rect 2881 4233 2915 4267
rect 3341 4233 3375 4267
rect 7665 4233 7699 4267
rect 7849 4233 7883 4267
rect 9689 4233 9723 4267
rect 10057 4233 10091 4267
rect 10793 4233 10827 4267
rect 11253 4233 11287 4267
rect 12173 4233 12207 4267
rect 16129 4233 16163 4267
rect 17509 4233 17543 4267
rect 18981 4233 19015 4267
rect 19717 4233 19751 4267
rect 21833 4233 21867 4267
rect 24777 4233 24811 4267
rect 6009 4097 6043 4131
rect 6929 4097 6963 4131
rect 7297 4097 7331 4131
rect 1869 4029 1903 4063
rect 2605 4029 2639 4063
rect 3433 4029 3467 4063
rect 3985 4029 4019 4063
rect 1777 3961 1811 3995
rect 4169 3961 4203 3995
rect 5089 3961 5123 3995
rect 5181 3961 5215 3995
rect 5733 3961 5767 3995
rect 7021 3961 7055 3995
rect 9919 4165 9953 4199
rect 15761 4165 15795 4199
rect 8309 4097 8343 4131
rect 8953 4097 8987 4131
rect 10149 4097 10183 4131
rect 13001 4097 13035 4131
rect 14013 4097 14047 4131
rect 14657 4097 14691 4131
rect 16497 4097 16531 4131
rect 17141 4097 17175 4131
rect 19901 4097 19935 4131
rect 22661 4097 22695 4131
rect 25789 4097 25823 4131
rect 8401 4029 8435 4063
rect 8585 4029 8619 4063
rect 9229 4029 9263 4063
rect 9781 4029 9815 4063
rect 11345 4029 11379 4063
rect 11805 4029 11839 4063
rect 12449 4029 12483 4063
rect 18061 4029 18095 4063
rect 23029 4029 23063 4063
rect 23489 4029 23523 4063
rect 23673 4029 23707 4063
rect 24133 4029 24167 4063
rect 25053 4029 25087 4063
rect 25237 4029 25271 4063
rect 14105 3961 14139 3995
rect 15393 3961 15427 3995
rect 16589 3961 16623 3995
rect 18382 3961 18416 3995
rect 19993 3961 20027 3995
rect 20545 3961 20579 3995
rect 22017 3961 22051 3995
rect 22109 3961 22143 3995
rect 4445 3893 4479 3927
rect 4905 3893 4939 3927
rect 6653 3893 6687 3927
rect 7665 3893 7699 3927
rect 10425 3893 10459 3927
rect 11529 3893 11563 3927
rect 12633 3893 12667 3927
rect 13553 3893 13587 3927
rect 14933 3893 14967 3927
rect 17877 3893 17911 3927
rect 19257 3893 19291 3927
rect 21097 3893 21131 3927
rect 23765 3893 23799 3927
rect 25421 3893 25455 3927
rect 2237 3689 2271 3723
rect 2881 3689 2915 3723
rect 3433 3689 3467 3723
rect 3801 3689 3835 3723
rect 4261 3689 4295 3723
rect 5365 3689 5399 3723
rect 5641 3689 5675 3723
rect 6377 3689 6411 3723
rect 8217 3689 8251 3723
rect 9413 3689 9447 3723
rect 9873 3689 9907 3723
rect 10241 3689 10275 3723
rect 12449 3689 12483 3723
rect 14657 3689 14691 3723
rect 16497 3689 16531 3723
rect 19993 3689 20027 3723
rect 20269 3689 20303 3723
rect 21189 3689 21223 3723
rect 22661 3689 22695 3723
rect 23489 3689 23523 3723
rect 24869 3689 24903 3723
rect 4807 3621 4841 3655
rect 7389 3621 7423 3655
rect 8677 3621 8711 3655
rect 10609 3621 10643 3655
rect 11621 3621 11655 3655
rect 12173 3621 12207 3655
rect 13829 3621 13863 3655
rect 14381 3621 14415 3655
rect 15485 3621 15519 3655
rect 16037 3621 16071 3655
rect 16865 3621 16899 3655
rect 18429 3621 18463 3655
rect 18981 3621 19015 3655
rect 21465 3621 21499 3655
rect 21833 3621 21867 3655
rect 23029 3621 23063 3655
rect 1476 3553 1510 3587
rect 2881 3553 2915 3587
rect 4445 3553 4479 3587
rect 6009 3553 6043 3587
rect 6193 3553 6227 3587
rect 10756 3553 10790 3587
rect 12357 3553 12391 3587
rect 17141 3553 17175 3587
rect 19809 3553 19843 3587
rect 23213 3553 23247 3587
rect 23673 3553 23707 3587
rect 25053 3553 25087 3587
rect 25237 3553 25271 3587
rect 7113 3485 7147 3519
rect 7297 3485 7331 3519
rect 7573 3485 7607 3519
rect 10977 3485 11011 3519
rect 13001 3485 13035 3519
rect 13737 3485 13771 3519
rect 15117 3485 15151 3519
rect 15393 3485 15427 3519
rect 17785 3485 17819 3519
rect 18337 3485 18371 3519
rect 19349 3485 19383 3519
rect 21741 3485 21775 3519
rect 22385 3485 22419 3519
rect 24593 3485 24627 3519
rect 11989 3417 12023 3451
rect 1547 3349 1581 3383
rect 1961 3349 1995 3383
rect 7021 3349 7055 3383
rect 7113 3349 7147 3383
rect 9045 3349 9079 3383
rect 10885 3349 10919 3383
rect 11253 3349 11287 3383
rect 13369 3349 13403 3383
rect 17325 3349 17359 3383
rect 18153 3349 18187 3383
rect 24225 3349 24259 3383
rect 1593 3145 1627 3179
rect 2881 3145 2915 3179
rect 6193 3145 6227 3179
rect 6653 3145 6687 3179
rect 7849 3145 7883 3179
rect 8125 3145 8159 3179
rect 9781 3145 9815 3179
rect 10057 3145 10091 3179
rect 10406 3145 10440 3179
rect 11253 3145 11287 3179
rect 12173 3145 12207 3179
rect 13737 3145 13771 3179
rect 14013 3145 14047 3179
rect 15485 3145 15519 3179
rect 15761 3145 15795 3179
rect 16037 3145 16071 3179
rect 16129 3145 16163 3179
rect 17325 3145 17359 3179
rect 19901 3145 19935 3179
rect 22707 3145 22741 3179
rect 23121 3145 23155 3179
rect 23489 3145 23523 3179
rect 23811 3145 23845 3179
rect 24685 3145 24719 3179
rect 25053 3145 25087 3179
rect 25789 3145 25823 3179
rect 5549 3077 5583 3111
rect 10517 3077 10551 3111
rect 10701 3077 10735 3111
rect 3157 3009 3191 3043
rect 4537 3009 4571 3043
rect 8585 3009 8619 3043
rect 10609 3009 10643 3043
rect 12817 3009 12851 3043
rect 1961 2941 1995 2975
rect 3433 2941 3467 2975
rect 3801 2941 3835 2975
rect 6929 2941 6963 2975
rect 8953 2941 8987 2975
rect 9229 2941 9263 2975
rect 10241 2941 10275 2975
rect 11713 2941 11747 2975
rect 14565 2941 14599 2975
rect 2513 2873 2547 2907
rect 4077 2873 4111 2907
rect 4997 2873 5031 2907
rect 5089 2873 5123 2907
rect 7250 2873 7284 2907
rect 13138 2873 13172 2907
rect 14381 2873 14415 2907
rect 14886 2873 14920 2907
rect 23949 3077 23983 3111
rect 16405 3009 16439 3043
rect 17049 3009 17083 3043
rect 18797 3009 18831 3043
rect 19073 3009 19107 3043
rect 20361 3009 20395 3043
rect 20821 3009 20855 3043
rect 22477 3009 22511 3043
rect 24041 3009 24075 3043
rect 22636 2941 22670 2975
rect 23673 2941 23707 2975
rect 25237 2941 25271 2975
rect 26157 2941 26191 2975
rect 16497 2873 16531 2907
rect 18337 2873 18371 2907
rect 18889 2873 18923 2907
rect 20729 2873 20763 2907
rect 21142 2873 21176 2907
rect 8769 2805 8803 2839
rect 12633 2805 12667 2839
rect 16037 2805 16071 2839
rect 17785 2805 17819 2839
rect 21741 2805 21775 2839
rect 22017 2805 22051 2839
rect 24317 2805 24351 2839
rect 25421 2805 25455 2839
rect 3801 2601 3835 2635
rect 4997 2601 5031 2635
rect 6009 2601 6043 2635
rect 6653 2601 6687 2635
rect 7941 2601 7975 2635
rect 9137 2601 9171 2635
rect 13645 2601 13679 2635
rect 14565 2601 14599 2635
rect 15669 2601 15703 2635
rect 16313 2601 16347 2635
rect 17417 2601 17451 2635
rect 19257 2601 19291 2635
rect 20223 2601 20257 2635
rect 22293 2601 22327 2635
rect 22753 2601 22787 2635
rect 23765 2601 23799 2635
rect 24133 2601 24167 2635
rect 25421 2601 25455 2635
rect 4537 2533 4571 2567
rect 5451 2533 5485 2567
rect 7113 2533 7147 2567
rect 7665 2533 7699 2567
rect 8309 2533 8343 2567
rect 11713 2533 11747 2567
rect 13046 2533 13080 2567
rect 16818 2533 16852 2567
rect 18061 2533 18095 2567
rect 18658 2533 18692 2567
rect 21005 2533 21039 2567
rect 21465 2533 21499 2567
rect 23489 2533 23523 2567
rect 1476 2465 1510 2499
rect 1869 2465 1903 2499
rect 2329 2465 2363 2499
rect 2697 2465 2731 2499
rect 2973 2465 3007 2499
rect 3433 2465 3467 2499
rect 4144 2465 4178 2499
rect 8677 2465 8711 2499
rect 9781 2465 9815 2499
rect 11161 2465 11195 2499
rect 11437 2465 11471 2499
rect 15485 2465 15519 2499
rect 15945 2465 15979 2499
rect 20152 2465 20186 2499
rect 20545 2465 20579 2499
rect 22845 2465 22879 2499
rect 24041 2465 24075 2499
rect 24593 2465 24627 2499
rect 25672 2465 25706 2499
rect 3157 2397 3191 2431
rect 5089 2397 5123 2431
rect 6285 2397 6319 2431
rect 7021 2397 7055 2431
rect 9505 2397 9539 2431
rect 10333 2397 10367 2431
rect 10701 2397 10735 2431
rect 11989 2397 12023 2431
rect 12725 2397 12759 2431
rect 13921 2397 13955 2431
rect 15301 2397 15335 2431
rect 16497 2397 16531 2431
rect 17785 2397 17819 2431
rect 18337 2397 18371 2431
rect 21373 2397 21407 2431
rect 21649 2397 21683 2431
rect 25053 2397 25087 2431
rect 1547 2261 1581 2295
rect 4215 2261 4249 2295
rect 8861 2261 8895 2295
rect 9965 2261 9999 2295
rect 12357 2261 12391 2295
rect 23029 2261 23063 2295
rect 25743 2261 25777 2295
rect 26157 2261 26191 2295
<< metal1 >>
rect 18322 26596 18328 26648
rect 18380 26636 18386 26648
rect 23474 26636 23480 26648
rect 18380 26608 23480 26636
rect 18380 26596 18386 26608
rect 23474 26596 23480 26608
rect 23532 26596 23538 26648
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 17126 24392 17132 24404
rect 17087 24364 17132 24392
rect 17126 24352 17132 24364
rect 17184 24352 17190 24404
rect 18230 24392 18236 24404
rect 18191 24364 18236 24392
rect 18230 24352 18236 24364
rect 18288 24352 18294 24404
rect 10686 24265 10692 24268
rect 10664 24259 10692 24265
rect 10664 24225 10676 24259
rect 10664 24219 10692 24225
rect 10686 24216 10692 24219
rect 10744 24216 10750 24268
rect 11606 24216 11612 24268
rect 11664 24265 11670 24268
rect 11664 24259 11702 24265
rect 11690 24225 11702 24259
rect 11664 24219 11702 24225
rect 16945 24259 17003 24265
rect 16945 24225 16957 24259
rect 16991 24256 17003 24259
rect 17310 24256 17316 24268
rect 16991 24228 17316 24256
rect 16991 24225 17003 24228
rect 16945 24219 17003 24225
rect 11664 24216 11670 24219
rect 17310 24216 17316 24228
rect 17368 24216 17374 24268
rect 18049 24259 18107 24265
rect 18049 24225 18061 24259
rect 18095 24256 18107 24259
rect 18690 24256 18696 24268
rect 18095 24228 18696 24256
rect 18095 24225 18107 24228
rect 18049 24219 18107 24225
rect 18690 24216 18696 24228
rect 18748 24216 18754 24268
rect 10042 24012 10048 24064
rect 10100 24052 10106 24064
rect 10735 24055 10793 24061
rect 10735 24052 10747 24055
rect 10100 24024 10747 24052
rect 10100 24012 10106 24024
rect 10735 24021 10747 24024
rect 10781 24021 10793 24055
rect 10735 24015 10793 24021
rect 11747 24055 11805 24061
rect 11747 24021 11759 24055
rect 11793 24052 11805 24055
rect 11882 24052 11888 24064
rect 11793 24024 11888 24052
rect 11793 24021 11805 24024
rect 11747 24015 11805 24021
rect 11882 24012 11888 24024
rect 11940 24012 11946 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 10686 23848 10692 23860
rect 10647 23820 10692 23848
rect 10686 23808 10692 23820
rect 10744 23808 10750 23860
rect 14550 23848 14556 23860
rect 14511 23820 14556 23848
rect 14550 23808 14556 23820
rect 14608 23808 14614 23860
rect 16206 23848 16212 23860
rect 16167 23820 16212 23848
rect 16206 23808 16212 23820
rect 16264 23808 16270 23860
rect 18230 23848 18236 23860
rect 18191 23820 18236 23848
rect 18230 23808 18236 23820
rect 18288 23808 18294 23860
rect 20346 23848 20352 23860
rect 20307 23820 20352 23848
rect 20346 23808 20352 23820
rect 20404 23808 20410 23860
rect 21450 23848 21456 23860
rect 21411 23820 21456 23848
rect 21450 23808 21456 23820
rect 21508 23808 21514 23860
rect 22554 23848 22560 23860
rect 22515 23820 22560 23848
rect 22554 23808 22560 23820
rect 22612 23808 22618 23860
rect 24762 23848 24768 23860
rect 24723 23820 24768 23848
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 8938 23644 8944 23656
rect 1443 23616 2084 23644
rect 8899 23616 8944 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 2056 23520 2084 23616
rect 8938 23604 8944 23616
rect 8996 23644 9002 23656
rect 11146 23653 11152 23656
rect 9401 23647 9459 23653
rect 9401 23644 9413 23647
rect 8996 23616 9413 23644
rect 8996 23604 9002 23616
rect 9401 23613 9413 23616
rect 9447 23613 9459 23647
rect 9401 23607 9459 23613
rect 11124 23647 11152 23653
rect 11124 23613 11136 23647
rect 11124 23607 11152 23613
rect 11146 23604 11152 23607
rect 11204 23604 11210 23656
rect 12434 23604 12440 23656
rect 12492 23653 12498 23656
rect 12492 23647 12530 23653
rect 12518 23644 12530 23647
rect 12897 23647 12955 23653
rect 12897 23644 12909 23647
rect 12518 23616 12909 23644
rect 12518 23613 12530 23616
rect 12492 23607 12530 23613
rect 12897 23613 12909 23616
rect 12943 23613 12955 23647
rect 12897 23607 12955 23613
rect 12492 23604 12498 23607
rect 13814 23604 13820 23656
rect 13872 23644 13878 23656
rect 14369 23647 14427 23653
rect 14369 23644 14381 23647
rect 13872 23616 14381 23644
rect 13872 23604 13878 23616
rect 14369 23613 14381 23616
rect 14415 23644 14427 23647
rect 14921 23647 14979 23653
rect 14921 23644 14933 23647
rect 14415 23616 14933 23644
rect 14415 23613 14427 23616
rect 14369 23607 14427 23613
rect 14921 23613 14933 23616
rect 14967 23613 14979 23647
rect 16022 23644 16028 23656
rect 15983 23616 16028 23644
rect 14921 23607 14979 23613
rect 16022 23604 16028 23616
rect 16080 23644 16086 23656
rect 16577 23647 16635 23653
rect 16577 23644 16589 23647
rect 16080 23616 16589 23644
rect 16080 23604 16086 23616
rect 16577 23613 16589 23616
rect 16623 23613 16635 23647
rect 16577 23607 16635 23613
rect 17865 23647 17923 23653
rect 17865 23613 17877 23647
rect 17911 23644 17923 23647
rect 18049 23647 18107 23653
rect 18049 23644 18061 23647
rect 17911 23616 18061 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 18049 23613 18061 23616
rect 18095 23644 18107 23647
rect 18138 23644 18144 23656
rect 18095 23616 18144 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 18138 23604 18144 23616
rect 18196 23604 18202 23656
rect 20165 23647 20223 23653
rect 20165 23613 20177 23647
rect 20211 23644 20223 23647
rect 21266 23644 21272 23656
rect 20211 23616 20852 23644
rect 21227 23616 21272 23644
rect 20211 23613 20223 23616
rect 20165 23607 20223 23613
rect 2038 23508 2044 23520
rect 1999 23480 2044 23508
rect 2038 23468 2044 23480
rect 2096 23468 2102 23520
rect 9122 23508 9128 23520
rect 9083 23480 9128 23508
rect 9122 23468 9128 23480
rect 9180 23468 9186 23520
rect 9950 23508 9956 23520
rect 9911 23480 9956 23508
rect 9950 23468 9956 23480
rect 10008 23468 10014 23520
rect 10962 23468 10968 23520
rect 11020 23508 11026 23520
rect 11195 23511 11253 23517
rect 11195 23508 11207 23511
rect 11020 23480 11207 23508
rect 11020 23468 11026 23480
rect 11195 23477 11207 23480
rect 11241 23477 11253 23511
rect 11606 23508 11612 23520
rect 11567 23480 11612 23508
rect 11195 23471 11253 23477
rect 11606 23468 11612 23480
rect 11664 23468 11670 23520
rect 12575 23511 12633 23517
rect 12575 23477 12587 23511
rect 12621 23508 12633 23511
rect 13354 23508 13360 23520
rect 12621 23480 13360 23508
rect 12621 23477 12633 23480
rect 12575 23471 12633 23477
rect 13354 23468 13360 23480
rect 13412 23468 13418 23520
rect 17037 23511 17095 23517
rect 17037 23477 17049 23511
rect 17083 23508 17095 23511
rect 17310 23508 17316 23520
rect 17083 23480 17316 23508
rect 17083 23477 17095 23480
rect 17037 23471 17095 23477
rect 17310 23468 17316 23480
rect 17368 23468 17374 23520
rect 18690 23508 18696 23520
rect 18651 23480 18696 23508
rect 18690 23468 18696 23480
rect 18748 23468 18754 23520
rect 20824 23517 20852 23616
rect 21266 23604 21272 23616
rect 21324 23644 21330 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 21324 23616 21833 23644
rect 21324 23604 21330 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 21821 23607 21879 23613
rect 22186 23604 22192 23656
rect 22244 23644 22250 23656
rect 22373 23647 22431 23653
rect 22373 23644 22385 23647
rect 22244 23616 22385 23644
rect 22244 23604 22250 23616
rect 22373 23613 22385 23616
rect 22419 23644 22431 23647
rect 22925 23647 22983 23653
rect 22925 23644 22937 23647
rect 22419 23616 22937 23644
rect 22419 23613 22431 23616
rect 22373 23607 22431 23613
rect 22925 23613 22937 23616
rect 22971 23613 22983 23647
rect 24578 23644 24584 23656
rect 24539 23616 24584 23644
rect 22925 23607 22983 23613
rect 24578 23604 24584 23616
rect 24636 23644 24642 23656
rect 25133 23647 25191 23653
rect 25133 23644 25145 23647
rect 24636 23616 25145 23644
rect 24636 23604 24642 23616
rect 25133 23613 25145 23616
rect 25179 23613 25191 23647
rect 25133 23607 25191 23613
rect 20809 23511 20867 23517
rect 20809 23477 20821 23511
rect 20855 23508 20867 23511
rect 21266 23508 21272 23520
rect 20855 23480 21272 23508
rect 20855 23477 20867 23480
rect 20809 23471 20867 23477
rect 21266 23468 21272 23480
rect 21324 23468 21330 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1394 23264 1400 23316
rect 1452 23304 1458 23316
rect 1581 23307 1639 23313
rect 1581 23304 1593 23307
rect 1452 23276 1593 23304
rect 1452 23264 1458 23276
rect 1581 23273 1593 23276
rect 1627 23273 1639 23307
rect 11146 23304 11152 23316
rect 11107 23276 11152 23304
rect 1581 23267 1639 23273
rect 11146 23264 11152 23276
rect 11204 23264 11210 23316
rect 13722 23313 13728 23316
rect 13679 23307 13728 23313
rect 13679 23273 13691 23307
rect 13725 23273 13728 23307
rect 13679 23267 13728 23273
rect 13722 23264 13728 23267
rect 13780 23264 13786 23316
rect 18233 23307 18291 23313
rect 18233 23273 18245 23307
rect 18279 23304 18291 23307
rect 18322 23304 18328 23316
rect 18279 23276 18328 23304
rect 18279 23273 18291 23276
rect 18233 23267 18291 23273
rect 18322 23264 18328 23276
rect 18380 23264 18386 23316
rect 24670 23264 24676 23316
rect 24728 23304 24734 23316
rect 24765 23307 24823 23313
rect 24765 23304 24777 23307
rect 24728 23276 24777 23304
rect 24728 23264 24734 23276
rect 24765 23273 24777 23276
rect 24811 23273 24823 23307
rect 24765 23267 24823 23273
rect 9858 23236 9864 23248
rect 9819 23208 9864 23236
rect 9858 23196 9864 23208
rect 9916 23196 9922 23248
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 1670 23168 1676 23180
rect 1443 23140 1676 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 1670 23128 1676 23140
rect 1728 23128 1734 23180
rect 7282 23128 7288 23180
rect 7340 23177 7346 23180
rect 7340 23171 7378 23177
rect 7366 23137 7378 23171
rect 7340 23131 7378 23137
rect 7340 23128 7346 23131
rect 8570 23128 8576 23180
rect 8628 23177 8634 23180
rect 11330 23177 11336 23180
rect 8628 23171 8666 23177
rect 8654 23137 8666 23171
rect 8628 23131 8666 23137
rect 11308 23171 11336 23177
rect 11308 23137 11320 23171
rect 11308 23131 11336 23137
rect 8628 23128 8634 23131
rect 11330 23128 11336 23131
rect 11388 23128 11394 23180
rect 12250 23128 12256 23180
rect 12308 23177 12314 23180
rect 12308 23171 12346 23177
rect 12334 23137 12346 23171
rect 12308 23131 12346 23137
rect 12308 23128 12314 23131
rect 13538 23128 13544 23180
rect 13596 23177 13602 23180
rect 15562 23177 15568 23180
rect 13596 23171 13634 23177
rect 13622 23137 13634 23171
rect 13596 23131 13634 23137
rect 15540 23171 15568 23177
rect 15540 23137 15552 23171
rect 15540 23131 15568 23137
rect 13596 23128 13602 23131
rect 15562 23128 15568 23131
rect 15620 23128 15626 23180
rect 16758 23128 16764 23180
rect 16816 23177 16822 23180
rect 16816 23171 16854 23177
rect 16842 23137 16854 23171
rect 18046 23168 18052 23180
rect 18007 23140 18052 23168
rect 16816 23131 16854 23137
rect 16816 23128 16822 23131
rect 18046 23128 18052 23140
rect 18104 23128 18110 23180
rect 24118 23128 24124 23180
rect 24176 23168 24182 23180
rect 24581 23171 24639 23177
rect 24581 23168 24593 23171
rect 24176 23140 24593 23168
rect 24176 23128 24182 23140
rect 24581 23137 24593 23140
rect 24627 23137 24639 23171
rect 24581 23131 24639 23137
rect 7466 23060 7472 23112
rect 7524 23100 7530 23112
rect 7745 23103 7803 23109
rect 7745 23100 7757 23103
rect 7524 23072 7757 23100
rect 7524 23060 7530 23072
rect 7745 23069 7757 23072
rect 7791 23069 7803 23103
rect 9766 23100 9772 23112
rect 9727 23072 9772 23100
rect 7745 23063 7803 23069
rect 9766 23060 9772 23072
rect 9824 23060 9830 23112
rect 10134 23100 10140 23112
rect 10095 23072 10140 23100
rect 10134 23060 10140 23072
rect 10192 23060 10198 23112
rect 7423 22967 7481 22973
rect 7423 22933 7435 22967
rect 7469 22964 7481 22967
rect 7650 22964 7656 22976
rect 7469 22936 7656 22964
rect 7469 22933 7481 22936
rect 7423 22927 7481 22933
rect 7650 22924 7656 22936
rect 7708 22924 7714 22976
rect 8754 22973 8760 22976
rect 8711 22967 8760 22973
rect 8711 22933 8723 22967
rect 8757 22933 8760 22967
rect 8711 22927 8760 22933
rect 8754 22924 8760 22927
rect 8812 22924 8818 22976
rect 11146 22924 11152 22976
rect 11204 22964 11210 22976
rect 11379 22967 11437 22973
rect 11379 22964 11391 22967
rect 11204 22936 11391 22964
rect 11204 22924 11210 22936
rect 11379 22933 11391 22936
rect 11425 22933 11437 22967
rect 11379 22927 11437 22933
rect 12342 22924 12348 22976
rect 12400 22973 12406 22976
rect 12400 22967 12449 22973
rect 12400 22933 12403 22967
rect 12437 22933 12449 22967
rect 12400 22927 12449 22933
rect 15611 22967 15669 22973
rect 15611 22933 15623 22967
rect 15657 22964 15669 22967
rect 15930 22964 15936 22976
rect 15657 22936 15936 22964
rect 15657 22933 15669 22936
rect 15611 22927 15669 22933
rect 12400 22924 12406 22927
rect 15930 22924 15936 22936
rect 15988 22924 15994 22976
rect 16899 22967 16957 22973
rect 16899 22933 16911 22967
rect 16945 22964 16957 22967
rect 17402 22964 17408 22976
rect 16945 22936 17408 22964
rect 16945 22933 16957 22936
rect 16899 22927 16957 22933
rect 17402 22924 17408 22936
rect 17460 22924 17466 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1486 22720 1492 22772
rect 1544 22760 1550 22772
rect 1581 22763 1639 22769
rect 1581 22760 1593 22763
rect 1544 22732 1593 22760
rect 1544 22720 1550 22732
rect 1581 22729 1593 22732
rect 1627 22729 1639 22763
rect 6270 22760 6276 22772
rect 6231 22732 6276 22760
rect 1581 22723 1639 22729
rect 6270 22720 6276 22732
rect 6328 22720 6334 22772
rect 8570 22760 8576 22772
rect 8531 22732 8576 22760
rect 8570 22720 8576 22732
rect 8628 22760 8634 22772
rect 9582 22760 9588 22772
rect 8628 22732 9588 22760
rect 8628 22720 8634 22732
rect 9582 22720 9588 22732
rect 9640 22720 9646 22772
rect 9766 22720 9772 22772
rect 9824 22760 9830 22772
rect 10597 22763 10655 22769
rect 10597 22760 10609 22763
rect 9824 22732 10609 22760
rect 9824 22720 9830 22732
rect 10597 22729 10609 22732
rect 10643 22729 10655 22763
rect 10597 22723 10655 22729
rect 13538 22720 13544 22772
rect 13596 22760 13602 22772
rect 14277 22763 14335 22769
rect 14277 22760 14289 22763
rect 13596 22732 14289 22760
rect 13596 22720 13602 22732
rect 14277 22729 14289 22732
rect 14323 22729 14335 22763
rect 15562 22760 15568 22772
rect 15523 22732 15568 22760
rect 14277 22723 14335 22729
rect 15562 22720 15568 22732
rect 15620 22720 15626 22772
rect 16758 22760 16764 22772
rect 16719 22732 16764 22760
rect 16758 22720 16764 22732
rect 16816 22720 16822 22772
rect 7193 22695 7251 22701
rect 7193 22661 7205 22695
rect 7239 22692 7251 22695
rect 7282 22692 7288 22704
rect 7239 22664 7288 22692
rect 7239 22661 7251 22664
rect 7193 22655 7251 22661
rect 7282 22652 7288 22664
rect 7340 22692 7346 22704
rect 7834 22692 7840 22704
rect 7340 22664 7840 22692
rect 7340 22652 7346 22664
rect 7834 22652 7840 22664
rect 7892 22652 7898 22704
rect 13814 22652 13820 22704
rect 13872 22692 13878 22704
rect 14599 22695 14657 22701
rect 14599 22692 14611 22695
rect 13872 22664 14611 22692
rect 13872 22652 13878 22664
rect 14599 22661 14611 22664
rect 14645 22661 14657 22695
rect 14599 22655 14657 22661
rect 17083 22695 17141 22701
rect 17083 22661 17095 22695
rect 17129 22692 17141 22695
rect 18046 22692 18052 22704
rect 17129 22664 18052 22692
rect 17129 22661 17141 22664
rect 17083 22655 17141 22661
rect 18046 22652 18052 22664
rect 18104 22692 18110 22704
rect 18233 22695 18291 22701
rect 18233 22692 18245 22695
rect 18104 22664 18245 22692
rect 18104 22652 18110 22664
rect 18233 22661 18245 22664
rect 18279 22661 18291 22695
rect 18233 22655 18291 22661
rect 7377 22627 7435 22633
rect 7377 22593 7389 22627
rect 7423 22624 7435 22627
rect 7466 22624 7472 22636
rect 7423 22596 7472 22624
rect 7423 22593 7435 22596
rect 7377 22587 7435 22593
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 7558 22584 7564 22636
rect 7616 22624 7622 22636
rect 7653 22627 7711 22633
rect 7653 22624 7665 22627
rect 7616 22596 7665 22624
rect 7616 22584 7622 22596
rect 7653 22593 7665 22596
rect 7699 22593 7711 22627
rect 7653 22587 7711 22593
rect 9674 22584 9680 22636
rect 9732 22624 9738 22636
rect 9953 22627 10011 22633
rect 9953 22624 9965 22627
rect 9732 22596 9965 22624
rect 9732 22584 9738 22596
rect 9953 22593 9965 22596
rect 9999 22624 10011 22627
rect 10134 22624 10140 22636
rect 9999 22596 10140 22624
rect 9999 22593 10011 22596
rect 9953 22587 10011 22593
rect 10134 22584 10140 22596
rect 10192 22584 10198 22636
rect 12250 22624 12256 22636
rect 11624 22596 12256 22624
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 1443 22528 2084 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 2056 22429 2084 22528
rect 5534 22516 5540 22568
rect 5592 22556 5598 22568
rect 5772 22559 5830 22565
rect 5772 22556 5784 22559
rect 5592 22528 5784 22556
rect 5592 22516 5598 22528
rect 5772 22525 5784 22528
rect 5818 22556 5830 22559
rect 6270 22556 6276 22568
rect 5818 22528 6276 22556
rect 5818 22525 5830 22528
rect 5772 22519 5830 22525
rect 6270 22516 6276 22528
rect 6328 22516 6334 22568
rect 6641 22559 6699 22565
rect 6641 22525 6653 22559
rect 6687 22556 6699 22559
rect 6687 22528 7236 22556
rect 6687 22525 6699 22528
rect 6641 22519 6699 22525
rect 5859 22491 5917 22497
rect 5859 22457 5871 22491
rect 5905 22488 5917 22491
rect 6730 22488 6736 22500
rect 5905 22460 6736 22488
rect 5905 22457 5917 22460
rect 5859 22451 5917 22457
rect 6730 22448 6736 22460
rect 6788 22448 6794 22500
rect 2041 22423 2099 22429
rect 2041 22389 2053 22423
rect 2087 22420 2099 22423
rect 2222 22420 2228 22432
rect 2087 22392 2228 22420
rect 2087 22389 2099 22392
rect 2041 22383 2099 22389
rect 2222 22380 2228 22392
rect 2280 22380 2286 22432
rect 7208 22420 7236 22528
rect 10778 22516 10784 22568
rect 10836 22565 10842 22568
rect 11624 22565 11652 22596
rect 12250 22584 12256 22596
rect 12308 22624 12314 22636
rect 12897 22627 12955 22633
rect 12897 22624 12909 22627
rect 12308 22596 12909 22624
rect 12308 22584 12314 22596
rect 12897 22593 12909 22596
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 10836 22559 10874 22565
rect 10862 22556 10874 22559
rect 11609 22559 11667 22565
rect 11609 22556 11621 22559
rect 10862 22528 11621 22556
rect 10862 22525 10874 22528
rect 10836 22519 10874 22525
rect 11609 22525 11621 22528
rect 11655 22525 11667 22559
rect 11609 22519 11667 22525
rect 10836 22516 10842 22519
rect 12434 22516 12440 22568
rect 12492 22556 12498 22568
rect 13265 22559 13323 22565
rect 13265 22556 13277 22559
rect 12492 22528 13277 22556
rect 12492 22516 12498 22528
rect 13265 22525 13277 22528
rect 13311 22525 13323 22559
rect 13265 22519 13323 22525
rect 13500 22559 13558 22565
rect 13500 22525 13512 22559
rect 13546 22556 13558 22559
rect 14458 22556 14464 22568
rect 13546 22528 14044 22556
rect 14422 22528 14464 22556
rect 13546 22525 13558 22528
rect 13500 22519 13558 22525
rect 14016 22500 14044 22528
rect 14458 22516 14464 22528
rect 14516 22565 14522 22568
rect 14516 22559 14570 22565
rect 14516 22525 14524 22559
rect 14558 22556 14570 22559
rect 14921 22559 14979 22565
rect 14921 22556 14933 22559
rect 14558 22528 14933 22556
rect 14558 22525 14570 22528
rect 14516 22519 14570 22525
rect 14921 22525 14933 22528
rect 14967 22525 14979 22559
rect 14921 22519 14979 22525
rect 14516 22516 14522 22519
rect 16666 22516 16672 22568
rect 16724 22556 16730 22568
rect 17012 22559 17070 22565
rect 17012 22556 17024 22559
rect 16724 22528 17024 22556
rect 16724 22516 16730 22528
rect 17012 22525 17024 22528
rect 17058 22556 17070 22559
rect 17405 22559 17463 22565
rect 17405 22556 17417 22559
rect 17058 22528 17417 22556
rect 17058 22525 17070 22528
rect 17012 22519 17070 22525
rect 17405 22525 17417 22528
rect 17451 22525 17463 22559
rect 17405 22519 17463 22525
rect 7469 22491 7527 22497
rect 7469 22457 7481 22491
rect 7515 22457 7527 22491
rect 9306 22488 9312 22500
rect 9267 22460 9312 22488
rect 7469 22451 7527 22457
rect 7484 22420 7512 22451
rect 9306 22448 9312 22460
rect 9364 22448 9370 22500
rect 9401 22491 9459 22497
rect 9401 22457 9413 22491
rect 9447 22457 9459 22491
rect 9401 22451 9459 22457
rect 7742 22420 7748 22432
rect 7208 22392 7748 22420
rect 7742 22380 7748 22392
rect 7800 22380 7806 22432
rect 8662 22380 8668 22432
rect 8720 22420 8726 22432
rect 9033 22423 9091 22429
rect 9033 22420 9045 22423
rect 8720 22392 9045 22420
rect 8720 22380 8726 22392
rect 9033 22389 9045 22392
rect 9079 22420 9091 22423
rect 9416 22420 9444 22451
rect 12802 22448 12808 22500
rect 12860 22488 12866 22500
rect 13587 22491 13645 22497
rect 13587 22488 13599 22491
rect 12860 22460 13599 22488
rect 12860 22448 12866 22460
rect 13587 22457 13599 22460
rect 13633 22457 13645 22491
rect 13998 22488 14004 22500
rect 13959 22460 14004 22488
rect 13587 22451 13645 22457
rect 13998 22448 14004 22460
rect 14056 22448 14062 22500
rect 9079 22392 9444 22420
rect 9079 22389 9091 22392
rect 9033 22383 9091 22389
rect 9858 22380 9864 22432
rect 9916 22420 9922 22432
rect 10229 22423 10287 22429
rect 10229 22420 10241 22423
rect 9916 22392 10241 22420
rect 9916 22380 9922 22392
rect 10229 22389 10241 22392
rect 10275 22389 10287 22423
rect 10229 22383 10287 22389
rect 10686 22380 10692 22432
rect 10744 22420 10750 22432
rect 10919 22423 10977 22429
rect 10919 22420 10931 22423
rect 10744 22392 10931 22420
rect 10744 22380 10750 22392
rect 10919 22389 10931 22392
rect 10965 22389 10977 22423
rect 11330 22420 11336 22432
rect 11291 22392 11336 22420
rect 10919 22383 10977 22389
rect 11330 22380 11336 22392
rect 11388 22380 11394 22432
rect 12621 22423 12679 22429
rect 12621 22389 12633 22423
rect 12667 22420 12679 22423
rect 13078 22420 13084 22432
rect 12667 22392 13084 22420
rect 12667 22389 12679 22392
rect 12621 22383 12679 22389
rect 13078 22380 13084 22392
rect 13136 22380 13142 22432
rect 15654 22420 15660 22432
rect 15615 22392 15660 22420
rect 15654 22380 15660 22392
rect 15712 22380 15718 22432
rect 24118 22380 24124 22432
rect 24176 22420 24182 22432
rect 24581 22423 24639 22429
rect 24581 22420 24593 22423
rect 24176 22392 24593 22420
rect 24176 22380 24182 22392
rect 24581 22389 24593 22392
rect 24627 22389 24639 22423
rect 24581 22383 24639 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 7466 22176 7472 22228
rect 7524 22216 7530 22228
rect 8754 22216 8760 22228
rect 7524 22188 8248 22216
rect 8715 22188 8760 22216
rect 7524 22176 7530 22188
rect 5166 22148 5172 22160
rect 5127 22120 5172 22148
rect 5166 22108 5172 22120
rect 5224 22108 5230 22160
rect 6914 22108 6920 22160
rect 6972 22148 6978 22160
rect 7377 22151 7435 22157
rect 7377 22148 7389 22151
rect 6972 22120 7389 22148
rect 6972 22108 6978 22120
rect 7377 22117 7389 22120
rect 7423 22117 7435 22151
rect 7377 22111 7435 22117
rect 6178 22040 6184 22092
rect 6236 22089 6242 22092
rect 6236 22083 6274 22089
rect 6262 22049 6274 22083
rect 8220 22080 8248 22188
rect 8754 22176 8760 22188
rect 8812 22176 8818 22228
rect 11057 22219 11115 22225
rect 11057 22185 11069 22219
rect 11103 22216 11115 22219
rect 11146 22216 11152 22228
rect 11103 22188 11152 22216
rect 11103 22185 11115 22188
rect 11057 22179 11115 22185
rect 11146 22176 11152 22188
rect 11204 22176 11210 22228
rect 12342 22216 12348 22228
rect 12303 22188 12348 22216
rect 12342 22176 12348 22188
rect 12400 22216 12406 22228
rect 12400 22188 13216 22216
rect 12400 22176 12406 22188
rect 10134 22148 10140 22160
rect 10095 22120 10140 22148
rect 10134 22108 10140 22120
rect 10192 22108 10198 22160
rect 13188 22157 13216 22188
rect 13173 22151 13231 22157
rect 13173 22117 13185 22151
rect 13219 22117 13231 22151
rect 13173 22111 13231 22117
rect 13265 22151 13323 22157
rect 13265 22117 13277 22151
rect 13311 22148 13323 22151
rect 13630 22148 13636 22160
rect 13311 22120 13636 22148
rect 13311 22117 13323 22120
rect 13265 22111 13323 22117
rect 13630 22108 13636 22120
rect 13688 22108 13694 22160
rect 15562 22108 15568 22160
rect 15620 22148 15626 22160
rect 16117 22151 16175 22157
rect 16117 22148 16129 22151
rect 15620 22120 16129 22148
rect 15620 22108 15626 22120
rect 16117 22117 16129 22120
rect 16163 22117 16175 22151
rect 16117 22111 16175 22117
rect 9122 22080 9128 22092
rect 8220 22052 9128 22080
rect 6236 22043 6274 22049
rect 6236 22040 6242 22043
rect 9122 22040 9128 22052
rect 9180 22040 9186 22092
rect 11514 22040 11520 22092
rect 11572 22089 11578 22092
rect 11572 22083 11610 22089
rect 11598 22049 11610 22083
rect 11572 22043 11610 22049
rect 11572 22040 11578 22043
rect 1670 22012 1676 22024
rect 1631 21984 1676 22012
rect 1670 21972 1676 21984
rect 1728 21972 1734 22024
rect 5534 21972 5540 22024
rect 5592 22012 5598 22024
rect 6319 22015 6377 22021
rect 6319 22012 6331 22015
rect 5592 21984 6331 22012
rect 5592 21972 5598 21984
rect 6319 21981 6331 21984
rect 6365 21981 6377 22015
rect 6319 21975 6377 21981
rect 7285 22015 7343 22021
rect 7285 21981 7297 22015
rect 7331 21981 7343 22015
rect 7558 22012 7564 22024
rect 7519 21984 7564 22012
rect 7285 21975 7343 21981
rect 7300 21944 7328 21975
rect 7558 21972 7564 21984
rect 7616 21972 7622 22024
rect 9490 21972 9496 22024
rect 9548 22012 9554 22024
rect 10045 22015 10103 22021
rect 10045 22012 10057 22015
rect 9548 21984 10057 22012
rect 9548 21972 9554 21984
rect 10045 21981 10057 21984
rect 10091 22012 10103 22015
rect 10686 22012 10692 22024
rect 10091 21984 10692 22012
rect 10091 21981 10103 21984
rect 10045 21975 10103 21981
rect 10686 21972 10692 21984
rect 10744 21972 10750 22024
rect 13446 22012 13452 22024
rect 13407 21984 13452 22012
rect 13446 21972 13452 21984
rect 13504 22012 13510 22024
rect 14277 22015 14335 22021
rect 14277 22012 14289 22015
rect 13504 21984 14289 22012
rect 13504 21972 13510 21984
rect 14277 21981 14289 21984
rect 14323 21981 14335 22015
rect 14277 21975 14335 21981
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 22012 16083 22015
rect 16942 22012 16948 22024
rect 16071 21984 16948 22012
rect 16071 21981 16083 21984
rect 16025 21975 16083 21981
rect 16942 21972 16948 21984
rect 17000 21972 17006 22024
rect 8018 21944 8024 21956
rect 7300 21916 8024 21944
rect 8018 21904 8024 21916
rect 8076 21904 8082 21956
rect 9674 21904 9680 21956
rect 9732 21944 9738 21956
rect 10597 21947 10655 21953
rect 10597 21944 10609 21947
rect 9732 21916 10609 21944
rect 9732 21904 9738 21916
rect 10597 21913 10609 21916
rect 10643 21913 10655 21947
rect 10597 21907 10655 21913
rect 15746 21904 15752 21956
rect 15804 21944 15810 21956
rect 16577 21947 16635 21953
rect 16577 21944 16589 21947
rect 15804 21916 16589 21944
rect 15804 21904 15810 21916
rect 16577 21913 16589 21916
rect 16623 21913 16635 21947
rect 16577 21907 16635 21913
rect 9306 21876 9312 21888
rect 9219 21848 9312 21876
rect 9306 21836 9312 21848
rect 9364 21876 9370 21888
rect 11655 21879 11713 21885
rect 11655 21876 11667 21879
rect 9364 21848 11667 21876
rect 9364 21836 9370 21848
rect 11655 21845 11667 21848
rect 11701 21845 11713 21879
rect 11655 21839 11713 21845
rect 12805 21879 12863 21885
rect 12805 21845 12817 21879
rect 12851 21876 12863 21879
rect 12894 21876 12900 21888
rect 12851 21848 12900 21876
rect 12851 21845 12863 21848
rect 12805 21839 12863 21845
rect 12894 21836 12900 21848
rect 12952 21836 12958 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1578 21672 1584 21684
rect 1539 21644 1584 21672
rect 1578 21632 1584 21644
rect 1636 21632 1642 21684
rect 5629 21675 5687 21681
rect 5629 21641 5641 21675
rect 5675 21672 5687 21675
rect 6178 21672 6184 21684
rect 5675 21644 6184 21672
rect 5675 21641 5687 21644
rect 5629 21635 5687 21641
rect 6178 21632 6184 21644
rect 6236 21632 6242 21684
rect 7282 21632 7288 21684
rect 7340 21672 7346 21684
rect 8297 21675 8355 21681
rect 8297 21672 8309 21675
rect 7340 21644 8309 21672
rect 7340 21632 7346 21644
rect 8297 21641 8309 21644
rect 8343 21672 8355 21675
rect 9674 21672 9680 21684
rect 8343 21644 9680 21672
rect 8343 21641 8355 21644
rect 8297 21635 8355 21641
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 9858 21632 9864 21684
rect 9916 21672 9922 21684
rect 10686 21672 10692 21684
rect 9916 21644 10692 21672
rect 9916 21632 9922 21644
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 11514 21672 11520 21684
rect 11475 21644 11520 21672
rect 11514 21632 11520 21644
rect 11572 21632 11578 21684
rect 13630 21632 13636 21684
rect 13688 21672 13694 21684
rect 13817 21675 13875 21681
rect 13817 21672 13829 21675
rect 13688 21644 13829 21672
rect 13688 21632 13694 21644
rect 13817 21641 13829 21644
rect 13863 21672 13875 21675
rect 15838 21672 15844 21684
rect 13863 21644 15844 21672
rect 13863 21641 13875 21644
rect 13817 21635 13875 21641
rect 15838 21632 15844 21644
rect 15896 21632 15902 21684
rect 24762 21672 24768 21684
rect 24723 21644 24768 21672
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 6196 21536 6224 21632
rect 8754 21564 8760 21616
rect 8812 21604 8818 21616
rect 10965 21607 11023 21613
rect 10965 21604 10977 21607
rect 8812 21576 8892 21604
rect 8812 21564 8818 21576
rect 7558 21536 7564 21548
rect 6196 21508 7564 21536
rect 7558 21496 7564 21508
rect 7616 21496 7622 21548
rect 8864 21545 8892 21576
rect 9140 21576 10977 21604
rect 9140 21548 9168 21576
rect 10965 21573 10977 21576
rect 11011 21573 11023 21607
rect 10965 21567 11023 21573
rect 13906 21564 13912 21616
rect 13964 21604 13970 21616
rect 15289 21607 15347 21613
rect 15289 21604 15301 21607
rect 13964 21576 15301 21604
rect 13964 21564 13970 21576
rect 15289 21573 15301 21576
rect 15335 21573 15347 21607
rect 15289 21567 15347 21573
rect 8849 21539 8907 21545
rect 8849 21505 8861 21539
rect 8895 21505 8907 21539
rect 9122 21536 9128 21548
rect 9083 21508 9128 21536
rect 8849 21499 8907 21505
rect 9122 21496 9128 21508
rect 9180 21496 9186 21548
rect 9858 21496 9864 21548
rect 9916 21536 9922 21548
rect 10042 21536 10048 21548
rect 9916 21508 10048 21536
rect 9916 21496 9922 21508
rect 10042 21496 10048 21508
rect 10100 21496 10106 21548
rect 10413 21539 10471 21545
rect 10413 21505 10425 21539
rect 10459 21536 10471 21539
rect 11146 21536 11152 21548
rect 10459 21508 11152 21536
rect 10459 21505 10471 21508
rect 10413 21499 10471 21505
rect 11146 21496 11152 21508
rect 11204 21496 11210 21548
rect 12253 21539 12311 21545
rect 12253 21505 12265 21539
rect 12299 21536 12311 21539
rect 12802 21536 12808 21548
rect 12299 21508 12808 21536
rect 12299 21505 12311 21508
rect 12253 21499 12311 21505
rect 12802 21496 12808 21508
rect 12860 21496 12866 21548
rect 13446 21536 13452 21548
rect 13407 21508 13452 21536
rect 13446 21496 13452 21508
rect 13504 21536 13510 21548
rect 14366 21536 14372 21548
rect 13504 21508 14372 21536
rect 13504 21496 13510 21508
rect 14366 21496 14372 21508
rect 14424 21496 14430 21548
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21468 1455 21471
rect 2038 21468 2044 21480
rect 1443 21440 2044 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 2038 21428 2044 21440
rect 2096 21428 2102 21480
rect 4592 21471 4650 21477
rect 4592 21437 4604 21471
rect 4638 21468 4650 21471
rect 5788 21471 5846 21477
rect 4638 21440 5120 21468
rect 4638 21437 4650 21440
rect 4592 21431 4650 21437
rect 5092 21344 5120 21440
rect 5788 21437 5800 21471
rect 5834 21468 5846 21471
rect 5834 21440 6316 21468
rect 5834 21437 5846 21440
rect 5788 21431 5846 21437
rect 6288 21412 6316 21440
rect 6270 21400 6276 21412
rect 6231 21372 6276 21400
rect 6270 21360 6276 21372
rect 6328 21360 6334 21412
rect 7282 21400 7288 21412
rect 7243 21372 7288 21400
rect 7282 21360 7288 21372
rect 7340 21360 7346 21412
rect 7374 21360 7380 21412
rect 7432 21400 7438 21412
rect 8941 21403 8999 21409
rect 7432 21372 7525 21400
rect 7432 21360 7466 21372
rect 8941 21369 8953 21403
rect 8987 21369 8999 21403
rect 10505 21403 10563 21409
rect 10505 21400 10517 21403
rect 8941 21363 8999 21369
rect 10152 21372 10517 21400
rect 4430 21292 4436 21344
rect 4488 21332 4494 21344
rect 4663 21335 4721 21341
rect 4663 21332 4675 21335
rect 4488 21304 4675 21332
rect 4488 21292 4494 21304
rect 4663 21301 4675 21304
rect 4709 21301 4721 21335
rect 5074 21332 5080 21344
rect 5035 21304 5080 21332
rect 4663 21295 4721 21301
rect 5074 21292 5080 21304
rect 5132 21292 5138 21344
rect 5859 21335 5917 21341
rect 5859 21301 5871 21335
rect 5905 21332 5917 21335
rect 5994 21332 6000 21344
rect 5905 21304 6000 21332
rect 5905 21301 5917 21304
rect 5859 21295 5917 21301
rect 5994 21292 6000 21304
rect 6052 21292 6058 21344
rect 6641 21335 6699 21341
rect 6641 21301 6653 21335
rect 6687 21332 6699 21335
rect 6822 21332 6828 21344
rect 6687 21304 6828 21332
rect 6687 21301 6699 21304
rect 6641 21295 6699 21301
rect 6822 21292 6828 21304
rect 6880 21292 6886 21344
rect 7101 21335 7159 21341
rect 7101 21301 7113 21335
rect 7147 21332 7159 21335
rect 7438 21332 7466 21360
rect 8662 21332 8668 21344
rect 7147 21304 7466 21332
rect 8623 21304 8668 21332
rect 7147 21301 7159 21304
rect 7101 21295 7159 21301
rect 8662 21292 8668 21304
rect 8720 21332 8726 21344
rect 8956 21332 8984 21363
rect 8720 21304 8984 21332
rect 9861 21335 9919 21341
rect 8720 21292 8726 21304
rect 9861 21301 9873 21335
rect 9907 21332 9919 21335
rect 10042 21332 10048 21344
rect 9907 21304 10048 21332
rect 9907 21301 9919 21304
rect 9861 21295 9919 21301
rect 10042 21292 10048 21304
rect 10100 21332 10106 21344
rect 10152 21341 10180 21372
rect 10505 21369 10517 21372
rect 10551 21369 10563 21403
rect 12894 21400 12900 21412
rect 12807 21372 12900 21400
rect 10505 21363 10563 21369
rect 12894 21360 12900 21372
rect 12952 21400 12958 21412
rect 13538 21400 13544 21412
rect 12952 21372 13544 21400
rect 12952 21360 12958 21372
rect 13538 21360 13544 21372
rect 13596 21360 13602 21412
rect 14461 21403 14519 21409
rect 14461 21369 14473 21403
rect 14507 21369 14519 21403
rect 15010 21400 15016 21412
rect 14971 21372 15016 21400
rect 14461 21363 14519 21369
rect 10137 21335 10195 21341
rect 10137 21332 10149 21335
rect 10100 21304 10149 21332
rect 10100 21292 10106 21304
rect 10137 21301 10149 21304
rect 10183 21301 10195 21335
rect 14182 21332 14188 21344
rect 14095 21304 14188 21332
rect 10137 21295 10195 21301
rect 14182 21292 14188 21304
rect 14240 21332 14246 21344
rect 14476 21332 14504 21363
rect 15010 21360 15016 21372
rect 15068 21360 15074 21412
rect 15304 21400 15332 21567
rect 16114 21564 16120 21616
rect 16172 21604 16178 21616
rect 16485 21607 16543 21613
rect 16485 21604 16497 21607
rect 16172 21576 16497 21604
rect 16172 21564 16178 21576
rect 16485 21573 16497 21576
rect 16531 21573 16543 21607
rect 16485 21567 16543 21573
rect 15930 21536 15936 21548
rect 15843 21508 15936 21536
rect 15930 21496 15936 21508
rect 15988 21536 15994 21548
rect 17221 21539 17279 21545
rect 17221 21536 17233 21539
rect 15988 21508 17233 21536
rect 15988 21496 15994 21508
rect 17221 21505 17233 21508
rect 17267 21505 17279 21539
rect 17221 21499 17279 21505
rect 18138 21477 18144 21480
rect 18116 21471 18144 21477
rect 18116 21468 18128 21471
rect 18051 21440 18128 21468
rect 18116 21437 18128 21440
rect 18196 21468 18202 21480
rect 24581 21471 24639 21477
rect 18196 21440 18644 21468
rect 18116 21431 18144 21437
rect 18138 21428 18144 21431
rect 18196 21428 18202 21440
rect 16025 21403 16083 21409
rect 16025 21400 16037 21403
rect 15304 21372 16037 21400
rect 16025 21369 16037 21372
rect 16071 21400 16083 21403
rect 16758 21400 16764 21412
rect 16071 21372 16764 21400
rect 16071 21369 16083 21372
rect 16025 21363 16083 21369
rect 16758 21360 16764 21372
rect 16816 21360 16822 21412
rect 16942 21400 16948 21412
rect 16855 21372 16948 21400
rect 16942 21360 16948 21372
rect 17000 21400 17006 21412
rect 17862 21400 17868 21412
rect 17000 21372 17868 21400
rect 17000 21360 17006 21372
rect 17862 21360 17868 21372
rect 17920 21360 17926 21412
rect 14240 21304 14504 21332
rect 14240 21292 14246 21304
rect 15562 21292 15568 21344
rect 15620 21332 15626 21344
rect 15749 21335 15807 21341
rect 15749 21332 15761 21335
rect 15620 21304 15761 21332
rect 15620 21292 15626 21304
rect 15749 21301 15761 21304
rect 15795 21332 15807 21335
rect 16850 21332 16856 21344
rect 15795 21304 16856 21332
rect 15795 21301 15807 21304
rect 15749 21295 15807 21301
rect 16850 21292 16856 21304
rect 16908 21292 16914 21344
rect 17494 21292 17500 21344
rect 17552 21332 17558 21344
rect 18616 21341 18644 21440
rect 24581 21437 24593 21471
rect 24627 21437 24639 21471
rect 24581 21431 24639 21437
rect 18187 21335 18245 21341
rect 18187 21332 18199 21335
rect 17552 21304 18199 21332
rect 17552 21292 17558 21304
rect 18187 21301 18199 21304
rect 18233 21301 18245 21335
rect 18187 21295 18245 21301
rect 18601 21335 18659 21341
rect 18601 21301 18613 21335
rect 18647 21332 18659 21335
rect 18782 21332 18788 21344
rect 18647 21304 18788 21332
rect 18647 21301 18659 21304
rect 18601 21295 18659 21301
rect 18782 21292 18788 21304
rect 18840 21292 18846 21344
rect 24210 21292 24216 21344
rect 24268 21332 24274 21344
rect 24596 21332 24624 21431
rect 25133 21335 25191 21341
rect 25133 21332 25145 21335
rect 24268 21304 25145 21332
rect 24268 21292 24274 21304
rect 25133 21301 25145 21304
rect 25179 21301 25191 21335
rect 25133 21295 25191 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 5258 21128 5264 21140
rect 5219 21100 5264 21128
rect 5258 21088 5264 21100
rect 5316 21088 5322 21140
rect 7374 21128 7380 21140
rect 7335 21100 7380 21128
rect 7374 21088 7380 21100
rect 7432 21088 7438 21140
rect 8018 21128 8024 21140
rect 7979 21100 8024 21128
rect 8018 21088 8024 21100
rect 8076 21088 8082 21140
rect 8711 21131 8769 21137
rect 8711 21097 8723 21131
rect 8757 21128 8769 21131
rect 9766 21128 9772 21140
rect 8757 21100 9772 21128
rect 8757 21097 8769 21100
rect 8711 21091 8769 21097
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 15838 21088 15844 21140
rect 15896 21128 15902 21140
rect 15896 21100 16068 21128
rect 15896 21088 15902 21100
rect 6638 21020 6644 21072
rect 6696 21060 6702 21072
rect 6778 21063 6836 21069
rect 6778 21060 6790 21063
rect 6696 21032 6790 21060
rect 6696 21020 6702 21032
rect 6778 21029 6790 21032
rect 6824 21029 6836 21063
rect 9490 21060 9496 21072
rect 9451 21032 9496 21060
rect 6778 21023 6836 21029
rect 9490 21020 9496 21032
rect 9548 21020 9554 21072
rect 10597 21063 10655 21069
rect 10597 21029 10609 21063
rect 10643 21060 10655 21063
rect 10686 21060 10692 21072
rect 10643 21032 10692 21060
rect 10643 21029 10655 21032
rect 10597 21023 10655 21029
rect 10686 21020 10692 21032
rect 10744 21020 10750 21072
rect 13817 21063 13875 21069
rect 13817 21029 13829 21063
rect 13863 21060 13875 21063
rect 13906 21060 13912 21072
rect 13863 21032 13912 21060
rect 13863 21029 13875 21032
rect 13817 21023 13875 21029
rect 13906 21020 13912 21032
rect 13964 21020 13970 21072
rect 14366 21060 14372 21072
rect 14327 21032 14372 21060
rect 14366 21020 14372 21032
rect 14424 21020 14430 21072
rect 15654 21020 15660 21072
rect 15712 21060 15718 21072
rect 16040 21069 16068 21100
rect 16758 21088 16764 21140
rect 16816 21128 16822 21140
rect 16816 21100 17632 21128
rect 16816 21088 16822 21100
rect 15933 21063 15991 21069
rect 15933 21060 15945 21063
rect 15712 21032 15945 21060
rect 15712 21020 15718 21032
rect 15933 21029 15945 21032
rect 15979 21029 15991 21063
rect 15933 21023 15991 21029
rect 16025 21063 16083 21069
rect 16025 21029 16037 21063
rect 16071 21029 16083 21063
rect 17494 21060 17500 21072
rect 17455 21032 17500 21060
rect 16025 21023 16083 21029
rect 17494 21020 17500 21032
rect 17552 21020 17558 21072
rect 17604 21069 17632 21100
rect 17589 21063 17647 21069
rect 17589 21029 17601 21063
rect 17635 21029 17647 21063
rect 17589 21023 17647 21029
rect 4433 20995 4491 21001
rect 4433 20961 4445 20995
rect 4479 20992 4491 20995
rect 4706 20992 4712 21004
rect 4479 20964 4712 20992
rect 4479 20961 4491 20964
rect 4433 20955 4491 20961
rect 4706 20952 4712 20964
rect 4764 20952 4770 21004
rect 5074 20952 5080 21004
rect 5132 20992 5138 21004
rect 5512 20995 5570 21001
rect 5512 20992 5524 20995
rect 5132 20964 5524 20992
rect 5132 20952 5138 20964
rect 5512 20961 5524 20964
rect 5558 20992 5570 20995
rect 6086 20992 6092 21004
rect 5558 20964 6092 20992
rect 5558 20961 5570 20964
rect 5512 20955 5570 20961
rect 6086 20952 6092 20964
rect 6144 20952 6150 21004
rect 8640 20995 8698 21001
rect 8640 20961 8652 20995
rect 8686 20992 8698 20995
rect 8846 20992 8852 21004
rect 8686 20964 8852 20992
rect 8686 20961 8698 20964
rect 8640 20955 8698 20961
rect 8846 20952 8852 20964
rect 8904 20952 8910 21004
rect 11146 20952 11152 21004
rect 11204 20992 11210 21004
rect 12066 20992 12072 21004
rect 11204 20964 11249 20992
rect 12027 20964 12072 20992
rect 11204 20952 11210 20964
rect 12066 20952 12072 20964
rect 12124 20952 12130 21004
rect 12618 20992 12624 21004
rect 12579 20964 12624 20992
rect 12618 20952 12624 20964
rect 12676 20952 12682 21004
rect 5626 20884 5632 20936
rect 5684 20924 5690 20936
rect 6273 20927 6331 20933
rect 6273 20924 6285 20927
rect 5684 20896 6285 20924
rect 5684 20884 5690 20896
rect 6273 20893 6285 20896
rect 6319 20924 6331 20927
rect 6457 20927 6515 20933
rect 6457 20924 6469 20927
rect 6319 20896 6469 20924
rect 6319 20893 6331 20896
rect 6273 20887 6331 20893
rect 6457 20893 6469 20896
rect 6503 20893 6515 20927
rect 6457 20887 6515 20893
rect 10505 20927 10563 20933
rect 10505 20893 10517 20927
rect 10551 20924 10563 20927
rect 10686 20924 10692 20936
rect 10551 20896 10692 20924
rect 10551 20893 10563 20896
rect 10505 20887 10563 20893
rect 10686 20884 10692 20896
rect 10744 20884 10750 20936
rect 12805 20927 12863 20933
rect 12805 20893 12817 20927
rect 12851 20924 12863 20927
rect 13262 20924 13268 20936
rect 12851 20896 13268 20924
rect 12851 20893 12863 20896
rect 12805 20887 12863 20893
rect 13262 20884 13268 20896
rect 13320 20884 13326 20936
rect 13722 20924 13728 20936
rect 13683 20896 13728 20924
rect 13722 20884 13728 20896
rect 13780 20884 13786 20936
rect 16114 20884 16120 20936
rect 16172 20924 16178 20936
rect 16209 20927 16267 20933
rect 16209 20924 16221 20927
rect 16172 20896 16221 20924
rect 16172 20884 16178 20896
rect 16209 20893 16221 20896
rect 16255 20893 16267 20927
rect 16209 20887 16267 20893
rect 17773 20927 17831 20933
rect 17773 20893 17785 20927
rect 17819 20893 17831 20927
rect 17773 20887 17831 20893
rect 17788 20856 17816 20887
rect 15764 20828 17816 20856
rect 15764 20800 15792 20828
rect 4154 20748 4160 20800
rect 4212 20788 4218 20800
rect 4617 20791 4675 20797
rect 4617 20788 4629 20791
rect 4212 20760 4629 20788
rect 4212 20748 4218 20760
rect 4617 20757 4629 20760
rect 4663 20757 4675 20791
rect 4617 20751 4675 20757
rect 5583 20791 5641 20797
rect 5583 20757 5595 20791
rect 5629 20788 5641 20791
rect 6546 20788 6552 20800
rect 5629 20760 6552 20788
rect 5629 20757 5641 20760
rect 5583 20751 5641 20757
rect 6546 20748 6552 20760
rect 6604 20748 6610 20800
rect 7006 20748 7012 20800
rect 7064 20788 7070 20800
rect 7653 20791 7711 20797
rect 7653 20788 7665 20791
rect 7064 20760 7665 20788
rect 7064 20748 7070 20760
rect 7653 20757 7665 20760
rect 7699 20757 7711 20791
rect 9030 20788 9036 20800
rect 8991 20760 9036 20788
rect 7653 20751 7711 20757
rect 9030 20748 9036 20760
rect 9088 20748 9094 20800
rect 10042 20748 10048 20800
rect 10100 20788 10106 20800
rect 10137 20791 10195 20797
rect 10137 20788 10149 20791
rect 10100 20760 10149 20788
rect 10100 20748 10106 20760
rect 10137 20757 10149 20760
rect 10183 20757 10195 20791
rect 15746 20788 15752 20800
rect 15707 20760 15752 20788
rect 10137 20751 10195 20757
rect 15746 20748 15752 20760
rect 15804 20748 15810 20800
rect 16574 20748 16580 20800
rect 16632 20788 16638 20800
rect 16853 20791 16911 20797
rect 16853 20788 16865 20791
rect 16632 20760 16865 20788
rect 16632 20748 16638 20760
rect 16853 20757 16865 20760
rect 16899 20757 16911 20791
rect 16853 20751 16911 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 3329 20587 3387 20593
rect 3329 20553 3341 20587
rect 3375 20584 3387 20587
rect 6362 20584 6368 20596
rect 3375 20556 6368 20584
rect 3375 20553 3387 20556
rect 3329 20547 3387 20553
rect 1811 20519 1869 20525
rect 1811 20485 1823 20519
rect 1857 20516 1869 20519
rect 2406 20516 2412 20528
rect 1857 20488 2412 20516
rect 1857 20485 1869 20488
rect 1811 20479 1869 20485
rect 2406 20476 2412 20488
rect 2464 20476 2470 20528
rect 1740 20383 1798 20389
rect 1740 20349 1752 20383
rect 1786 20380 1798 20383
rect 2844 20383 2902 20389
rect 1786 20352 1992 20380
rect 1786 20349 1798 20352
rect 1740 20343 1798 20349
rect 1964 20256 1992 20352
rect 2844 20349 2856 20383
rect 2890 20380 2902 20383
rect 3344 20380 3372 20547
rect 6362 20544 6368 20556
rect 6420 20544 6426 20596
rect 7742 20584 7748 20596
rect 7703 20556 7748 20584
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 8481 20587 8539 20593
rect 8481 20553 8493 20587
rect 8527 20584 8539 20587
rect 8846 20584 8852 20596
rect 8527 20556 8852 20584
rect 8527 20553 8539 20556
rect 8481 20547 8539 20553
rect 8846 20544 8852 20556
rect 8904 20544 8910 20596
rect 9950 20584 9956 20596
rect 9911 20556 9956 20584
rect 9950 20544 9956 20556
rect 10008 20544 10014 20596
rect 10778 20544 10784 20596
rect 10836 20584 10842 20596
rect 11149 20587 11207 20593
rect 11149 20584 11161 20587
rect 10836 20556 11161 20584
rect 10836 20544 10842 20556
rect 11149 20553 11161 20556
rect 11195 20553 11207 20587
rect 12066 20584 12072 20596
rect 12027 20556 12072 20584
rect 11149 20547 11207 20553
rect 12066 20544 12072 20556
rect 12124 20544 12130 20596
rect 12618 20584 12624 20596
rect 12579 20556 12624 20584
rect 12618 20544 12624 20556
rect 12676 20544 12682 20596
rect 14182 20584 14188 20596
rect 14143 20556 14188 20584
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 15654 20544 15660 20596
rect 15712 20584 15718 20596
rect 15841 20587 15899 20593
rect 15841 20584 15853 20587
rect 15712 20556 15853 20584
rect 15712 20544 15718 20556
rect 15841 20553 15853 20556
rect 15887 20553 15899 20587
rect 15841 20547 15899 20553
rect 16758 20544 16764 20596
rect 16816 20584 16822 20596
rect 17405 20587 17463 20593
rect 17405 20584 17417 20587
rect 16816 20556 17417 20584
rect 16816 20544 16822 20556
rect 17405 20553 17417 20556
rect 17451 20553 17463 20587
rect 17405 20547 17463 20553
rect 17494 20544 17500 20596
rect 17552 20584 17558 20596
rect 17773 20587 17831 20593
rect 17773 20584 17785 20587
rect 17552 20556 17785 20584
rect 17552 20544 17558 20556
rect 17773 20553 17785 20556
rect 17819 20553 17831 20587
rect 17773 20547 17831 20553
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 18187 20587 18245 20593
rect 18187 20584 18199 20587
rect 18012 20556 18199 20584
rect 18012 20544 18018 20556
rect 18187 20553 18199 20556
rect 18233 20553 18245 20587
rect 18187 20547 18245 20553
rect 6086 20476 6092 20528
rect 6144 20516 6150 20528
rect 6273 20519 6331 20525
rect 6273 20516 6285 20519
rect 6144 20488 6285 20516
rect 6144 20476 6150 20488
rect 6273 20485 6285 20488
rect 6319 20516 6331 20519
rect 6822 20516 6828 20528
rect 6319 20488 6828 20516
rect 6319 20485 6331 20488
rect 6273 20479 6331 20485
rect 6822 20476 6828 20488
rect 6880 20476 6886 20528
rect 8665 20451 8723 20457
rect 8665 20417 8677 20451
rect 8711 20448 8723 20451
rect 9030 20448 9036 20460
rect 8711 20420 9036 20448
rect 8711 20417 8723 20420
rect 8665 20411 8723 20417
rect 9030 20408 9036 20420
rect 9088 20408 9094 20460
rect 9122 20408 9128 20460
rect 9180 20448 9186 20460
rect 9968 20448 9996 20544
rect 10229 20451 10287 20457
rect 10229 20448 10241 20451
rect 9180 20420 9225 20448
rect 9968 20420 10241 20448
rect 9180 20408 9186 20420
rect 10229 20417 10241 20420
rect 10275 20417 10287 20451
rect 10502 20448 10508 20460
rect 10463 20420 10508 20448
rect 10229 20411 10287 20417
rect 10502 20408 10508 20420
rect 10560 20448 10566 20460
rect 10870 20448 10876 20460
rect 10560 20420 10876 20448
rect 10560 20408 10566 20420
rect 10870 20408 10876 20420
rect 10928 20408 10934 20460
rect 13262 20448 13268 20460
rect 13223 20420 13268 20448
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 15562 20448 15568 20460
rect 15523 20420 15568 20448
rect 15562 20408 15568 20420
rect 15620 20408 15626 20460
rect 16666 20448 16672 20460
rect 16627 20420 16672 20448
rect 16666 20408 16672 20420
rect 16724 20408 16730 20460
rect 2890 20352 3372 20380
rect 2890 20349 2902 20352
rect 2844 20343 2902 20349
rect 3786 20340 3792 20392
rect 3844 20389 3850 20392
rect 3844 20383 3882 20389
rect 3870 20380 3882 20383
rect 4249 20383 4307 20389
rect 4249 20380 4261 20383
rect 3870 20352 4261 20380
rect 3870 20349 3882 20352
rect 3844 20343 3882 20349
rect 4249 20349 4261 20352
rect 4295 20349 4307 20383
rect 4249 20343 4307 20349
rect 3844 20340 3850 20343
rect 4890 20340 4896 20392
rect 4948 20380 4954 20392
rect 5077 20383 5135 20389
rect 5077 20380 5089 20383
rect 4948 20352 5089 20380
rect 4948 20340 4954 20352
rect 5077 20349 5089 20352
rect 5123 20380 5135 20383
rect 5169 20383 5227 20389
rect 5169 20380 5181 20383
rect 5123 20352 5181 20380
rect 5123 20349 5135 20352
rect 5077 20343 5135 20349
rect 5169 20349 5181 20352
rect 5215 20349 5227 20383
rect 5169 20343 5227 20349
rect 5258 20340 5264 20392
rect 5316 20380 5322 20392
rect 5629 20383 5687 20389
rect 5629 20380 5641 20383
rect 5316 20352 5641 20380
rect 5316 20340 5322 20352
rect 5629 20349 5641 20352
rect 5675 20349 5687 20383
rect 5629 20343 5687 20349
rect 6086 20340 6092 20392
rect 6144 20380 6150 20392
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 6144 20352 6837 20380
rect 6144 20340 6150 20352
rect 6825 20349 6837 20352
rect 6871 20380 6883 20383
rect 7006 20380 7012 20392
rect 6871 20352 7012 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 7006 20340 7012 20352
rect 7064 20340 7070 20392
rect 14734 20340 14740 20392
rect 14792 20380 14798 20392
rect 15080 20383 15138 20389
rect 15080 20380 15092 20383
rect 14792 20352 15092 20380
rect 14792 20340 14798 20352
rect 15080 20349 15092 20352
rect 15126 20380 15138 20383
rect 15580 20380 15608 20408
rect 15126 20352 15608 20380
rect 18116 20383 18174 20389
rect 15126 20349 15138 20352
rect 15080 20343 15138 20349
rect 18116 20349 18128 20383
rect 18162 20380 18174 20383
rect 18690 20380 18696 20392
rect 18162 20352 18696 20380
rect 18162 20349 18174 20352
rect 18116 20343 18174 20349
rect 5902 20312 5908 20324
rect 5863 20284 5908 20312
rect 5902 20272 5908 20284
rect 5960 20272 5966 20324
rect 7146 20315 7204 20321
rect 7146 20312 7158 20315
rect 6656 20284 7158 20312
rect 6656 20256 6684 20284
rect 7146 20281 7158 20284
rect 7192 20312 7204 20315
rect 8021 20315 8079 20321
rect 8021 20312 8033 20315
rect 7192 20284 8033 20312
rect 7192 20281 7204 20284
rect 7146 20275 7204 20281
rect 8021 20281 8033 20284
rect 8067 20281 8079 20315
rect 8754 20312 8760 20324
rect 8715 20284 8760 20312
rect 8021 20275 8079 20281
rect 8754 20272 8760 20284
rect 8812 20272 8818 20324
rect 10042 20272 10048 20324
rect 10100 20312 10106 20324
rect 10321 20315 10379 20321
rect 10321 20312 10333 20315
rect 10100 20284 10333 20312
rect 10100 20272 10106 20284
rect 10321 20281 10333 20284
rect 10367 20281 10379 20315
rect 13586 20315 13644 20321
rect 13586 20312 13598 20315
rect 10321 20275 10379 20281
rect 13464 20284 13598 20312
rect 13464 20256 13492 20284
rect 13586 20281 13598 20284
rect 13632 20281 13644 20315
rect 13586 20275 13644 20281
rect 15746 20272 15752 20324
rect 15804 20312 15810 20324
rect 16209 20315 16267 20321
rect 16209 20312 16221 20315
rect 15804 20284 16221 20312
rect 15804 20272 15810 20284
rect 16209 20281 16221 20284
rect 16255 20281 16267 20315
rect 16209 20275 16267 20281
rect 16301 20315 16359 20321
rect 16301 20281 16313 20315
rect 16347 20312 16359 20315
rect 16482 20312 16488 20324
rect 16347 20284 16488 20312
rect 16347 20281 16359 20284
rect 16301 20275 16359 20281
rect 1946 20204 1952 20256
rect 2004 20244 2010 20256
rect 2133 20247 2191 20253
rect 2133 20244 2145 20247
rect 2004 20216 2145 20244
rect 2004 20204 2010 20216
rect 2133 20213 2145 20216
rect 2179 20213 2191 20247
rect 2133 20207 2191 20213
rect 2915 20247 2973 20253
rect 2915 20213 2927 20247
rect 2961 20244 2973 20247
rect 3142 20244 3148 20256
rect 2961 20216 3148 20244
rect 2961 20213 2973 20216
rect 2915 20207 2973 20213
rect 3142 20204 3148 20216
rect 3200 20204 3206 20256
rect 3878 20204 3884 20256
rect 3936 20253 3942 20256
rect 3936 20247 3985 20253
rect 3936 20213 3939 20247
rect 3973 20213 3985 20247
rect 4706 20244 4712 20256
rect 4619 20216 4712 20244
rect 3936 20207 3985 20213
rect 3936 20204 3942 20207
rect 4706 20204 4712 20216
rect 4764 20244 4770 20256
rect 5442 20244 5448 20256
rect 4764 20216 5448 20244
rect 4764 20204 4770 20216
rect 5442 20204 5448 20216
rect 5500 20204 5506 20256
rect 6638 20244 6644 20256
rect 6599 20216 6644 20244
rect 6638 20204 6644 20216
rect 6696 20204 6702 20256
rect 9677 20247 9735 20253
rect 9677 20213 9689 20247
rect 9723 20244 9735 20247
rect 10686 20244 10692 20256
rect 9723 20216 10692 20244
rect 9723 20213 9735 20216
rect 9677 20207 9735 20213
rect 10686 20204 10692 20216
rect 10744 20204 10750 20256
rect 13173 20247 13231 20253
rect 13173 20213 13185 20247
rect 13219 20244 13231 20247
rect 13446 20244 13452 20256
rect 13219 20216 13452 20244
rect 13219 20213 13231 20216
rect 13173 20207 13231 20213
rect 13446 20204 13452 20216
rect 13504 20204 13510 20256
rect 14458 20244 14464 20256
rect 14419 20216 14464 20244
rect 14458 20204 14464 20216
rect 14516 20204 14522 20256
rect 14826 20204 14832 20256
rect 14884 20244 14890 20256
rect 15151 20247 15209 20253
rect 15151 20244 15163 20247
rect 14884 20216 15163 20244
rect 14884 20204 14890 20216
rect 15151 20213 15163 20216
rect 15197 20213 15209 20247
rect 16224 20244 16252 20275
rect 16482 20272 16488 20284
rect 16540 20272 16546 20324
rect 18524 20256 18552 20352
rect 18690 20340 18696 20352
rect 18748 20340 18754 20392
rect 19058 20340 19064 20392
rect 19116 20389 19122 20392
rect 19116 20383 19154 20389
rect 19142 20380 19154 20383
rect 19521 20383 19579 20389
rect 19521 20380 19533 20383
rect 19142 20352 19533 20380
rect 19142 20349 19154 20352
rect 19116 20343 19154 20349
rect 19521 20349 19533 20352
rect 19567 20349 19579 20383
rect 19521 20343 19579 20349
rect 19116 20340 19122 20343
rect 16574 20244 16580 20256
rect 16224 20216 16580 20244
rect 15151 20207 15209 20213
rect 16574 20204 16580 20216
rect 16632 20204 16638 20256
rect 18506 20244 18512 20256
rect 18467 20216 18512 20244
rect 18506 20204 18512 20216
rect 18564 20204 18570 20256
rect 19199 20247 19257 20253
rect 19199 20213 19211 20247
rect 19245 20244 19257 20247
rect 19978 20244 19984 20256
rect 19245 20216 19984 20244
rect 19245 20213 19257 20216
rect 19199 20207 19257 20213
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 6914 20000 6920 20052
rect 6972 20040 6978 20052
rect 7285 20043 7343 20049
rect 7285 20040 7297 20043
rect 6972 20012 7297 20040
rect 6972 20000 6978 20012
rect 7285 20009 7297 20012
rect 7331 20009 7343 20043
rect 7285 20003 7343 20009
rect 8711 20043 8769 20049
rect 8711 20009 8723 20043
rect 8757 20040 8769 20043
rect 9030 20040 9036 20052
rect 8757 20012 9036 20040
rect 8757 20009 8769 20012
rect 8711 20003 8769 20009
rect 9030 20000 9036 20012
rect 9088 20000 9094 20052
rect 10686 20000 10692 20052
rect 10744 20040 10750 20052
rect 11563 20043 11621 20049
rect 11563 20040 11575 20043
rect 10744 20012 11575 20040
rect 10744 20000 10750 20012
rect 11563 20009 11575 20012
rect 11609 20009 11621 20043
rect 11563 20003 11621 20009
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 14093 20043 14151 20049
rect 14093 20040 14105 20043
rect 13872 20012 14105 20040
rect 13872 20000 13878 20012
rect 14093 20009 14105 20012
rect 14139 20009 14151 20043
rect 15838 20040 15844 20052
rect 15799 20012 15844 20040
rect 14093 20003 14151 20009
rect 15838 20000 15844 20012
rect 15896 20000 15902 20052
rect 5534 19972 5540 19984
rect 5495 19944 5540 19972
rect 5534 19932 5540 19944
rect 5592 19932 5598 19984
rect 6638 19932 6644 19984
rect 6696 19981 6702 19984
rect 6696 19975 6744 19981
rect 6696 19941 6698 19975
rect 6732 19941 6744 19975
rect 6696 19935 6744 19941
rect 6696 19932 6702 19935
rect 9950 19932 9956 19984
rect 10008 19981 10014 19984
rect 10008 19975 10056 19981
rect 10008 19941 10010 19975
rect 10044 19941 10056 19975
rect 10008 19935 10056 19941
rect 13259 19975 13317 19981
rect 13259 19941 13271 19975
rect 13305 19972 13317 19975
rect 13446 19972 13452 19984
rect 13305 19944 13452 19972
rect 13305 19941 13317 19944
rect 13259 19935 13317 19941
rect 10008 19932 10014 19935
rect 13446 19932 13452 19944
rect 13504 19932 13510 19984
rect 16206 19972 16212 19984
rect 16167 19944 16212 19972
rect 16206 19932 16212 19944
rect 16264 19932 16270 19984
rect 16850 19932 16856 19984
rect 16908 19972 16914 19984
rect 17773 19975 17831 19981
rect 17773 19972 17785 19975
rect 16908 19944 17785 19972
rect 16908 19932 16914 19944
rect 17773 19941 17785 19944
rect 17819 19972 17831 19975
rect 17862 19972 17868 19984
rect 17819 19944 17868 19972
rect 17819 19941 17831 19944
rect 17773 19935 17831 19941
rect 17862 19932 17868 19944
rect 17920 19932 17926 19984
rect 1464 19907 1522 19913
rect 1464 19873 1476 19907
rect 1510 19904 1522 19907
rect 1854 19904 1860 19916
rect 1510 19876 1860 19904
rect 1510 19873 1522 19876
rect 1464 19867 1522 19873
rect 1854 19864 1860 19876
rect 1912 19864 1918 19916
rect 2961 19907 3019 19913
rect 2961 19873 2973 19907
rect 3007 19904 3019 19907
rect 3050 19904 3056 19916
rect 3007 19876 3056 19904
rect 3007 19873 3019 19876
rect 2961 19867 3019 19873
rect 3050 19864 3056 19876
rect 3108 19904 3114 19916
rect 4154 19904 4160 19916
rect 3108 19876 4160 19904
rect 3108 19864 3114 19876
rect 4154 19864 4160 19876
rect 4212 19864 4218 19916
rect 5074 19904 5080 19916
rect 5035 19876 5080 19904
rect 5074 19864 5080 19876
rect 5132 19864 5138 19916
rect 5258 19904 5264 19916
rect 5219 19876 5264 19904
rect 5258 19864 5264 19876
rect 5316 19904 5322 19916
rect 5813 19907 5871 19913
rect 5813 19904 5825 19907
rect 5316 19876 5825 19904
rect 5316 19864 5322 19876
rect 5813 19873 5825 19876
rect 5859 19873 5871 19907
rect 5813 19867 5871 19873
rect 8640 19907 8698 19913
rect 8640 19873 8652 19907
rect 8686 19904 8698 19907
rect 9398 19904 9404 19916
rect 8686 19876 9404 19904
rect 8686 19873 8698 19876
rect 8640 19867 8698 19873
rect 9398 19864 9404 19876
rect 9456 19864 9462 19916
rect 9674 19904 9680 19916
rect 9635 19876 9680 19904
rect 9674 19864 9680 19876
rect 9732 19864 9738 19916
rect 10597 19907 10655 19913
rect 10597 19873 10609 19907
rect 10643 19904 10655 19907
rect 10778 19904 10784 19916
rect 10643 19876 10784 19904
rect 10643 19873 10655 19876
rect 10597 19867 10655 19873
rect 6178 19796 6184 19848
rect 6236 19836 6242 19848
rect 6365 19839 6423 19845
rect 6365 19836 6377 19839
rect 6236 19808 6377 19836
rect 6236 19796 6242 19808
rect 6365 19805 6377 19808
rect 6411 19805 6423 19839
rect 6365 19799 6423 19805
rect 8754 19796 8760 19848
rect 8812 19836 8818 19848
rect 9125 19839 9183 19845
rect 9125 19836 9137 19839
rect 8812 19808 9137 19836
rect 8812 19796 8818 19808
rect 9125 19805 9137 19808
rect 9171 19836 9183 19839
rect 10612 19836 10640 19867
rect 10778 19864 10784 19876
rect 10836 19864 10842 19916
rect 11492 19907 11550 19913
rect 11492 19873 11504 19907
rect 11538 19904 11550 19907
rect 11974 19904 11980 19916
rect 11538 19876 11980 19904
rect 11538 19873 11550 19876
rect 11492 19867 11550 19873
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 13817 19907 13875 19913
rect 13817 19873 13829 19907
rect 13863 19904 13875 19907
rect 13906 19904 13912 19916
rect 13863 19876 13912 19904
rect 13863 19873 13875 19876
rect 13817 19867 13875 19873
rect 13906 19864 13912 19876
rect 13964 19904 13970 19916
rect 14458 19904 14464 19916
rect 13964 19876 14464 19904
rect 13964 19864 13970 19876
rect 14458 19864 14464 19876
rect 14516 19864 14522 19916
rect 19242 19913 19248 19916
rect 19220 19907 19248 19913
rect 19220 19873 19232 19907
rect 19220 19867 19248 19873
rect 19242 19864 19248 19867
rect 19300 19864 19306 19916
rect 9171 19808 10640 19836
rect 9171 19805 9183 19808
rect 9125 19799 9183 19805
rect 12434 19796 12440 19848
rect 12492 19836 12498 19848
rect 12897 19839 12955 19845
rect 12897 19836 12909 19839
rect 12492 19808 12909 19836
rect 12492 19796 12498 19808
rect 12897 19805 12909 19808
rect 12943 19805 12955 19839
rect 16114 19836 16120 19848
rect 16075 19808 16120 19836
rect 12897 19799 12955 19805
rect 16114 19796 16120 19808
rect 16172 19796 16178 19848
rect 17678 19836 17684 19848
rect 17639 19808 17684 19836
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 17770 19796 17776 19848
rect 17828 19836 17834 19848
rect 17957 19839 18015 19845
rect 17957 19836 17969 19839
rect 17828 19808 17969 19836
rect 17828 19796 17834 19808
rect 17957 19805 17969 19808
rect 18003 19805 18015 19839
rect 17957 19799 18015 19805
rect 16666 19768 16672 19780
rect 16627 19740 16672 19768
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 1535 19703 1593 19709
rect 1535 19669 1547 19703
rect 1581 19700 1593 19703
rect 2590 19700 2596 19712
rect 1581 19672 2596 19700
rect 1581 19669 1593 19672
rect 1535 19663 1593 19669
rect 2590 19660 2596 19672
rect 2648 19660 2654 19712
rect 3145 19703 3203 19709
rect 3145 19669 3157 19703
rect 3191 19700 3203 19703
rect 3510 19700 3516 19712
rect 3191 19672 3516 19700
rect 3191 19669 3203 19672
rect 3145 19663 3203 19669
rect 3510 19660 3516 19672
rect 3568 19660 3574 19712
rect 7742 19700 7748 19712
rect 7703 19672 7748 19700
rect 7742 19660 7748 19672
rect 7800 19660 7806 19712
rect 12526 19700 12532 19712
rect 12487 19672 12532 19700
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 17954 19660 17960 19712
rect 18012 19700 18018 19712
rect 19291 19703 19349 19709
rect 19291 19700 19303 19703
rect 18012 19672 19303 19700
rect 18012 19660 18018 19672
rect 19291 19669 19303 19672
rect 19337 19669 19349 19703
rect 19291 19663 19349 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2501 19499 2559 19505
rect 2501 19465 2513 19499
rect 2547 19496 2559 19499
rect 3050 19496 3056 19508
rect 2547 19468 3056 19496
rect 2547 19465 2559 19468
rect 2501 19459 2559 19465
rect 3050 19456 3056 19468
rect 3108 19456 3114 19508
rect 4614 19456 4620 19508
rect 4672 19496 4678 19508
rect 4709 19499 4767 19505
rect 4709 19496 4721 19499
rect 4672 19468 4721 19496
rect 4672 19456 4678 19468
rect 4709 19465 4721 19468
rect 4755 19496 4767 19499
rect 5074 19496 5080 19508
rect 4755 19468 5080 19496
rect 4755 19465 4767 19468
rect 4709 19459 4767 19465
rect 5074 19456 5080 19468
rect 5132 19456 5138 19508
rect 10042 19456 10048 19508
rect 10100 19496 10106 19508
rect 10413 19499 10471 19505
rect 10413 19496 10425 19499
rect 10100 19468 10425 19496
rect 10100 19456 10106 19468
rect 10413 19465 10425 19468
rect 10459 19465 10471 19499
rect 10413 19459 10471 19465
rect 15841 19499 15899 19505
rect 15841 19465 15853 19499
rect 15887 19496 15899 19499
rect 16206 19496 16212 19508
rect 15887 19468 16212 19496
rect 15887 19465 15899 19468
rect 15841 19459 15899 19465
rect 16206 19456 16212 19468
rect 16264 19456 16270 19508
rect 17681 19499 17739 19505
rect 17681 19465 17693 19499
rect 17727 19496 17739 19499
rect 17862 19496 17868 19508
rect 17727 19468 17868 19496
rect 17727 19465 17739 19468
rect 17681 19459 17739 19465
rect 17862 19456 17868 19468
rect 17920 19456 17926 19508
rect 24762 19496 24768 19508
rect 24723 19468 24768 19496
rect 24762 19456 24768 19468
rect 24820 19456 24826 19508
rect 9674 19388 9680 19440
rect 9732 19428 9738 19440
rect 10689 19431 10747 19437
rect 10689 19428 10701 19431
rect 9732 19400 10701 19428
rect 9732 19388 9738 19400
rect 10689 19397 10701 19400
rect 10735 19397 10747 19431
rect 14734 19428 14740 19440
rect 10689 19391 10747 19397
rect 14292 19400 14740 19428
rect 2314 19320 2320 19372
rect 2372 19360 2378 19372
rect 2731 19363 2789 19369
rect 2731 19360 2743 19363
rect 2372 19332 2743 19360
rect 2372 19320 2378 19332
rect 2731 19329 2743 19332
rect 2777 19329 2789 19363
rect 2731 19323 2789 19329
rect 5905 19363 5963 19369
rect 5905 19329 5917 19363
rect 5951 19360 5963 19363
rect 6178 19360 6184 19372
rect 5951 19332 6184 19360
rect 5951 19329 5963 19332
rect 5905 19323 5963 19329
rect 6178 19320 6184 19332
rect 6236 19360 6242 19372
rect 9033 19363 9091 19369
rect 6236 19332 6408 19360
rect 6236 19320 6242 19332
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 2644 19295 2702 19301
rect 1443 19264 2084 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 2056 19165 2084 19264
rect 2644 19261 2656 19295
rect 2690 19292 2702 19295
rect 3513 19295 3571 19301
rect 2690 19264 3096 19292
rect 2690 19261 2702 19264
rect 2644 19255 2702 19261
rect 2041 19159 2099 19165
rect 2041 19125 2053 19159
rect 2087 19156 2099 19159
rect 2130 19156 2136 19168
rect 2087 19128 2136 19156
rect 2087 19125 2099 19128
rect 2041 19119 2099 19125
rect 2130 19116 2136 19128
rect 2188 19116 2194 19168
rect 3068 19165 3096 19264
rect 3513 19261 3525 19295
rect 3559 19292 3571 19295
rect 3602 19292 3608 19304
rect 3559 19264 3608 19292
rect 3559 19261 3571 19264
rect 3513 19255 3571 19261
rect 3602 19252 3608 19264
rect 3660 19252 3666 19304
rect 4157 19295 4215 19301
rect 4157 19261 4169 19295
rect 4203 19261 4215 19295
rect 4157 19255 4215 19261
rect 5077 19295 5135 19301
rect 5077 19261 5089 19295
rect 5123 19292 5135 19295
rect 5166 19292 5172 19304
rect 5123 19264 5172 19292
rect 5123 19261 5135 19264
rect 5077 19255 5135 19261
rect 4172 19224 4200 19255
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 5258 19252 5264 19304
rect 5316 19292 5322 19304
rect 5629 19295 5687 19301
rect 5629 19292 5641 19295
rect 5316 19264 5641 19292
rect 5316 19252 5322 19264
rect 5629 19261 5641 19264
rect 5675 19292 5687 19295
rect 5810 19292 5816 19304
rect 5675 19264 5816 19292
rect 5675 19261 5687 19264
rect 5629 19255 5687 19261
rect 5810 19252 5816 19264
rect 5868 19252 5874 19304
rect 6380 19292 6408 19332
rect 9033 19329 9045 19363
rect 9079 19360 9091 19363
rect 9398 19360 9404 19372
rect 9079 19332 9404 19360
rect 9079 19329 9091 19332
rect 9033 19323 9091 19329
rect 9398 19320 9404 19332
rect 9456 19320 9462 19372
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 14292 19360 14320 19400
rect 14734 19388 14740 19400
rect 14792 19388 14798 19440
rect 14366 19360 14372 19372
rect 12492 19332 13768 19360
rect 14292 19332 14372 19360
rect 12492 19320 12498 19332
rect 7009 19295 7067 19301
rect 7009 19292 7021 19295
rect 6380 19264 7021 19292
rect 7009 19261 7021 19264
rect 7055 19261 7067 19295
rect 7742 19292 7748 19304
rect 7703 19264 7748 19292
rect 7009 19255 7067 19261
rect 7742 19252 7748 19264
rect 7800 19252 7806 19304
rect 8662 19292 8668 19304
rect 8575 19264 8668 19292
rect 8662 19252 8668 19264
rect 8720 19252 8726 19304
rect 9490 19292 9496 19304
rect 9451 19264 9496 19292
rect 9490 19252 9496 19264
rect 9548 19252 9554 19304
rect 11333 19295 11391 19301
rect 11333 19292 11345 19295
rect 11164 19264 11345 19292
rect 5276 19224 5304 19252
rect 8066 19227 8124 19233
rect 8066 19224 8078 19227
rect 4172 19196 5304 19224
rect 7576 19196 8078 19224
rect 3053 19159 3111 19165
rect 3053 19125 3065 19159
rect 3099 19156 3111 19159
rect 3234 19156 3240 19168
rect 3099 19128 3240 19156
rect 3099 19125 3111 19128
rect 3053 19119 3111 19125
rect 3234 19116 3240 19128
rect 3292 19116 3298 19168
rect 3878 19156 3884 19168
rect 3839 19128 3884 19156
rect 3878 19116 3884 19128
rect 3936 19116 3942 19168
rect 6178 19116 6184 19168
rect 6236 19156 6242 19168
rect 6365 19159 6423 19165
rect 6365 19156 6377 19159
rect 6236 19128 6377 19156
rect 6236 19116 6242 19128
rect 6365 19125 6377 19128
rect 6411 19156 6423 19159
rect 6638 19156 6644 19168
rect 6411 19128 6644 19156
rect 6411 19125 6423 19128
rect 6365 19119 6423 19125
rect 6638 19116 6644 19128
rect 6696 19156 6702 19168
rect 7576 19165 7604 19196
rect 8066 19193 8078 19196
rect 8112 19193 8124 19227
rect 8680 19224 8708 19252
rect 9855 19227 9913 19233
rect 8680 19196 9444 19224
rect 8066 19187 8124 19193
rect 7561 19159 7619 19165
rect 7561 19156 7573 19159
rect 6696 19128 7573 19156
rect 6696 19116 6702 19128
rect 7561 19125 7573 19128
rect 7607 19125 7619 19159
rect 9306 19156 9312 19168
rect 9267 19128 9312 19156
rect 7561 19119 7619 19125
rect 9306 19116 9312 19128
rect 9364 19116 9370 19168
rect 9416 19156 9444 19196
rect 9855 19193 9867 19227
rect 9901 19224 9913 19227
rect 9950 19224 9956 19236
rect 9901 19196 9956 19224
rect 9901 19193 9913 19196
rect 9855 19187 9913 19193
rect 9950 19184 9956 19196
rect 10008 19184 10014 19236
rect 11164 19168 11192 19264
rect 11333 19261 11345 19264
rect 11379 19261 11391 19295
rect 12526 19292 12532 19304
rect 12487 19264 12532 19292
rect 11333 19255 11391 19261
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 13449 19295 13507 19301
rect 13449 19261 13461 19295
rect 13495 19292 13507 19295
rect 13630 19292 13636 19304
rect 13495 19264 13636 19292
rect 13495 19261 13507 19264
rect 13449 19255 13507 19261
rect 13630 19252 13636 19264
rect 13688 19252 13694 19304
rect 13740 19292 13768 19332
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 16114 19320 16120 19372
rect 16172 19360 16178 19372
rect 16485 19363 16543 19369
rect 16485 19360 16497 19363
rect 16172 19332 16497 19360
rect 16172 19320 16178 19332
rect 16485 19329 16497 19332
rect 16531 19360 16543 19363
rect 16531 19332 16896 19360
rect 16531 19329 16543 19332
rect 16485 19323 16543 19329
rect 14093 19295 14151 19301
rect 14093 19292 14105 19295
rect 13740 19264 14105 19292
rect 14093 19261 14105 19264
rect 14139 19261 14151 19295
rect 14093 19255 14151 19261
rect 14734 19252 14740 19304
rect 14792 19292 14798 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14792 19264 14933 19292
rect 14792 19252 14798 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 16704 19295 16762 19301
rect 16704 19292 16716 19295
rect 14921 19255 14979 19261
rect 16684 19261 16716 19292
rect 16750 19261 16762 19295
rect 16868 19292 16896 19332
rect 18322 19320 18328 19372
rect 18380 19360 18386 19372
rect 19242 19360 19248 19372
rect 18380 19332 19248 19360
rect 18380 19320 18386 19332
rect 19242 19320 19248 19332
rect 19300 19320 19306 19372
rect 17770 19292 17776 19304
rect 16868 19264 17776 19292
rect 16684 19255 16762 19261
rect 12891 19227 12949 19233
rect 12891 19193 12903 19227
rect 12937 19224 12949 19227
rect 15242 19227 15300 19233
rect 12937 19196 12971 19224
rect 12937 19193 12949 19196
rect 12891 19187 12949 19193
rect 15242 19193 15254 19227
rect 15288 19193 15300 19227
rect 15242 19187 15300 19193
rect 10134 19156 10140 19168
rect 9416 19128 10140 19156
rect 10134 19116 10140 19128
rect 10192 19116 10198 19168
rect 11146 19156 11152 19168
rect 11107 19128 11152 19156
rect 11146 19116 11152 19128
rect 11204 19116 11210 19168
rect 11422 19116 11428 19168
rect 11480 19156 11486 19168
rect 11517 19159 11575 19165
rect 11517 19156 11529 19159
rect 11480 19128 11529 19156
rect 11480 19116 11486 19128
rect 11517 19125 11529 19128
rect 11563 19125 11575 19159
rect 11517 19119 11575 19125
rect 11885 19159 11943 19165
rect 11885 19125 11897 19159
rect 11931 19156 11943 19159
rect 11974 19156 11980 19168
rect 11931 19128 11980 19156
rect 11931 19125 11943 19128
rect 11885 19119 11943 19125
rect 11974 19116 11980 19128
rect 12032 19116 12038 19168
rect 12253 19159 12311 19165
rect 12253 19125 12265 19159
rect 12299 19156 12311 19159
rect 12906 19156 12934 19187
rect 13446 19156 13452 19168
rect 12299 19128 13452 19156
rect 12299 19125 12311 19128
rect 12253 19119 12311 19125
rect 13446 19116 13452 19128
rect 13504 19156 13510 19168
rect 13725 19159 13783 19165
rect 13725 19156 13737 19159
rect 13504 19128 13737 19156
rect 13504 19116 13510 19128
rect 13725 19125 13737 19128
rect 13771 19156 13783 19159
rect 14737 19159 14795 19165
rect 14737 19156 14749 19159
rect 13771 19128 14749 19156
rect 13771 19125 13783 19128
rect 13725 19119 13783 19125
rect 14737 19125 14749 19128
rect 14783 19156 14795 19159
rect 15257 19156 15285 19187
rect 14783 19128 15285 19156
rect 16684 19156 16712 19255
rect 17770 19252 17776 19264
rect 17828 19252 17834 19304
rect 18046 19252 18052 19304
rect 18104 19301 18110 19304
rect 18104 19295 18142 19301
rect 18130 19292 18142 19295
rect 18509 19295 18567 19301
rect 18509 19292 18521 19295
rect 18130 19264 18521 19292
rect 18130 19261 18142 19264
rect 18104 19255 18142 19261
rect 18509 19261 18521 19264
rect 18555 19261 18567 19295
rect 19058 19292 19064 19304
rect 19019 19264 19064 19292
rect 18509 19255 18567 19261
rect 18104 19252 18110 19255
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 19260 19292 19288 19320
rect 19521 19295 19579 19301
rect 19521 19292 19533 19295
rect 19260 19264 19533 19292
rect 19521 19261 19533 19264
rect 19567 19261 19579 19295
rect 19886 19292 19892 19304
rect 19847 19264 19892 19292
rect 19521 19255 19579 19261
rect 19886 19252 19892 19264
rect 19944 19252 19950 19304
rect 24578 19292 24584 19304
rect 24539 19264 24584 19292
rect 24578 19252 24584 19264
rect 24636 19292 24642 19304
rect 25133 19295 25191 19301
rect 25133 19292 25145 19295
rect 24636 19264 25145 19292
rect 24636 19252 24642 19264
rect 25133 19261 25145 19264
rect 25179 19261 25191 19295
rect 25133 19255 25191 19261
rect 16807 19227 16865 19233
rect 16807 19193 16819 19227
rect 16853 19224 16865 19227
rect 17678 19224 17684 19236
rect 16853 19196 17684 19224
rect 16853 19193 16865 19196
rect 16807 19187 16865 19193
rect 17678 19184 17684 19196
rect 17736 19184 17742 19236
rect 19334 19184 19340 19236
rect 19392 19224 19398 19236
rect 20073 19227 20131 19233
rect 20073 19224 20085 19227
rect 19392 19196 20085 19224
rect 19392 19184 19398 19196
rect 20073 19193 20085 19196
rect 20119 19193 20131 19227
rect 20073 19187 20131 19193
rect 17218 19156 17224 19168
rect 16684 19128 17224 19156
rect 14783 19125 14795 19128
rect 14737 19119 14795 19125
rect 17218 19116 17224 19128
rect 17276 19116 17282 19168
rect 17954 19116 17960 19168
rect 18012 19156 18018 19168
rect 18187 19159 18245 19165
rect 18187 19156 18199 19159
rect 18012 19128 18199 19156
rect 18012 19116 18018 19128
rect 18187 19125 18199 19128
rect 18233 19125 18245 19159
rect 19242 19156 19248 19168
rect 19203 19128 19248 19156
rect 18187 19119 18245 19125
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 3697 18955 3755 18961
rect 3697 18921 3709 18955
rect 3743 18952 3755 18955
rect 4154 18952 4160 18964
rect 3743 18924 4160 18952
rect 3743 18921 3755 18924
rect 3697 18915 3755 18921
rect 4154 18912 4160 18924
rect 4212 18952 4218 18964
rect 4893 18955 4951 18961
rect 4893 18952 4905 18955
rect 4212 18924 4905 18952
rect 4212 18912 4218 18924
rect 4893 18921 4905 18924
rect 4939 18952 4951 18955
rect 5258 18952 5264 18964
rect 4939 18924 5264 18952
rect 4939 18921 4951 18924
rect 4893 18915 4951 18921
rect 5258 18912 5264 18924
rect 5316 18912 5322 18964
rect 9490 18952 9496 18964
rect 9451 18924 9496 18952
rect 9490 18912 9496 18924
rect 9548 18912 9554 18964
rect 11238 18952 11244 18964
rect 10244 18924 11244 18952
rect 6086 18884 6092 18896
rect 6047 18856 6092 18884
rect 6086 18844 6092 18856
rect 6144 18844 6150 18896
rect 8938 18844 8944 18896
rect 8996 18884 9002 18896
rect 9306 18884 9312 18896
rect 8996 18856 9312 18884
rect 8996 18844 9002 18856
rect 9306 18844 9312 18856
rect 9364 18884 9370 18896
rect 9950 18884 9956 18896
rect 9364 18856 9956 18884
rect 9364 18844 9370 18856
rect 9950 18844 9956 18856
rect 10008 18844 10014 18896
rect 10244 18893 10272 18924
rect 11238 18912 11244 18924
rect 11296 18912 11302 18964
rect 12529 18955 12587 18961
rect 12529 18921 12541 18955
rect 12575 18952 12587 18955
rect 12618 18952 12624 18964
rect 12575 18924 12624 18952
rect 12575 18921 12587 18924
rect 12529 18915 12587 18921
rect 12618 18912 12624 18924
rect 12676 18952 12682 18964
rect 14001 18955 14059 18961
rect 14001 18952 14013 18955
rect 12676 18924 14013 18952
rect 12676 18912 12682 18924
rect 14001 18921 14013 18924
rect 14047 18921 14059 18955
rect 14001 18915 14059 18921
rect 16209 18955 16267 18961
rect 16209 18921 16221 18955
rect 16255 18952 16267 18955
rect 16482 18952 16488 18964
rect 16255 18924 16488 18952
rect 16255 18921 16267 18924
rect 16209 18915 16267 18921
rect 16482 18912 16488 18924
rect 16540 18912 16546 18964
rect 17126 18952 17132 18964
rect 17087 18924 17132 18952
rect 17126 18912 17132 18924
rect 17184 18912 17190 18964
rect 17678 18912 17684 18964
rect 17736 18952 17742 18964
rect 18049 18955 18107 18961
rect 18049 18952 18061 18955
rect 17736 18924 18061 18952
rect 17736 18912 17742 18924
rect 18049 18921 18061 18924
rect 18095 18921 18107 18955
rect 18049 18915 18107 18921
rect 24670 18912 24676 18964
rect 24728 18952 24734 18964
rect 24765 18955 24823 18961
rect 24765 18952 24777 18955
rect 24728 18924 24777 18952
rect 24728 18912 24734 18924
rect 24765 18921 24777 18924
rect 24811 18921 24823 18955
rect 24765 18915 24823 18921
rect 10229 18887 10287 18893
rect 10229 18853 10241 18887
rect 10275 18853 10287 18887
rect 10229 18847 10287 18853
rect 10318 18844 10324 18896
rect 10376 18884 10382 18896
rect 10870 18884 10876 18896
rect 10376 18856 10421 18884
rect 10831 18856 10876 18884
rect 10376 18844 10382 18856
rect 10870 18844 10876 18856
rect 10928 18844 10934 18896
rect 13167 18887 13225 18893
rect 13167 18853 13179 18887
rect 13213 18884 13225 18887
rect 13446 18884 13452 18896
rect 13213 18856 13452 18884
rect 13213 18853 13225 18856
rect 13167 18847 13225 18853
rect 13446 18844 13452 18856
rect 13504 18844 13510 18896
rect 15562 18844 15568 18896
rect 15620 18893 15626 18896
rect 15620 18887 15668 18893
rect 15620 18853 15622 18887
rect 15656 18853 15668 18887
rect 15620 18847 15668 18853
rect 15620 18844 15626 18847
rect 16022 18844 16028 18896
rect 16080 18884 16086 18896
rect 16577 18887 16635 18893
rect 16577 18884 16589 18887
rect 16080 18856 16589 18884
rect 16080 18844 16086 18856
rect 16577 18853 16589 18856
rect 16623 18884 16635 18887
rect 17862 18884 17868 18896
rect 16623 18856 17868 18884
rect 16623 18853 16635 18856
rect 16577 18847 16635 18853
rect 17862 18844 17868 18856
rect 17920 18844 17926 18896
rect 2016 18819 2074 18825
rect 2016 18785 2028 18819
rect 2062 18816 2074 18819
rect 2222 18816 2228 18828
rect 2062 18788 2228 18816
rect 2062 18785 2074 18788
rect 2016 18779 2074 18785
rect 2222 18776 2228 18788
rect 2280 18816 2286 18828
rect 3028 18819 3086 18825
rect 3028 18816 3040 18819
rect 2280 18788 3040 18816
rect 2280 18776 2286 18788
rect 3028 18785 3040 18788
rect 3074 18816 3086 18819
rect 3142 18816 3148 18828
rect 3074 18788 3148 18816
rect 3074 18785 3086 18788
rect 3028 18779 3086 18785
rect 3142 18776 3148 18788
rect 3200 18776 3206 18828
rect 5445 18819 5503 18825
rect 5445 18785 5457 18819
rect 5491 18785 5503 18819
rect 5445 18779 5503 18785
rect 2682 18748 2688 18760
rect 2240 18720 2688 18748
rect 2240 18692 2268 18720
rect 2682 18708 2688 18720
rect 2740 18708 2746 18760
rect 3878 18708 3884 18760
rect 3936 18748 3942 18760
rect 4065 18751 4123 18757
rect 4065 18748 4077 18751
rect 3936 18720 4077 18748
rect 3936 18708 3942 18720
rect 4065 18717 4077 18720
rect 4111 18717 4123 18751
rect 5460 18748 5488 18779
rect 5534 18776 5540 18828
rect 5592 18816 5598 18828
rect 5810 18816 5816 18828
rect 5592 18788 5816 18816
rect 5592 18776 5598 18788
rect 5810 18776 5816 18788
rect 5868 18776 5874 18828
rect 7006 18816 7012 18828
rect 6967 18788 7012 18816
rect 7006 18776 7012 18788
rect 7064 18776 7070 18828
rect 7469 18819 7527 18825
rect 7469 18785 7481 18819
rect 7515 18816 7527 18819
rect 7742 18816 7748 18828
rect 7515 18788 7748 18816
rect 7515 18785 7527 18788
rect 7469 18779 7527 18785
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 8662 18825 8668 18828
rect 8640 18819 8668 18825
rect 8640 18785 8652 18819
rect 8640 18779 8668 18785
rect 8662 18776 8668 18779
rect 8720 18776 8726 18828
rect 11790 18825 11796 18828
rect 11768 18819 11796 18825
rect 11768 18785 11780 18819
rect 11768 18779 11796 18785
rect 11790 18776 11796 18779
rect 11848 18776 11854 18828
rect 13538 18776 13544 18828
rect 13596 18816 13602 18828
rect 13725 18819 13783 18825
rect 13725 18816 13737 18819
rect 13596 18788 13737 18816
rect 13596 18776 13602 18788
rect 13725 18785 13737 18788
rect 13771 18785 13783 18819
rect 17034 18816 17040 18828
rect 16995 18788 17040 18816
rect 13725 18779 13783 18785
rect 17034 18776 17040 18788
rect 17092 18776 17098 18828
rect 17589 18819 17647 18825
rect 17589 18785 17601 18819
rect 17635 18816 17647 18819
rect 17770 18816 17776 18828
rect 17635 18788 17776 18816
rect 17635 18785 17647 18788
rect 17589 18779 17647 18785
rect 17770 18776 17776 18788
rect 17828 18776 17834 18828
rect 18690 18825 18696 18828
rect 18668 18819 18696 18825
rect 18668 18785 18680 18819
rect 18668 18779 18696 18785
rect 18690 18776 18696 18779
rect 18748 18776 18754 18828
rect 19648 18819 19706 18825
rect 19648 18816 19660 18819
rect 18800 18788 19660 18816
rect 6362 18748 6368 18760
rect 5460 18720 6368 18748
rect 4065 18711 4123 18717
rect 6362 18708 6368 18720
rect 6420 18708 6426 18760
rect 7653 18751 7711 18757
rect 7653 18717 7665 18751
rect 7699 18748 7711 18751
rect 8018 18748 8024 18760
rect 7699 18720 8024 18748
rect 7699 18717 7711 18720
rect 7653 18711 7711 18717
rect 8018 18708 8024 18720
rect 8076 18708 8082 18760
rect 12805 18751 12863 18757
rect 12805 18717 12817 18751
rect 12851 18748 12863 18751
rect 13170 18748 13176 18760
rect 12851 18720 13176 18748
rect 12851 18717 12863 18720
rect 12805 18711 12863 18717
rect 13170 18708 13176 18720
rect 13228 18708 13234 18760
rect 15286 18748 15292 18760
rect 15247 18720 15292 18748
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 18046 18708 18052 18760
rect 18104 18748 18110 18760
rect 18800 18748 18828 18788
rect 19648 18785 19660 18788
rect 19694 18816 19706 18819
rect 20070 18816 20076 18828
rect 19694 18788 20076 18816
rect 19694 18785 19706 18788
rect 19648 18779 19706 18785
rect 20070 18776 20076 18788
rect 20128 18776 20134 18828
rect 24581 18819 24639 18825
rect 24581 18785 24593 18819
rect 24627 18816 24639 18819
rect 24670 18816 24676 18828
rect 24627 18788 24676 18816
rect 24627 18785 24639 18788
rect 24581 18779 24639 18785
rect 24670 18776 24676 18788
rect 24728 18776 24734 18828
rect 20898 18748 20904 18760
rect 18104 18720 18828 18748
rect 20859 18720 20904 18748
rect 18104 18708 18110 18720
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 2222 18640 2228 18692
rect 2280 18640 2286 18692
rect 4890 18640 4896 18692
rect 4948 18680 4954 18692
rect 9030 18680 9036 18692
rect 4948 18652 9036 18680
rect 4948 18640 4954 18652
rect 9030 18640 9036 18652
rect 9088 18640 9094 18692
rect 1673 18615 1731 18621
rect 1673 18581 1685 18615
rect 1719 18612 1731 18615
rect 1854 18612 1860 18624
rect 1719 18584 1860 18612
rect 1719 18581 1731 18584
rect 1673 18575 1731 18581
rect 1854 18572 1860 18584
rect 1912 18572 1918 18624
rect 2087 18615 2145 18621
rect 2087 18581 2099 18615
rect 2133 18612 2145 18615
rect 2682 18612 2688 18624
rect 2133 18584 2688 18612
rect 2133 18581 2145 18584
rect 2087 18575 2145 18581
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 3099 18615 3157 18621
rect 3099 18581 3111 18615
rect 3145 18612 3157 18615
rect 3418 18612 3424 18624
rect 3145 18584 3424 18612
rect 3145 18581 3157 18584
rect 3099 18575 3157 18581
rect 3418 18572 3424 18584
rect 3476 18572 3482 18624
rect 5258 18612 5264 18624
rect 5219 18584 5264 18612
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 8021 18615 8079 18621
rect 8021 18581 8033 18615
rect 8067 18612 8079 18615
rect 8110 18612 8116 18624
rect 8067 18584 8116 18612
rect 8067 18581 8079 18584
rect 8021 18575 8079 18581
rect 8110 18572 8116 18584
rect 8168 18572 8174 18624
rect 8711 18615 8769 18621
rect 8711 18581 8723 18615
rect 8757 18612 8769 18615
rect 9582 18612 9588 18624
rect 8757 18584 9588 18612
rect 8757 18581 8769 18584
rect 8711 18575 8769 18581
rect 9582 18572 9588 18584
rect 9640 18572 9646 18624
rect 11839 18615 11897 18621
rect 11839 18581 11851 18615
rect 11885 18612 11897 18615
rect 12066 18612 12072 18624
rect 11885 18584 12072 18612
rect 11885 18581 11897 18584
rect 11839 18575 11897 18581
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 14734 18572 14740 18624
rect 14792 18612 14798 18624
rect 14921 18615 14979 18621
rect 14921 18612 14933 18615
rect 14792 18584 14933 18612
rect 14792 18572 14798 18584
rect 14921 18581 14933 18584
rect 14967 18581 14979 18615
rect 14921 18575 14979 18581
rect 18598 18572 18604 18624
rect 18656 18612 18662 18624
rect 18739 18615 18797 18621
rect 18739 18612 18751 18615
rect 18656 18584 18751 18612
rect 18656 18572 18662 18584
rect 18739 18581 18751 18584
rect 18785 18581 18797 18615
rect 18739 18575 18797 18581
rect 19751 18615 19809 18621
rect 19751 18581 19763 18615
rect 19797 18612 19809 18615
rect 20346 18612 20352 18624
rect 19797 18584 20352 18612
rect 19797 18581 19809 18584
rect 19751 18575 19809 18581
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2498 18408 2504 18420
rect 2459 18380 2504 18408
rect 2498 18368 2504 18380
rect 2556 18368 2562 18420
rect 7006 18408 7012 18420
rect 6967 18380 7012 18408
rect 7006 18368 7012 18380
rect 7064 18368 7070 18420
rect 9030 18408 9036 18420
rect 8991 18380 9036 18408
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 11514 18368 11520 18420
rect 11572 18408 11578 18420
rect 11790 18408 11796 18420
rect 11572 18380 11796 18408
rect 11572 18368 11578 18380
rect 11790 18368 11796 18380
rect 11848 18368 11854 18420
rect 15838 18408 15844 18420
rect 15799 18380 15844 18408
rect 15838 18368 15844 18380
rect 15896 18368 15902 18420
rect 20070 18408 20076 18420
rect 20031 18380 20076 18408
rect 20070 18368 20076 18380
rect 20128 18368 20134 18420
rect 1648 18207 1706 18213
rect 1648 18173 1660 18207
rect 1694 18204 1706 18207
rect 2516 18204 2544 18368
rect 6641 18343 6699 18349
rect 6641 18340 6653 18343
rect 3896 18312 6653 18340
rect 3142 18204 3148 18216
rect 1694 18176 2544 18204
rect 2675 18176 3148 18204
rect 1694 18173 1706 18176
rect 1648 18167 1706 18173
rect 2133 18139 2191 18145
rect 2133 18105 2145 18139
rect 2179 18136 2191 18139
rect 2675 18136 2703 18176
rect 3142 18164 3148 18176
rect 3200 18164 3206 18216
rect 3896 18213 3924 18312
rect 6641 18309 6653 18312
rect 6687 18340 6699 18343
rect 7098 18340 7104 18352
rect 6687 18312 7104 18340
rect 6687 18309 6699 18312
rect 6641 18303 6699 18309
rect 7098 18300 7104 18312
rect 7156 18340 7162 18352
rect 7742 18340 7748 18352
rect 7156 18312 7748 18340
rect 7156 18300 7162 18312
rect 7742 18300 7748 18312
rect 7800 18300 7806 18352
rect 12250 18300 12256 18352
rect 12308 18340 12314 18352
rect 16574 18340 16580 18352
rect 12308 18312 12480 18340
rect 16535 18312 16580 18340
rect 12308 18300 12314 18312
rect 5258 18232 5264 18284
rect 5316 18272 5322 18284
rect 5316 18244 5764 18272
rect 5316 18232 5322 18244
rect 3513 18207 3571 18213
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 3881 18207 3939 18213
rect 3881 18204 3893 18207
rect 3559 18176 3893 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 3881 18173 3893 18176
rect 3927 18173 3939 18207
rect 4154 18204 4160 18216
rect 4115 18176 4160 18204
rect 3881 18167 3939 18173
rect 4154 18164 4160 18176
rect 4212 18164 4218 18216
rect 4706 18164 4712 18216
rect 4764 18204 4770 18216
rect 5077 18207 5135 18213
rect 5077 18204 5089 18207
rect 4764 18176 5089 18204
rect 4764 18164 4770 18176
rect 5077 18173 5089 18176
rect 5123 18204 5135 18207
rect 5350 18204 5356 18216
rect 5123 18176 5356 18204
rect 5123 18173 5135 18176
rect 5077 18167 5135 18173
rect 5350 18164 5356 18176
rect 5408 18164 5414 18216
rect 5736 18213 5764 18244
rect 6914 18232 6920 18284
rect 6972 18272 6978 18284
rect 8021 18275 8079 18281
rect 8021 18272 8033 18275
rect 6972 18244 8033 18272
rect 6972 18232 6978 18244
rect 8021 18241 8033 18244
rect 8067 18272 8079 18275
rect 8202 18272 8208 18284
rect 8067 18244 8208 18272
rect 8067 18241 8079 18244
rect 8021 18235 8079 18241
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 11422 18272 11428 18284
rect 10367 18244 11428 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 5721 18207 5779 18213
rect 5721 18173 5733 18207
rect 5767 18204 5779 18207
rect 6270 18204 6276 18216
rect 5767 18176 6276 18204
rect 5767 18173 5779 18176
rect 5721 18167 5779 18173
rect 6270 18164 6276 18176
rect 6328 18164 6334 18216
rect 8662 18204 8668 18216
rect 8623 18176 8668 18204
rect 8662 18164 8668 18176
rect 8720 18164 8726 18216
rect 9030 18164 9036 18216
rect 9088 18204 9094 18216
rect 9214 18204 9220 18216
rect 9088 18176 9220 18204
rect 9088 18164 9094 18176
rect 9214 18164 9220 18176
rect 9272 18164 9278 18216
rect 9766 18204 9772 18216
rect 9727 18176 9772 18204
rect 9766 18164 9772 18176
rect 9824 18164 9830 18216
rect 11256 18213 11284 18244
rect 11422 18232 11428 18244
rect 11480 18232 11486 18284
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 12342 18272 12348 18284
rect 11563 18244 12348 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 12452 18213 12480 18312
rect 16574 18300 16580 18312
rect 16632 18300 16638 18352
rect 24578 18340 24584 18352
rect 24539 18312 24584 18340
rect 24578 18300 24584 18312
rect 24636 18300 24642 18352
rect 14734 18272 14740 18284
rect 14695 18244 14740 18272
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 16022 18272 16028 18284
rect 15983 18244 16028 18272
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 18739 18275 18797 18281
rect 18739 18241 18751 18275
rect 18785 18272 18797 18275
rect 19242 18272 19248 18284
rect 18785 18244 19248 18272
rect 18785 18241 18797 18244
rect 18739 18235 18797 18241
rect 19242 18232 19248 18244
rect 19300 18232 19306 18284
rect 20441 18275 20499 18281
rect 20441 18272 20453 18275
rect 19663 18244 20453 18272
rect 19663 18216 19691 18244
rect 20441 18241 20453 18244
rect 20487 18272 20499 18275
rect 21910 18272 21916 18284
rect 20487 18244 21916 18272
rect 20487 18241 20499 18244
rect 20441 18235 20499 18241
rect 21910 18232 21916 18244
rect 21968 18232 21974 18284
rect 10965 18207 11023 18213
rect 10965 18173 10977 18207
rect 11011 18173 11023 18207
rect 10965 18167 11023 18173
rect 11241 18207 11299 18213
rect 11241 18173 11253 18207
rect 11287 18173 11299 18207
rect 11241 18167 11299 18173
rect 12437 18207 12495 18213
rect 12437 18173 12449 18207
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 12897 18207 12955 18213
rect 12897 18173 12909 18207
rect 12943 18173 12955 18207
rect 14001 18207 14059 18213
rect 14001 18204 14013 18207
rect 12897 18167 12955 18173
rect 13832 18176 14013 18204
rect 2179 18108 2703 18136
rect 5905 18139 5963 18145
rect 2179 18105 2191 18108
rect 2133 18099 2191 18105
rect 5905 18105 5917 18139
rect 5951 18136 5963 18139
rect 6638 18136 6644 18148
rect 5951 18108 6644 18136
rect 5951 18105 5963 18108
rect 5905 18099 5963 18105
rect 6638 18096 6644 18108
rect 6696 18096 6702 18148
rect 7377 18139 7435 18145
rect 7377 18105 7389 18139
rect 7423 18105 7435 18139
rect 7377 18099 7435 18105
rect 1762 18077 1768 18080
rect 1719 18071 1768 18077
rect 1719 18037 1731 18071
rect 1765 18037 1768 18071
rect 1719 18031 1768 18037
rect 1762 18028 1768 18031
rect 1820 18028 1826 18080
rect 2590 18068 2596 18080
rect 2551 18040 2596 18068
rect 2590 18028 2596 18040
rect 2648 18028 2654 18080
rect 3142 18028 3148 18080
rect 3200 18068 3206 18080
rect 3881 18071 3939 18077
rect 3200 18040 3245 18068
rect 3200 18028 3206 18040
rect 3881 18037 3893 18071
rect 3927 18068 3939 18071
rect 4062 18068 4068 18080
rect 3927 18040 4068 18068
rect 3927 18037 3939 18040
rect 3881 18031 3939 18037
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 6273 18071 6331 18077
rect 6273 18037 6285 18071
rect 6319 18068 6331 18071
rect 6362 18068 6368 18080
rect 6319 18040 6368 18068
rect 6319 18037 6331 18040
rect 6273 18031 6331 18037
rect 6362 18028 6368 18040
rect 6420 18028 6426 18080
rect 7392 18068 7420 18099
rect 7466 18096 7472 18148
rect 7524 18136 7530 18148
rect 9953 18139 10011 18145
rect 7524 18108 7569 18136
rect 7524 18096 7530 18108
rect 9953 18105 9965 18139
rect 9999 18136 10011 18139
rect 10870 18136 10876 18148
rect 9999 18108 10876 18136
rect 9999 18105 10011 18108
rect 9953 18099 10011 18105
rect 10870 18096 10876 18108
rect 10928 18096 10934 18148
rect 8110 18068 8116 18080
rect 7392 18040 8116 18068
rect 8110 18028 8116 18040
rect 8168 18028 8174 18080
rect 10042 18028 10048 18080
rect 10100 18068 10106 18080
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 10100 18040 10701 18068
rect 10100 18028 10106 18040
rect 10689 18037 10701 18040
rect 10735 18068 10747 18071
rect 10980 18068 11008 18167
rect 11256 18136 11284 18167
rect 12618 18136 12624 18148
rect 11256 18108 12624 18136
rect 12618 18096 12624 18108
rect 12676 18136 12682 18148
rect 12912 18136 12940 18167
rect 13170 18136 13176 18148
rect 12676 18108 12940 18136
rect 13131 18108 13176 18136
rect 12676 18096 12682 18108
rect 13170 18096 13176 18108
rect 13228 18096 13234 18148
rect 13832 18080 13860 18176
rect 14001 18173 14013 18176
rect 14047 18173 14059 18207
rect 14001 18167 14059 18173
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14461 18207 14519 18213
rect 14461 18204 14473 18207
rect 14240 18176 14473 18204
rect 14240 18164 14246 18176
rect 14461 18173 14473 18176
rect 14507 18173 14519 18207
rect 14461 18167 14519 18173
rect 18414 18164 18420 18216
rect 18472 18204 18478 18216
rect 18636 18207 18694 18213
rect 18636 18204 18648 18207
rect 18472 18176 18648 18204
rect 18472 18164 18478 18176
rect 18636 18173 18648 18176
rect 18682 18204 18694 18207
rect 19429 18207 19487 18213
rect 19429 18204 19441 18207
rect 18682 18176 19441 18204
rect 18682 18173 18694 18176
rect 18636 18167 18694 18173
rect 19429 18173 19441 18176
rect 19475 18173 19487 18207
rect 19645 18204 19651 18216
rect 19606 18176 19651 18204
rect 19429 18167 19487 18173
rect 19645 18164 19651 18176
rect 19703 18164 19709 18216
rect 15838 18096 15844 18148
rect 15896 18136 15902 18148
rect 16117 18139 16175 18145
rect 16117 18136 16129 18139
rect 15896 18108 16129 18136
rect 15896 18096 15902 18108
rect 16117 18105 16129 18108
rect 16163 18105 16175 18139
rect 16117 18099 16175 18105
rect 11698 18068 11704 18080
rect 10735 18040 11704 18068
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 12250 18068 12256 18080
rect 12211 18040 12256 18068
rect 12250 18028 12256 18040
rect 12308 18028 12314 18080
rect 13446 18068 13452 18080
rect 13407 18040 13452 18068
rect 13446 18028 13452 18040
rect 13504 18028 13510 18080
rect 13814 18068 13820 18080
rect 13775 18040 13820 18068
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 15289 18071 15347 18077
rect 15289 18068 15301 18071
rect 14792 18040 15301 18068
rect 14792 18028 14798 18040
rect 15289 18037 15301 18040
rect 15335 18068 15347 18071
rect 15562 18068 15568 18080
rect 15335 18040 15568 18068
rect 15335 18037 15347 18040
rect 15289 18031 15347 18037
rect 15562 18028 15568 18040
rect 15620 18028 15626 18080
rect 17034 18068 17040 18080
rect 16995 18040 17040 18068
rect 17034 18028 17040 18040
rect 17092 18028 17098 18080
rect 17497 18071 17555 18077
rect 17497 18037 17509 18071
rect 17543 18068 17555 18071
rect 17770 18068 17776 18080
rect 17543 18040 17776 18068
rect 17543 18037 17555 18040
rect 17497 18031 17555 18037
rect 17770 18028 17776 18040
rect 17828 18028 17834 18080
rect 18690 18028 18696 18080
rect 18748 18068 18754 18080
rect 19153 18071 19211 18077
rect 19153 18068 19165 18071
rect 18748 18040 19165 18068
rect 18748 18028 18754 18040
rect 19153 18037 19165 18040
rect 19199 18068 19211 18071
rect 19242 18068 19248 18080
rect 19199 18040 19248 18068
rect 19199 18037 19211 18040
rect 19153 18031 19211 18037
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 19751 18071 19809 18077
rect 19751 18037 19763 18071
rect 19797 18068 19809 18071
rect 20254 18068 20260 18080
rect 19797 18040 20260 18068
rect 19797 18037 19809 18040
rect 19751 18031 19809 18037
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 20622 18068 20628 18080
rect 20583 18040 20628 18068
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 21174 18028 21180 18080
rect 21232 18068 21238 18080
rect 21637 18071 21695 18077
rect 21637 18068 21649 18071
rect 21232 18040 21649 18068
rect 21232 18028 21238 18040
rect 21637 18037 21649 18040
rect 21683 18037 21695 18071
rect 21637 18031 21695 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 3697 17867 3755 17873
rect 3697 17833 3709 17867
rect 3743 17864 3755 17867
rect 4062 17864 4068 17876
rect 3743 17836 4068 17864
rect 3743 17833 3755 17836
rect 3697 17827 3755 17833
rect 4062 17824 4068 17836
rect 4120 17824 4126 17876
rect 5534 17864 5540 17876
rect 5495 17836 5540 17864
rect 5534 17824 5540 17836
rect 5592 17824 5598 17876
rect 6917 17867 6975 17873
rect 6917 17833 6929 17867
rect 6963 17864 6975 17867
rect 7377 17867 7435 17873
rect 7377 17864 7389 17867
rect 6963 17836 7389 17864
rect 6963 17833 6975 17836
rect 6917 17827 6975 17833
rect 7377 17833 7389 17836
rect 7423 17864 7435 17867
rect 7466 17864 7472 17876
rect 7423 17836 7472 17864
rect 7423 17833 7435 17836
rect 7377 17827 7435 17833
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 9309 17867 9367 17873
rect 9309 17833 9321 17867
rect 9355 17864 9367 17867
rect 9766 17864 9772 17876
rect 9355 17836 9772 17864
rect 9355 17833 9367 17836
rect 9309 17827 9367 17833
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 10134 17864 10140 17876
rect 10095 17836 10140 17864
rect 10134 17824 10140 17836
rect 10192 17824 10198 17876
rect 13081 17867 13139 17873
rect 13081 17833 13093 17867
rect 13127 17864 13139 17867
rect 13170 17864 13176 17876
rect 13127 17836 13176 17864
rect 13127 17833 13139 17836
rect 13081 17827 13139 17833
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 16114 17824 16120 17876
rect 16172 17864 16178 17876
rect 16485 17867 16543 17873
rect 16485 17864 16497 17867
rect 16172 17836 16497 17864
rect 16172 17824 16178 17836
rect 16485 17833 16497 17836
rect 16531 17864 16543 17867
rect 18417 17867 18475 17873
rect 18417 17864 18429 17867
rect 16531 17836 18429 17864
rect 16531 17833 16543 17836
rect 16485 17827 16543 17833
rect 18417 17833 18429 17836
rect 18463 17833 18475 17867
rect 18417 17827 18475 17833
rect 6178 17756 6184 17808
rect 6236 17796 6242 17808
rect 6318 17799 6376 17805
rect 6318 17796 6330 17799
rect 6236 17768 6330 17796
rect 6236 17756 6242 17768
rect 6318 17765 6330 17768
rect 6364 17765 6376 17799
rect 7926 17796 7932 17808
rect 7887 17768 7932 17796
rect 6318 17759 6376 17765
rect 7926 17756 7932 17768
rect 7984 17756 7990 17808
rect 8294 17756 8300 17808
rect 8352 17796 8358 17808
rect 8481 17799 8539 17805
rect 8481 17796 8493 17799
rect 8352 17768 8493 17796
rect 8352 17756 8358 17768
rect 8481 17765 8493 17768
rect 8527 17765 8539 17799
rect 8481 17759 8539 17765
rect 10597 17799 10655 17805
rect 10597 17765 10609 17799
rect 10643 17796 10655 17799
rect 10778 17796 10784 17808
rect 10643 17768 10784 17796
rect 10643 17765 10655 17768
rect 10597 17759 10655 17765
rect 10778 17756 10784 17768
rect 10836 17756 10842 17808
rect 14182 17796 14188 17808
rect 12636 17768 14188 17796
rect 12636 17740 12664 17768
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17728 2007 17731
rect 2130 17728 2136 17740
rect 1995 17700 2136 17728
rect 1995 17697 2007 17700
rect 1949 17691 2007 17697
rect 2130 17688 2136 17700
rect 2188 17688 2194 17740
rect 4706 17728 4712 17740
rect 4667 17700 4712 17728
rect 4706 17688 4712 17700
rect 4764 17688 4770 17740
rect 4985 17731 5043 17737
rect 4985 17697 4997 17731
rect 5031 17728 5043 17731
rect 5258 17728 5264 17740
rect 5031 17700 5264 17728
rect 5031 17697 5043 17700
rect 4985 17691 5043 17697
rect 5258 17688 5264 17700
rect 5316 17688 5322 17740
rect 11422 17688 11428 17740
rect 11480 17728 11486 17740
rect 11977 17731 12035 17737
rect 11977 17728 11989 17731
rect 11480 17700 11989 17728
rect 11480 17688 11486 17700
rect 11977 17697 11989 17700
rect 12023 17697 12035 17731
rect 11977 17691 12035 17697
rect 12437 17731 12495 17737
rect 12437 17697 12449 17731
rect 12483 17728 12495 17731
rect 12618 17728 12624 17740
rect 12483 17700 12624 17728
rect 12483 17697 12495 17700
rect 12437 17691 12495 17697
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 12894 17688 12900 17740
rect 12952 17728 12958 17740
rect 13538 17728 13544 17740
rect 12952 17700 13544 17728
rect 12952 17688 12958 17700
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 14016 17737 14044 17768
rect 14182 17756 14188 17768
rect 14240 17756 14246 17808
rect 14277 17799 14335 17805
rect 14277 17765 14289 17799
rect 14323 17796 14335 17799
rect 15286 17796 15292 17808
rect 14323 17768 15292 17796
rect 14323 17765 14335 17768
rect 14277 17759 14335 17765
rect 15286 17756 15292 17768
rect 15344 17796 15350 17808
rect 16942 17805 16948 17808
rect 16025 17799 16083 17805
rect 16025 17796 16037 17799
rect 15344 17768 16037 17796
rect 15344 17756 15350 17768
rect 16025 17765 16037 17768
rect 16071 17765 16083 17799
rect 16939 17796 16948 17805
rect 16903 17768 16948 17796
rect 16025 17759 16083 17765
rect 16939 17759 16948 17768
rect 16942 17756 16948 17759
rect 17000 17756 17006 17808
rect 17770 17756 17776 17808
rect 17828 17796 17834 17808
rect 17828 17768 18828 17796
rect 17828 17756 17834 17768
rect 14001 17731 14059 17737
rect 14001 17697 14013 17731
rect 14047 17697 14059 17731
rect 14001 17691 14059 17697
rect 15632 17731 15690 17737
rect 15632 17697 15644 17731
rect 15678 17728 15690 17731
rect 15746 17728 15752 17740
rect 15678 17700 15752 17728
rect 15678 17697 15690 17700
rect 15632 17691 15690 17697
rect 15746 17688 15752 17700
rect 15804 17688 15810 17740
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17728 16635 17731
rect 16666 17728 16672 17740
rect 16623 17700 16672 17728
rect 16623 17697 16635 17700
rect 16577 17691 16635 17697
rect 16666 17688 16672 17700
rect 16724 17728 16730 17740
rect 17126 17728 17132 17740
rect 16724 17700 17132 17728
rect 16724 17688 16730 17700
rect 17126 17688 17132 17700
rect 17184 17688 17190 17740
rect 18601 17731 18659 17737
rect 18601 17697 18613 17731
rect 18647 17728 18659 17731
rect 18690 17728 18696 17740
rect 18647 17700 18696 17728
rect 18647 17697 18659 17700
rect 18601 17691 18659 17697
rect 18690 17688 18696 17700
rect 18748 17688 18754 17740
rect 18800 17737 18828 17768
rect 18785 17731 18843 17737
rect 18785 17697 18797 17731
rect 18831 17697 18843 17731
rect 18785 17691 18843 17697
rect 20806 17688 20812 17740
rect 20864 17728 20870 17740
rect 20936 17731 20994 17737
rect 20936 17728 20948 17731
rect 20864 17700 20948 17728
rect 20864 17688 20870 17700
rect 20936 17697 20948 17700
rect 20982 17697 20994 17731
rect 20936 17691 20994 17697
rect 22256 17731 22314 17737
rect 22256 17697 22268 17731
rect 22302 17728 22314 17731
rect 22830 17728 22836 17740
rect 22302 17700 22836 17728
rect 22302 17697 22314 17700
rect 22256 17691 22314 17697
rect 22830 17688 22836 17700
rect 22888 17688 22894 17740
rect 23268 17731 23326 17737
rect 23268 17697 23280 17731
rect 23314 17728 23326 17731
rect 23382 17728 23388 17740
rect 23314 17700 23388 17728
rect 23314 17697 23326 17700
rect 23268 17691 23326 17697
rect 23382 17688 23388 17700
rect 23440 17688 23446 17740
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17660 3019 17663
rect 3234 17660 3240 17672
rect 3007 17632 3240 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 5169 17663 5227 17669
rect 5169 17629 5181 17663
rect 5215 17660 5227 17663
rect 5997 17663 6055 17669
rect 5997 17660 6009 17663
rect 5215 17632 6009 17660
rect 5215 17629 5227 17632
rect 5169 17623 5227 17629
rect 5997 17629 6009 17632
rect 6043 17660 6055 17663
rect 6822 17660 6828 17672
rect 6043 17632 6828 17660
rect 6043 17629 6055 17632
rect 5997 17623 6055 17629
rect 6822 17620 6828 17632
rect 6880 17620 6886 17672
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17660 7895 17663
rect 8662 17660 8668 17672
rect 7883 17632 8668 17660
rect 7883 17629 7895 17632
rect 7837 17623 7895 17629
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 10505 17663 10563 17669
rect 10505 17629 10517 17663
rect 10551 17660 10563 17663
rect 10962 17660 10968 17672
rect 10551 17632 10968 17660
rect 10551 17629 10563 17632
rect 10505 17623 10563 17629
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 12526 17660 12532 17672
rect 12487 17632 12532 17660
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 11054 17592 11060 17604
rect 11015 17564 11060 17592
rect 11054 17552 11060 17564
rect 11112 17592 11118 17604
rect 11698 17592 11704 17604
rect 11112 17564 11704 17592
rect 11112 17552 11118 17564
rect 11698 17552 11704 17564
rect 11756 17552 11762 17604
rect 1486 17484 1492 17536
rect 1544 17524 1550 17536
rect 2133 17527 2191 17533
rect 2133 17524 2145 17527
rect 1544 17496 2145 17524
rect 1544 17484 1550 17496
rect 2133 17493 2145 17496
rect 2179 17493 2191 17527
rect 2133 17487 2191 17493
rect 4341 17527 4399 17533
rect 4341 17493 4353 17527
rect 4387 17524 4399 17527
rect 4798 17524 4804 17536
rect 4387 17496 4804 17524
rect 4387 17493 4399 17496
rect 4341 17487 4399 17493
rect 4798 17484 4804 17496
rect 4856 17484 4862 17536
rect 14550 17524 14556 17536
rect 14511 17496 14556 17524
rect 14550 17484 14556 17496
rect 14608 17484 14614 17536
rect 15703 17527 15761 17533
rect 15703 17493 15715 17527
rect 15749 17524 15761 17527
rect 16482 17524 16488 17536
rect 15749 17496 16488 17524
rect 15749 17493 15761 17496
rect 15703 17487 15761 17493
rect 16482 17484 16488 17496
rect 16540 17484 16546 17536
rect 17494 17524 17500 17536
rect 17455 17496 17500 17524
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 18141 17527 18199 17533
rect 18141 17493 18153 17527
rect 18187 17524 18199 17527
rect 18230 17524 18236 17536
rect 18187 17496 18236 17524
rect 18187 17493 18199 17496
rect 18141 17487 18199 17493
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 21039 17527 21097 17533
rect 21039 17493 21051 17527
rect 21085 17524 21097 17527
rect 21358 17524 21364 17536
rect 21085 17496 21364 17524
rect 21085 17493 21097 17496
rect 21039 17487 21097 17493
rect 21358 17484 21364 17496
rect 21416 17484 21422 17536
rect 22370 17533 22376 17536
rect 22327 17527 22376 17533
rect 22327 17493 22339 17527
rect 22373 17493 22376 17527
rect 22327 17487 22376 17493
rect 22370 17484 22376 17487
rect 22428 17484 22434 17536
rect 22462 17484 22468 17536
rect 22520 17524 22526 17536
rect 23339 17527 23397 17533
rect 23339 17524 23351 17527
rect 22520 17496 23351 17524
rect 22520 17484 22526 17496
rect 23339 17493 23351 17496
rect 23385 17493 23397 17527
rect 23339 17487 23397 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 4525 17323 4583 17329
rect 4525 17289 4537 17323
rect 4571 17320 4583 17323
rect 4706 17320 4712 17332
rect 4571 17292 4712 17320
rect 4571 17289 4583 17292
rect 4525 17283 4583 17289
rect 4706 17280 4712 17292
rect 4764 17320 4770 17332
rect 5074 17320 5080 17332
rect 4764 17292 5080 17320
rect 4764 17280 4770 17292
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 5258 17280 5264 17332
rect 5316 17320 5322 17332
rect 5534 17320 5540 17332
rect 5316 17292 5540 17320
rect 5316 17280 5322 17292
rect 5534 17280 5540 17292
rect 5592 17320 5598 17332
rect 5721 17323 5779 17329
rect 5721 17320 5733 17323
rect 5592 17292 5733 17320
rect 5592 17280 5598 17292
rect 5721 17289 5733 17292
rect 5767 17320 5779 17323
rect 6362 17320 6368 17332
rect 5767 17292 6368 17320
rect 5767 17289 5779 17292
rect 5721 17283 5779 17289
rect 6362 17280 6368 17292
rect 6420 17280 6426 17332
rect 7745 17323 7803 17329
rect 7745 17289 7757 17323
rect 7791 17320 7803 17323
rect 7926 17320 7932 17332
rect 7791 17292 7932 17320
rect 7791 17289 7803 17292
rect 7745 17283 7803 17289
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 8018 17280 8024 17332
rect 8076 17320 8082 17332
rect 8076 17292 8121 17320
rect 8076 17280 8082 17292
rect 20806 17280 20812 17332
rect 20864 17320 20870 17332
rect 21085 17323 21143 17329
rect 21085 17320 21097 17323
rect 20864 17292 21097 17320
rect 20864 17280 20870 17292
rect 21085 17289 21097 17292
rect 21131 17289 21143 17323
rect 24762 17320 24768 17332
rect 24723 17292 24768 17320
rect 21085 17283 21143 17289
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 1578 17144 1584 17196
rect 1636 17184 1642 17196
rect 2038 17184 2044 17196
rect 1636 17156 2044 17184
rect 1636 17144 1642 17156
rect 2038 17144 2044 17156
rect 2096 17144 2102 17196
rect 3145 17187 3203 17193
rect 3145 17184 3157 17187
rect 2608 17156 3157 17184
rect 2608 17125 2636 17156
rect 3145 17153 3157 17156
rect 3191 17184 3203 17187
rect 3786 17184 3792 17196
rect 3191 17156 3792 17184
rect 3191 17153 3203 17156
rect 3145 17147 3203 17153
rect 3786 17144 3792 17156
rect 3844 17144 3850 17196
rect 4706 17184 4712 17196
rect 4667 17156 4712 17184
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 6638 17144 6644 17196
rect 6696 17184 6702 17196
rect 6825 17187 6883 17193
rect 6825 17184 6837 17187
rect 6696 17156 6837 17184
rect 6696 17144 6702 17156
rect 6825 17153 6837 17156
rect 6871 17153 6883 17187
rect 8036 17184 8064 17280
rect 10134 17212 10140 17264
rect 10192 17252 10198 17264
rect 10965 17255 11023 17261
rect 10965 17252 10977 17255
rect 10192 17224 10977 17252
rect 10192 17212 10198 17224
rect 10965 17221 10977 17224
rect 11011 17221 11023 17255
rect 10965 17215 11023 17221
rect 11701 17255 11759 17261
rect 11701 17221 11713 17255
rect 11747 17252 11759 17255
rect 12618 17252 12624 17264
rect 11747 17224 12624 17252
rect 11747 17221 11759 17224
rect 11701 17215 11759 17221
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 13814 17252 13820 17264
rect 12820 17224 13820 17252
rect 8573 17187 8631 17193
rect 8573 17184 8585 17187
rect 8036 17156 8585 17184
rect 6825 17147 6883 17153
rect 8573 17153 8585 17156
rect 8619 17153 8631 17187
rect 8573 17147 8631 17153
rect 10413 17187 10471 17193
rect 10413 17153 10425 17187
rect 10459 17184 10471 17187
rect 11054 17184 11060 17196
rect 10459 17156 11060 17184
rect 10459 17153 10471 17156
rect 10413 17147 10471 17153
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 2593 17119 2651 17125
rect 1443 17088 2084 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 2056 16992 2084 17088
rect 2593 17085 2605 17119
rect 2639 17085 2651 17119
rect 2593 17079 2651 17085
rect 3672 17119 3730 17125
rect 3672 17085 3684 17119
rect 3718 17116 3730 17119
rect 4065 17119 4123 17125
rect 4065 17116 4077 17119
rect 3718 17088 4077 17116
rect 3718 17085 3730 17088
rect 3672 17079 3730 17085
rect 4065 17085 4077 17088
rect 4111 17085 4123 17119
rect 4065 17079 4123 17085
rect 2038 16980 2044 16992
rect 1999 16952 2044 16980
rect 2038 16940 2044 16952
rect 2096 16940 2102 16992
rect 2130 16940 2136 16992
rect 2188 16980 2194 16992
rect 2409 16983 2467 16989
rect 2409 16980 2421 16983
rect 2188 16952 2421 16980
rect 2188 16940 2194 16952
rect 2409 16949 2421 16952
rect 2455 16980 2467 16983
rect 2590 16980 2596 16992
rect 2455 16952 2596 16980
rect 2455 16949 2467 16952
rect 2409 16943 2467 16949
rect 2590 16940 2596 16952
rect 2648 16940 2654 16992
rect 2774 16940 2780 16992
rect 2832 16980 2838 16992
rect 3743 16983 3801 16989
rect 2832 16952 2877 16980
rect 2832 16940 2838 16952
rect 3743 16949 3755 16983
rect 3789 16980 3801 16983
rect 3970 16980 3976 16992
rect 3789 16952 3976 16980
rect 3789 16949 3801 16952
rect 3743 16943 3801 16949
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 4080 16980 4108 17079
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 12820 17125 12848 17224
rect 13814 17212 13820 17224
rect 13872 17212 13878 17264
rect 17037 17255 17095 17261
rect 17037 17221 17049 17255
rect 17083 17252 17095 17255
rect 18230 17252 18236 17264
rect 17083 17224 18236 17252
rect 17083 17221 17095 17224
rect 17037 17215 17095 17221
rect 18230 17212 18236 17224
rect 18288 17212 18294 17264
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17184 13599 17187
rect 14369 17187 14427 17193
rect 14369 17184 14381 17187
rect 13587 17156 14381 17184
rect 13587 17153 13599 17156
rect 13541 17147 13599 17153
rect 14369 17153 14381 17156
rect 14415 17184 14427 17187
rect 14550 17184 14556 17196
rect 14415 17156 14556 17184
rect 14415 17153 14427 17156
rect 14369 17147 14427 17153
rect 14550 17144 14556 17156
rect 14608 17144 14614 17196
rect 16114 17184 16120 17196
rect 16075 17156 16120 17184
rect 16114 17144 16120 17156
rect 16172 17144 16178 17196
rect 18414 17184 18420 17196
rect 18375 17156 18420 17184
rect 18414 17144 18420 17156
rect 18472 17144 18478 17196
rect 9953 17119 10011 17125
rect 9953 17116 9965 17119
rect 9824 17088 9965 17116
rect 9824 17076 9830 17088
rect 9953 17085 9965 17088
rect 9999 17085 10011 17119
rect 12805 17119 12863 17125
rect 12805 17116 12817 17119
rect 9953 17079 10011 17085
rect 12636 17088 12817 17116
rect 4798 17008 4804 17060
rect 4856 17048 4862 17060
rect 5350 17048 5356 17060
rect 4856 17020 4901 17048
rect 5311 17020 5356 17048
rect 4856 17008 4862 17020
rect 5350 17008 5356 17020
rect 5408 17008 5414 17060
rect 8938 17057 8944 17060
rect 7146 17051 7204 17057
rect 7146 17017 7158 17051
rect 7192 17048 7204 17051
rect 8894 17051 8944 17057
rect 8894 17048 8906 17051
rect 7192 17020 7226 17048
rect 8404 17020 8906 17048
rect 7192 17017 7204 17020
rect 7146 17011 7204 17017
rect 4982 16980 4988 16992
rect 4080 16952 4988 16980
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 6089 16983 6147 16989
rect 6089 16949 6101 16983
rect 6135 16980 6147 16983
rect 6178 16980 6184 16992
rect 6135 16952 6184 16980
rect 6135 16949 6147 16952
rect 6089 16943 6147 16949
rect 6178 16940 6184 16952
rect 6236 16980 6242 16992
rect 6362 16980 6368 16992
rect 6236 16952 6368 16980
rect 6236 16940 6242 16952
rect 6362 16940 6368 16952
rect 6420 16980 6426 16992
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6420 16952 6561 16980
rect 6420 16940 6426 16952
rect 6549 16949 6561 16952
rect 6595 16980 6607 16983
rect 7161 16980 7189 17011
rect 8404 16989 8432 17020
rect 8894 17017 8906 17020
rect 8940 17017 8944 17051
rect 8894 17011 8944 17017
rect 8938 17008 8944 17011
rect 8996 17048 9002 17060
rect 9861 17051 9919 17057
rect 8996 17020 9042 17048
rect 8996 17008 9002 17020
rect 9861 17017 9873 17051
rect 9907 17048 9919 17051
rect 10229 17051 10287 17057
rect 10229 17048 10241 17051
rect 9907 17020 10241 17048
rect 9907 17017 9919 17020
rect 9861 17011 9919 17017
rect 10229 17017 10241 17020
rect 10275 17048 10287 17051
rect 10505 17051 10563 17057
rect 10505 17048 10517 17051
rect 10275 17020 10517 17048
rect 10275 17017 10287 17020
rect 10229 17011 10287 17017
rect 10505 17017 10517 17020
rect 10551 17048 10563 17051
rect 10778 17048 10784 17060
rect 10551 17020 10784 17048
rect 10551 17017 10563 17020
rect 10505 17011 10563 17017
rect 10778 17008 10784 17020
rect 10836 17008 10842 17060
rect 8389 16983 8447 16989
rect 8389 16980 8401 16983
rect 6595 16952 8401 16980
rect 6595 16949 6607 16952
rect 6549 16943 6607 16949
rect 8389 16949 8401 16952
rect 8435 16949 8447 16983
rect 9490 16980 9496 16992
rect 9451 16952 9496 16980
rect 8389 16943 8447 16949
rect 9490 16940 9496 16952
rect 9548 16980 9554 16992
rect 9766 16980 9772 16992
rect 9548 16952 9772 16980
rect 9548 16940 9554 16952
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 9950 16980 9956 16992
rect 9911 16952 9956 16980
rect 9950 16940 9956 16952
rect 10008 16940 10014 16992
rect 11422 16940 11428 16992
rect 11480 16980 11486 16992
rect 11977 16983 12035 16989
rect 11977 16980 11989 16983
rect 11480 16952 11989 16980
rect 11480 16940 11486 16952
rect 11977 16949 11989 16952
rect 12023 16949 12035 16983
rect 11977 16943 12035 16949
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 12636 16989 12664 17088
rect 12805 17085 12817 17088
rect 12851 17085 12863 17119
rect 13262 17116 13268 17128
rect 13223 17088 13268 17116
rect 12805 17079 12863 17085
rect 13262 17076 13268 17088
rect 13320 17076 13326 17128
rect 17770 17116 17776 17128
rect 17731 17088 17776 17116
rect 17770 17076 17776 17088
rect 17828 17076 17834 17128
rect 18874 17076 18880 17128
rect 18932 17116 18938 17128
rect 20714 17125 20720 17128
rect 19680 17119 19738 17125
rect 19680 17116 19692 17119
rect 18932 17088 19692 17116
rect 18932 17076 18938 17088
rect 19680 17085 19692 17088
rect 19726 17116 19738 17119
rect 20692 17119 20720 17125
rect 19726 17088 20208 17116
rect 19726 17085 19738 17088
rect 19680 17079 19738 17085
rect 13446 17008 13452 17060
rect 13504 17048 13510 17060
rect 14734 17057 14740 17060
rect 14185 17051 14243 17057
rect 14185 17048 14197 17051
rect 13504 17020 14197 17048
rect 13504 17008 13510 17020
rect 14185 17017 14197 17020
rect 14231 17048 14243 17051
rect 14690 17051 14740 17057
rect 14690 17048 14702 17051
rect 14231 17020 14702 17048
rect 14231 17017 14243 17020
rect 14185 17011 14243 17017
rect 14690 17017 14702 17020
rect 14736 17017 14740 17051
rect 14690 17011 14740 17017
rect 14734 17008 14740 17011
rect 14792 17048 14798 17060
rect 15933 17051 15991 17057
rect 15933 17048 15945 17051
rect 14792 17020 15945 17048
rect 14792 17008 14798 17020
rect 15933 17017 15945 17020
rect 15979 17048 15991 17051
rect 16438 17051 16496 17057
rect 16438 17048 16450 17051
rect 15979 17020 16450 17048
rect 15979 17017 15991 17020
rect 15933 17011 15991 17017
rect 16438 17017 16450 17020
rect 16484 17048 16496 17051
rect 16942 17048 16948 17060
rect 16484 17020 16948 17048
rect 16484 17017 16496 17020
rect 16438 17011 16496 17017
rect 16942 17008 16948 17020
rect 17000 17048 17006 17060
rect 17313 17051 17371 17057
rect 17313 17048 17325 17051
rect 17000 17020 17325 17048
rect 17000 17008 17006 17020
rect 17313 17017 17325 17020
rect 17359 17017 17371 17051
rect 18138 17048 18144 17060
rect 18099 17020 18144 17048
rect 17313 17011 17371 17017
rect 18138 17008 18144 17020
rect 18196 17008 18202 17060
rect 18230 17008 18236 17060
rect 18288 17048 18294 17060
rect 20180 17057 20208 17088
rect 20692 17085 20704 17119
rect 20772 17116 20778 17128
rect 21453 17119 21511 17125
rect 21453 17116 21465 17119
rect 20772 17088 21465 17116
rect 20692 17079 20720 17085
rect 20714 17076 20720 17079
rect 20772 17076 20778 17088
rect 21453 17085 21465 17088
rect 21499 17085 21511 17119
rect 21453 17079 21511 17085
rect 21704 17119 21762 17125
rect 21704 17085 21716 17119
rect 21750 17116 21762 17119
rect 22097 17119 22155 17125
rect 22097 17116 22109 17119
rect 21750 17088 22109 17116
rect 21750 17085 21762 17088
rect 21704 17079 21762 17085
rect 22097 17085 22109 17088
rect 22143 17116 22155 17119
rect 22186 17116 22192 17128
rect 22143 17088 22192 17116
rect 22143 17085 22155 17088
rect 22097 17079 22155 17085
rect 22186 17076 22192 17088
rect 22244 17076 22250 17128
rect 24118 17076 24124 17128
rect 24176 17116 24182 17128
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 24176 17088 24593 17116
rect 24176 17076 24182 17088
rect 24581 17085 24593 17088
rect 24627 17116 24639 17119
rect 25133 17119 25191 17125
rect 25133 17116 25145 17119
rect 24627 17088 25145 17116
rect 24627 17085 24639 17088
rect 24581 17079 24639 17085
rect 25133 17085 25145 17088
rect 25179 17085 25191 17119
rect 25133 17079 25191 17085
rect 20165 17051 20223 17057
rect 18288 17020 18333 17048
rect 18288 17008 18294 17020
rect 20165 17017 20177 17051
rect 20211 17048 20223 17051
rect 25038 17048 25044 17060
rect 20211 17020 25044 17048
rect 20211 17017 20223 17020
rect 20165 17011 20223 17017
rect 25038 17008 25044 17020
rect 25096 17008 25102 17060
rect 12621 16983 12679 16989
rect 12621 16980 12633 16983
rect 12584 16952 12633 16980
rect 12584 16940 12590 16952
rect 12621 16949 12633 16952
rect 12667 16949 12679 16983
rect 12621 16943 12679 16949
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 13817 16983 13875 16989
rect 13817 16980 13829 16983
rect 12952 16952 13829 16980
rect 12952 16940 12958 16952
rect 13817 16949 13829 16952
rect 13863 16949 13875 16983
rect 15286 16980 15292 16992
rect 15247 16952 15292 16980
rect 13817 16943 13875 16949
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 15657 16983 15715 16989
rect 15657 16949 15669 16983
rect 15703 16980 15715 16983
rect 15746 16980 15752 16992
rect 15703 16952 15752 16980
rect 15703 16949 15715 16952
rect 15657 16943 15715 16949
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 18690 16940 18696 16992
rect 18748 16980 18754 16992
rect 19061 16983 19119 16989
rect 19061 16980 19073 16983
rect 18748 16952 19073 16980
rect 18748 16940 18754 16952
rect 19061 16949 19073 16952
rect 19107 16949 19119 16983
rect 19061 16943 19119 16949
rect 19518 16940 19524 16992
rect 19576 16980 19582 16992
rect 19751 16983 19809 16989
rect 19751 16980 19763 16983
rect 19576 16952 19763 16980
rect 19576 16940 19582 16952
rect 19751 16949 19763 16952
rect 19797 16949 19809 16983
rect 19751 16943 19809 16949
rect 20714 16940 20720 16992
rect 20772 16989 20778 16992
rect 20772 16983 20821 16989
rect 20772 16949 20775 16983
rect 20809 16949 20821 16983
rect 20772 16943 20821 16949
rect 20772 16940 20778 16943
rect 21542 16940 21548 16992
rect 21600 16980 21606 16992
rect 21775 16983 21833 16989
rect 21775 16980 21787 16983
rect 21600 16952 21787 16980
rect 21600 16940 21606 16952
rect 21775 16949 21787 16952
rect 21821 16949 21833 16983
rect 21775 16943 21833 16949
rect 22557 16983 22615 16989
rect 22557 16949 22569 16983
rect 22603 16980 22615 16983
rect 22830 16980 22836 16992
rect 22603 16952 22836 16980
rect 22603 16949 22615 16952
rect 22557 16943 22615 16949
rect 22830 16940 22836 16952
rect 22888 16940 22894 16992
rect 23293 16983 23351 16989
rect 23293 16949 23305 16983
rect 23339 16980 23351 16983
rect 23382 16980 23388 16992
rect 23339 16952 23388 16980
rect 23339 16949 23351 16952
rect 23293 16943 23351 16949
rect 23382 16940 23388 16952
rect 23440 16940 23446 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 3099 16779 3157 16785
rect 3099 16745 3111 16779
rect 3145 16776 3157 16779
rect 4062 16776 4068 16788
rect 3145 16748 4068 16776
rect 3145 16745 3157 16748
rect 3099 16739 3157 16745
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 4985 16779 5043 16785
rect 4985 16745 4997 16779
rect 5031 16776 5043 16779
rect 6822 16776 6828 16788
rect 5031 16748 6040 16776
rect 6783 16748 6828 16776
rect 5031 16745 5043 16748
rect 4985 16739 5043 16745
rect 6012 16720 6040 16748
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 7561 16779 7619 16785
rect 7561 16745 7573 16779
rect 7607 16776 7619 16779
rect 7926 16776 7932 16788
rect 7607 16748 7932 16776
rect 7607 16745 7619 16748
rect 7561 16739 7619 16745
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 8662 16776 8668 16788
rect 8623 16748 8668 16776
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 11054 16776 11060 16788
rect 11015 16748 11060 16776
rect 11054 16736 11060 16748
rect 11112 16776 11118 16788
rect 12434 16776 12440 16788
rect 11112 16748 12440 16776
rect 11112 16736 11118 16748
rect 12434 16736 12440 16748
rect 12492 16736 12498 16788
rect 14182 16736 14188 16788
rect 14240 16776 14246 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 14240 16748 14381 16776
rect 14240 16736 14246 16748
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 16666 16776 16672 16788
rect 16627 16748 16672 16776
rect 14369 16739 14427 16745
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 18138 16736 18144 16788
rect 18196 16776 18202 16788
rect 18601 16779 18659 16785
rect 18601 16776 18613 16779
rect 18196 16748 18613 16776
rect 18196 16736 18202 16748
rect 18601 16745 18613 16748
rect 18647 16776 18659 16779
rect 21039 16779 21097 16785
rect 18647 16748 19932 16776
rect 18647 16745 18659 16748
rect 18601 16739 18659 16745
rect 19904 16720 19932 16748
rect 21039 16745 21051 16779
rect 21085 16776 21097 16779
rect 21266 16776 21272 16788
rect 21085 16748 21272 16776
rect 21085 16745 21097 16748
rect 21039 16739 21097 16745
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 4246 16668 4252 16720
rect 4304 16708 4310 16720
rect 4386 16711 4444 16717
rect 4386 16708 4398 16711
rect 4304 16680 4398 16708
rect 4304 16668 4310 16680
rect 4386 16677 4398 16680
rect 4432 16677 4444 16711
rect 4386 16671 4444 16677
rect 4706 16668 4712 16720
rect 4764 16708 4770 16720
rect 5261 16711 5319 16717
rect 5261 16708 5273 16711
rect 4764 16680 5273 16708
rect 4764 16668 4770 16680
rect 5261 16677 5273 16680
rect 5307 16677 5319 16711
rect 5994 16708 6000 16720
rect 5907 16680 6000 16708
rect 5261 16671 5319 16677
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 7834 16708 7840 16720
rect 7795 16680 7840 16708
rect 7834 16668 7840 16680
rect 7892 16668 7898 16720
rect 9582 16668 9588 16720
rect 9640 16708 9646 16720
rect 9769 16711 9827 16717
rect 9769 16708 9781 16711
rect 9640 16680 9781 16708
rect 9640 16668 9646 16680
rect 9769 16677 9781 16680
rect 9815 16677 9827 16711
rect 9769 16671 9827 16677
rect 9858 16668 9864 16720
rect 9916 16708 9922 16720
rect 10781 16711 10839 16717
rect 9916 16680 10732 16708
rect 9916 16668 9922 16680
rect 1949 16643 2007 16649
rect 1949 16609 1961 16643
rect 1995 16640 2007 16643
rect 2130 16640 2136 16652
rect 1995 16612 2136 16640
rect 1995 16609 2007 16612
rect 1949 16603 2007 16609
rect 2130 16600 2136 16612
rect 2188 16600 2194 16652
rect 2774 16600 2780 16652
rect 2832 16640 2838 16652
rect 3028 16643 3086 16649
rect 3028 16640 3040 16643
rect 2832 16612 3040 16640
rect 2832 16600 2838 16612
rect 3028 16609 3040 16612
rect 3074 16640 3086 16643
rect 3694 16640 3700 16652
rect 3074 16612 3700 16640
rect 3074 16609 3086 16612
rect 3028 16603 3086 16609
rect 3694 16600 3700 16612
rect 3752 16600 3758 16652
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 4080 16572 4108 16603
rect 5350 16600 5356 16652
rect 5408 16640 5414 16652
rect 10704 16640 10732 16680
rect 10781 16677 10793 16711
rect 10827 16708 10839 16711
rect 10962 16708 10968 16720
rect 10827 16680 10968 16708
rect 10827 16677 10839 16680
rect 10781 16671 10839 16677
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 11330 16708 11336 16720
rect 11164 16680 11336 16708
rect 11164 16640 11192 16680
rect 11330 16668 11336 16680
rect 11388 16708 11394 16720
rect 11425 16711 11483 16717
rect 11425 16708 11437 16711
rect 11388 16680 11437 16708
rect 11388 16668 11394 16680
rect 11425 16677 11437 16680
rect 11471 16677 11483 16711
rect 11425 16671 11483 16677
rect 12342 16668 12348 16720
rect 12400 16708 12406 16720
rect 12805 16711 12863 16717
rect 12805 16708 12817 16711
rect 12400 16680 12817 16708
rect 12400 16668 12406 16680
rect 12805 16677 12817 16680
rect 12851 16708 12863 16711
rect 13262 16708 13268 16720
rect 12851 16680 13268 16708
rect 12851 16677 12863 16680
rect 12805 16671 12863 16677
rect 13262 16668 13268 16680
rect 13320 16668 13326 16720
rect 13446 16668 13452 16720
rect 13504 16717 13510 16720
rect 13504 16711 13552 16717
rect 13504 16677 13506 16711
rect 13540 16677 13552 16711
rect 13504 16671 13552 16677
rect 13504 16668 13510 16671
rect 15286 16668 15292 16720
rect 15344 16708 15350 16720
rect 15749 16711 15807 16717
rect 15749 16708 15761 16711
rect 15344 16680 15761 16708
rect 15344 16668 15350 16680
rect 15749 16677 15761 16680
rect 15795 16708 15807 16711
rect 15838 16708 15844 16720
rect 15795 16680 15844 16708
rect 15795 16677 15807 16680
rect 15749 16671 15807 16677
rect 15838 16668 15844 16680
rect 15896 16668 15902 16720
rect 17494 16668 17500 16720
rect 17552 16708 17558 16720
rect 17773 16711 17831 16717
rect 17773 16708 17785 16711
rect 17552 16680 17785 16708
rect 17552 16668 17558 16680
rect 17773 16677 17785 16680
rect 17819 16677 17831 16711
rect 19337 16711 19395 16717
rect 19337 16708 19349 16711
rect 17773 16671 17831 16677
rect 19076 16680 19349 16708
rect 5408 16612 5488 16640
rect 10704 16612 11192 16640
rect 15105 16643 15163 16649
rect 5408 16600 5414 16612
rect 4338 16572 4344 16584
rect 4080 16544 4344 16572
rect 4338 16532 4344 16544
rect 4396 16532 4402 16584
rect 5460 16572 5488 16612
rect 15105 16609 15117 16643
rect 15151 16640 15163 16643
rect 15151 16612 15424 16640
rect 15151 16609 15163 16612
rect 15105 16603 15163 16609
rect 5902 16572 5908 16584
rect 5460 16544 5580 16572
rect 5863 16544 5908 16572
rect 3326 16464 3332 16516
rect 3384 16504 3390 16516
rect 4062 16504 4068 16516
rect 3384 16476 4068 16504
rect 3384 16464 3390 16476
rect 4062 16464 4068 16476
rect 4120 16464 4126 16516
rect 5552 16504 5580 16544
rect 5902 16532 5908 16544
rect 5960 16572 5966 16584
rect 6178 16572 6184 16584
rect 5960 16544 6184 16572
rect 5960 16532 5966 16544
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 6549 16575 6607 16581
rect 6549 16541 6561 16575
rect 6595 16572 6607 16575
rect 6822 16572 6828 16584
rect 6595 16544 6828 16572
rect 6595 16541 6607 16544
rect 6549 16535 6607 16541
rect 6564 16504 6592 16535
rect 6822 16532 6828 16544
rect 6880 16532 6886 16584
rect 7742 16572 7748 16584
rect 7703 16544 7748 16572
rect 7742 16532 7748 16544
rect 7800 16532 7806 16584
rect 8018 16572 8024 16584
rect 7979 16544 8024 16572
rect 8018 16532 8024 16544
rect 8076 16532 8082 16584
rect 8662 16532 8668 16584
rect 8720 16572 8726 16584
rect 10045 16575 10103 16581
rect 10045 16572 10057 16575
rect 8720 16544 10057 16572
rect 8720 16532 8726 16544
rect 10045 16541 10057 16544
rect 10091 16572 10103 16575
rect 10134 16572 10140 16584
rect 10091 16544 10140 16572
rect 10091 16541 10103 16544
rect 10045 16535 10103 16541
rect 10134 16532 10140 16544
rect 10192 16532 10198 16584
rect 11333 16575 11391 16581
rect 11333 16541 11345 16575
rect 11379 16572 11391 16575
rect 11514 16572 11520 16584
rect 11379 16544 11520 16572
rect 11379 16541 11391 16544
rect 11333 16535 11391 16541
rect 11514 16532 11520 16544
rect 11572 16532 11578 16584
rect 11698 16572 11704 16584
rect 11659 16544 11704 16572
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 13170 16572 13176 16584
rect 13131 16544 13176 16572
rect 13170 16532 13176 16544
rect 13228 16532 13234 16584
rect 15396 16572 15424 16612
rect 18966 16600 18972 16652
rect 19024 16600 19030 16652
rect 15470 16572 15476 16584
rect 15383 16544 15476 16572
rect 15470 16532 15476 16544
rect 15528 16572 15534 16584
rect 15657 16575 15715 16581
rect 15657 16572 15669 16575
rect 15528 16544 15669 16572
rect 15528 16532 15534 16544
rect 15657 16541 15669 16544
rect 15703 16541 15715 16575
rect 15657 16535 15715 16541
rect 17497 16575 17555 16581
rect 17497 16541 17509 16575
rect 17543 16572 17555 16575
rect 17678 16572 17684 16584
rect 17543 16544 17684 16572
rect 17543 16541 17555 16544
rect 17497 16535 17555 16541
rect 17678 16532 17684 16544
rect 17736 16532 17742 16584
rect 17957 16575 18015 16581
rect 17957 16541 17969 16575
rect 18003 16572 18015 16575
rect 18414 16572 18420 16584
rect 18003 16544 18420 16572
rect 18003 16541 18015 16544
rect 17957 16535 18015 16541
rect 5552 16476 6592 16504
rect 14093 16507 14151 16513
rect 14093 16473 14105 16507
rect 14139 16504 14151 16507
rect 14734 16504 14740 16516
rect 14139 16476 14740 16504
rect 14139 16473 14151 16476
rect 14093 16467 14151 16473
rect 14734 16464 14740 16476
rect 14792 16464 14798 16516
rect 16209 16507 16267 16513
rect 16209 16473 16221 16507
rect 16255 16504 16267 16507
rect 17972 16504 18000 16535
rect 18414 16532 18420 16544
rect 18472 16532 18478 16584
rect 16255 16476 18000 16504
rect 18984 16504 19012 16600
rect 19076 16584 19104 16680
rect 19337 16677 19349 16680
rect 19383 16677 19395 16711
rect 19886 16708 19892 16720
rect 19799 16680 19892 16708
rect 19337 16671 19395 16677
rect 19886 16668 19892 16680
rect 19944 16668 19950 16720
rect 24670 16668 24676 16720
rect 24728 16708 24734 16720
rect 25087 16711 25145 16717
rect 25087 16708 25099 16711
rect 24728 16680 25099 16708
rect 24728 16668 24734 16680
rect 25087 16677 25099 16680
rect 25133 16677 25145 16711
rect 25087 16671 25145 16677
rect 20968 16643 21026 16649
rect 20968 16609 20980 16643
rect 21014 16640 21026 16643
rect 21082 16640 21088 16652
rect 21014 16612 21088 16640
rect 21014 16609 21026 16612
rect 20968 16603 21026 16609
rect 21082 16600 21088 16612
rect 21140 16600 21146 16652
rect 21980 16643 22038 16649
rect 21980 16609 21992 16643
rect 22026 16640 22038 16643
rect 22026 16609 22048 16640
rect 21980 16603 22048 16609
rect 19058 16532 19064 16584
rect 19116 16532 19122 16584
rect 19245 16575 19303 16581
rect 19245 16541 19257 16575
rect 19291 16541 19303 16575
rect 22020 16572 22048 16603
rect 22922 16600 22928 16652
rect 22980 16649 22986 16652
rect 23106 16649 23112 16652
rect 22980 16643 23018 16649
rect 23006 16609 23018 16643
rect 22980 16603 23018 16609
rect 23063 16643 23112 16649
rect 23063 16609 23075 16643
rect 23109 16609 23112 16643
rect 23063 16603 23112 16609
rect 22980 16600 22986 16603
rect 23106 16600 23112 16603
rect 23164 16600 23170 16652
rect 23937 16643 23995 16649
rect 23937 16640 23949 16643
rect 23216 16612 23949 16640
rect 22278 16572 22284 16584
rect 22020 16544 22284 16572
rect 19245 16535 19303 16541
rect 19260 16504 19288 16535
rect 22278 16532 22284 16544
rect 22336 16532 22342 16584
rect 22646 16532 22652 16584
rect 22704 16572 22710 16584
rect 23216 16572 23244 16612
rect 23937 16609 23949 16612
rect 23983 16609 23995 16643
rect 23937 16603 23995 16609
rect 25000 16643 25058 16649
rect 25000 16609 25012 16643
rect 25046 16640 25058 16643
rect 25498 16640 25504 16652
rect 25046 16612 25504 16640
rect 25046 16609 25058 16612
rect 25000 16603 25058 16609
rect 25498 16600 25504 16612
rect 25556 16600 25562 16652
rect 22704 16544 23244 16572
rect 22704 16532 22710 16544
rect 20714 16504 20720 16516
rect 18984 16476 20720 16504
rect 16255 16473 16267 16476
rect 16209 16467 16267 16473
rect 20714 16464 20720 16476
rect 20772 16464 20778 16516
rect 1762 16396 1768 16448
rect 1820 16436 1826 16448
rect 1946 16436 1952 16448
rect 1820 16408 1952 16436
rect 1820 16396 1826 16408
rect 1946 16396 1952 16408
rect 2004 16396 2010 16448
rect 2038 16396 2044 16448
rect 2096 16436 2102 16448
rect 2133 16439 2191 16445
rect 2133 16436 2145 16439
rect 2096 16408 2145 16436
rect 2096 16396 2102 16408
rect 2133 16405 2145 16408
rect 2179 16405 2191 16439
rect 2133 16399 2191 16405
rect 3142 16396 3148 16448
rect 3200 16436 3206 16448
rect 8386 16436 8392 16448
rect 3200 16408 8392 16436
rect 3200 16396 3206 16408
rect 8386 16396 8392 16408
rect 8444 16396 8450 16448
rect 22051 16439 22109 16445
rect 22051 16405 22063 16439
rect 22097 16436 22109 16439
rect 25406 16436 25412 16448
rect 22097 16408 25412 16436
rect 22097 16405 22109 16408
rect 22051 16399 22109 16405
rect 25406 16396 25412 16408
rect 25464 16396 25470 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1394 16192 1400 16244
rect 1452 16232 1458 16244
rect 1581 16235 1639 16241
rect 1581 16232 1593 16235
rect 1452 16204 1593 16232
rect 1452 16192 1458 16204
rect 1581 16201 1593 16204
rect 1627 16201 1639 16235
rect 1581 16195 1639 16201
rect 4798 16192 4804 16244
rect 4856 16232 4862 16244
rect 5077 16235 5135 16241
rect 5077 16232 5089 16235
rect 4856 16204 5089 16232
rect 4856 16192 4862 16204
rect 5077 16201 5089 16204
rect 5123 16201 5135 16235
rect 5077 16195 5135 16201
rect 5905 16235 5963 16241
rect 5905 16201 5917 16235
rect 5951 16232 5963 16235
rect 5994 16232 6000 16244
rect 5951 16204 6000 16232
rect 5951 16201 5963 16204
rect 5905 16195 5963 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 6178 16232 6184 16244
rect 6139 16204 6184 16232
rect 6178 16192 6184 16204
rect 6236 16192 6242 16244
rect 6638 16232 6644 16244
rect 6599 16204 6644 16232
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 7193 16235 7251 16241
rect 7193 16201 7205 16235
rect 7239 16232 7251 16235
rect 7561 16235 7619 16241
rect 7561 16232 7573 16235
rect 7239 16204 7573 16232
rect 7239 16201 7251 16204
rect 7193 16195 7251 16201
rect 7561 16201 7573 16204
rect 7607 16232 7619 16235
rect 7834 16232 7840 16244
rect 7607 16204 7840 16232
rect 7607 16201 7619 16204
rect 7561 16195 7619 16201
rect 7834 16192 7840 16204
rect 7892 16192 7898 16244
rect 9033 16235 9091 16241
rect 9033 16201 9045 16235
rect 9079 16232 9091 16235
rect 9490 16232 9496 16244
rect 9079 16204 9496 16232
rect 9079 16201 9091 16204
rect 9033 16195 9091 16201
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 10778 16232 10784 16244
rect 10739 16204 10784 16232
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 11330 16232 11336 16244
rect 11291 16204 11336 16232
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 14001 16235 14059 16241
rect 14001 16201 14013 16235
rect 14047 16232 14059 16235
rect 15657 16235 15715 16241
rect 15657 16232 15669 16235
rect 14047 16204 15669 16232
rect 14047 16201 14059 16204
rect 14001 16195 14059 16201
rect 15657 16201 15669 16204
rect 15703 16201 15715 16235
rect 15838 16232 15844 16244
rect 15799 16204 15844 16232
rect 15657 16195 15715 16201
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 17494 16232 17500 16244
rect 17455 16204 17500 16232
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 24762 16232 24768 16244
rect 24723 16204 24768 16232
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 2314 16124 2320 16176
rect 2372 16164 2378 16176
rect 9122 16164 9128 16176
rect 2372 16136 9128 16164
rect 2372 16124 2378 16136
rect 9122 16124 9128 16136
rect 9180 16124 9186 16176
rect 15470 16164 15476 16176
rect 15431 16136 15476 16164
rect 15470 16124 15476 16136
rect 15528 16164 15534 16176
rect 15528 16136 16804 16164
rect 15528 16124 15534 16136
rect 2038 16096 2044 16108
rect 1412 16068 2044 16096
rect 1412 16037 1440 16068
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16096 4123 16099
rect 4111 16068 4292 16096
rect 4111 16065 4123 16068
rect 4065 16059 4123 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 1397 15991 1455 15997
rect 2501 16031 2559 16037
rect 2501 15997 2513 16031
rect 2547 16028 2559 16031
rect 2866 16028 2872 16040
rect 2547 16000 2872 16028
rect 2547 15997 2559 16000
rect 2501 15991 2559 15997
rect 2866 15988 2872 16000
rect 2924 15988 2930 16040
rect 3145 16031 3203 16037
rect 3145 15997 3157 16031
rect 3191 16028 3203 16031
rect 3602 16028 3608 16040
rect 3191 16000 3608 16028
rect 3191 15997 3203 16000
rect 3145 15991 3203 15997
rect 3602 15988 3608 16000
rect 3660 15988 3666 16040
rect 4157 16031 4215 16037
rect 4157 15997 4169 16031
rect 4203 15997 4215 16031
rect 4157 15991 4215 15997
rect 3326 15960 3332 15972
rect 3287 15932 3332 15960
rect 3326 15920 3332 15932
rect 3384 15920 3390 15972
rect 3694 15960 3700 15972
rect 3655 15932 3700 15960
rect 3694 15920 3700 15932
rect 3752 15920 3758 15972
rect 4172 15892 4200 15991
rect 4264 15972 4292 16068
rect 7466 16056 7472 16108
rect 7524 16096 7530 16108
rect 7745 16099 7803 16105
rect 7745 16096 7757 16099
rect 7524 16068 7757 16096
rect 7524 16056 7530 16068
rect 7745 16065 7757 16068
rect 7791 16096 7803 16099
rect 8110 16096 8116 16108
rect 7791 16068 8116 16096
rect 7791 16065 7803 16068
rect 7745 16059 7803 16065
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 8389 16099 8447 16105
rect 8389 16065 8401 16099
rect 8435 16096 8447 16099
rect 8662 16096 8668 16108
rect 8435 16068 8668 16096
rect 8435 16065 8447 16068
rect 8389 16059 8447 16065
rect 8662 16056 8668 16068
rect 8720 16056 8726 16108
rect 14642 16096 14648 16108
rect 14603 16068 14648 16096
rect 14642 16056 14648 16068
rect 14700 16096 14706 16108
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14700 16068 14933 16096
rect 14700 16056 14706 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15194 16056 15200 16108
rect 15252 16096 15258 16108
rect 16482 16096 16488 16108
rect 15252 16068 16488 16096
rect 15252 16056 15258 16068
rect 16482 16056 16488 16068
rect 16540 16056 16546 16108
rect 16776 16105 16804 16136
rect 19426 16124 19432 16176
rect 19484 16164 19490 16176
rect 19484 16136 19932 16164
rect 19484 16124 19490 16136
rect 19904 16108 19932 16136
rect 16761 16099 16819 16105
rect 16761 16065 16773 16099
rect 16807 16065 16819 16099
rect 16761 16059 16819 16065
rect 18141 16099 18199 16105
rect 18141 16065 18153 16099
rect 18187 16096 18199 16099
rect 18598 16096 18604 16108
rect 18187 16068 18604 16096
rect 18187 16065 18199 16068
rect 18141 16059 18199 16065
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 19518 16056 19524 16108
rect 19576 16096 19582 16108
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 19576 16068 19717 16096
rect 19576 16056 19582 16068
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 19705 16059 19763 16065
rect 19886 16056 19892 16108
rect 19944 16096 19950 16108
rect 19981 16099 20039 16105
rect 19981 16096 19993 16099
rect 19944 16068 19993 16096
rect 19944 16056 19950 16068
rect 19981 16065 19993 16068
rect 20027 16065 20039 16099
rect 21082 16096 21088 16108
rect 20995 16068 21088 16096
rect 19981 16059 20039 16065
rect 21082 16056 21088 16068
rect 21140 16096 21146 16108
rect 21726 16096 21732 16108
rect 21140 16068 21732 16096
rect 21140 16056 21146 16068
rect 21726 16056 21732 16068
rect 21784 16056 21790 16108
rect 9861 16031 9919 16037
rect 9861 16028 9873 16031
rect 9324 16000 9873 16028
rect 4246 15920 4252 15972
rect 4304 15960 4310 15972
rect 4519 15963 4577 15969
rect 4519 15960 4531 15963
rect 4304 15932 4531 15960
rect 4304 15920 4310 15932
rect 4519 15929 4531 15932
rect 4565 15960 4577 15963
rect 6362 15960 6368 15972
rect 4565 15932 6368 15960
rect 4565 15929 4577 15932
rect 4519 15923 4577 15929
rect 6362 15920 6368 15932
rect 6420 15920 6426 15972
rect 7834 15920 7840 15972
rect 7892 15960 7898 15972
rect 7892 15932 7937 15960
rect 7892 15920 7898 15932
rect 9324 15904 9352 16000
rect 9861 15997 9873 16000
rect 9907 15997 9919 16031
rect 13078 16028 13084 16040
rect 12991 16000 13084 16028
rect 9861 15991 9919 15997
rect 13078 15988 13084 16000
rect 13136 16028 13142 16040
rect 14277 16031 14335 16037
rect 14277 16028 14289 16031
rect 13136 16000 14289 16028
rect 13136 15988 13142 16000
rect 14277 15997 14289 16000
rect 14323 15997 14335 16031
rect 14277 15991 14335 15997
rect 15657 16031 15715 16037
rect 15657 15997 15669 16031
rect 15703 16028 15715 16031
rect 16209 16031 16267 16037
rect 16209 16028 16221 16031
rect 15703 16000 16221 16028
rect 15703 15997 15715 16000
rect 15657 15991 15715 15997
rect 16209 15997 16221 16000
rect 16255 16028 16267 16031
rect 16298 16028 16304 16040
rect 16255 16000 16304 16028
rect 16255 15997 16267 16000
rect 16209 15991 16267 15997
rect 16298 15988 16304 16000
rect 16356 15988 16362 16040
rect 21228 16031 21286 16037
rect 21228 15997 21240 16031
rect 21274 16028 21286 16031
rect 22224 16031 22282 16037
rect 21274 16000 21772 16028
rect 21274 15997 21286 16000
rect 21228 15991 21286 15997
rect 13446 15969 13452 15972
rect 10182 15963 10240 15969
rect 10182 15960 10194 15963
rect 9876 15932 10194 15960
rect 9876 15904 9904 15932
rect 10182 15929 10194 15932
rect 10228 15929 10240 15963
rect 13402 15963 13452 15969
rect 13402 15960 13414 15963
rect 10182 15923 10240 15929
rect 13280 15932 13414 15960
rect 13280 15904 13308 15932
rect 13402 15929 13414 15932
rect 13448 15929 13452 15963
rect 13402 15923 13452 15929
rect 13446 15920 13452 15923
rect 13504 15960 13510 15972
rect 15013 15963 15071 15969
rect 13504 15932 13550 15960
rect 13504 15920 13510 15932
rect 15013 15929 15025 15963
rect 15059 15960 15071 15963
rect 16574 15960 16580 15972
rect 15059 15932 16436 15960
rect 16535 15932 16580 15960
rect 15059 15929 15071 15932
rect 15013 15923 15071 15929
rect 5350 15892 5356 15904
rect 4172 15864 5356 15892
rect 5350 15852 5356 15864
rect 5408 15852 5414 15904
rect 9306 15892 9312 15904
rect 9267 15864 9312 15892
rect 9306 15852 9312 15864
rect 9364 15852 9370 15904
rect 9769 15895 9827 15901
rect 9769 15861 9781 15895
rect 9815 15892 9827 15895
rect 9858 15892 9864 15904
rect 9815 15864 9864 15892
rect 9815 15861 9827 15864
rect 9769 15855 9827 15861
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 11609 15895 11667 15901
rect 11609 15892 11621 15895
rect 11572 15864 11621 15892
rect 11572 15852 11578 15864
rect 11609 15861 11621 15864
rect 11655 15861 11667 15895
rect 11609 15855 11667 15861
rect 12253 15895 12311 15901
rect 12253 15861 12265 15895
rect 12299 15892 12311 15895
rect 12989 15895 13047 15901
rect 12989 15892 13001 15895
rect 12299 15864 13001 15892
rect 12299 15861 12311 15864
rect 12253 15855 12311 15861
rect 12989 15861 13001 15864
rect 13035 15892 13047 15895
rect 13262 15892 13268 15904
rect 13035 15864 13268 15892
rect 13035 15861 13047 15864
rect 12989 15855 13047 15861
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 14734 15852 14740 15904
rect 14792 15892 14798 15904
rect 15028 15892 15056 15923
rect 14792 15864 15056 15892
rect 16408 15892 16436 15932
rect 16574 15920 16580 15932
rect 16632 15920 16638 15972
rect 18233 15963 18291 15969
rect 18233 15929 18245 15963
rect 18279 15929 18291 15963
rect 18782 15960 18788 15972
rect 18743 15932 18788 15960
rect 18233 15923 18291 15929
rect 17773 15895 17831 15901
rect 17773 15892 17785 15895
rect 16408 15864 17785 15892
rect 14792 15852 14798 15864
rect 17773 15861 17785 15864
rect 17819 15892 17831 15895
rect 18248 15892 18276 15923
rect 18782 15920 18788 15932
rect 18840 15920 18846 15972
rect 19797 15963 19855 15969
rect 19797 15929 19809 15963
rect 19843 15929 19855 15963
rect 19797 15923 19855 15929
rect 19058 15892 19064 15904
rect 17819 15864 19064 15892
rect 17819 15861 17831 15864
rect 17773 15855 17831 15861
rect 19058 15852 19064 15864
rect 19116 15852 19122 15904
rect 19242 15852 19248 15904
rect 19300 15892 19306 15904
rect 19429 15895 19487 15901
rect 19429 15892 19441 15895
rect 19300 15864 19441 15892
rect 19300 15852 19306 15864
rect 19429 15861 19441 15864
rect 19475 15892 19487 15895
rect 19812 15892 19840 15923
rect 20714 15920 20720 15972
rect 20772 15960 20778 15972
rect 21315 15963 21373 15969
rect 21315 15960 21327 15963
rect 20772 15932 21327 15960
rect 20772 15920 20778 15932
rect 21315 15929 21327 15932
rect 21361 15929 21373 15963
rect 21315 15923 21373 15929
rect 21744 15901 21772 16000
rect 22224 15997 22236 16031
rect 22270 16028 22282 16031
rect 22270 16000 22304 16028
rect 22270 15997 22282 16000
rect 22224 15991 22282 15997
rect 22094 15960 22100 15972
rect 22007 15932 22100 15960
rect 22094 15920 22100 15932
rect 22152 15960 22158 15972
rect 22239 15960 22267 15991
rect 22922 15988 22928 16040
rect 22980 16028 22986 16040
rect 23017 16031 23075 16037
rect 23017 16028 23029 16031
rect 22980 16000 23029 16028
rect 22980 15988 22986 16000
rect 23017 15997 23029 16000
rect 23063 16028 23075 16031
rect 24581 16031 24639 16037
rect 24581 16028 24593 16031
rect 23063 16000 24593 16028
rect 23063 15997 23075 16000
rect 23017 15991 23075 15997
rect 24581 15997 24593 16000
rect 24627 16028 24639 16031
rect 25133 16031 25191 16037
rect 25133 16028 25145 16031
rect 24627 16000 25145 16028
rect 24627 15997 24639 16000
rect 24581 15991 24639 15997
rect 25133 15997 25145 16000
rect 25179 15997 25191 16031
rect 25133 15991 25191 15997
rect 22554 15960 22560 15972
rect 22152 15932 22560 15960
rect 22152 15920 22158 15932
rect 22554 15920 22560 15932
rect 22612 15920 22618 15972
rect 19475 15864 19840 15892
rect 21729 15895 21787 15901
rect 19475 15861 19487 15864
rect 19429 15855 19487 15861
rect 21729 15861 21741 15895
rect 21775 15892 21787 15895
rect 21818 15892 21824 15904
rect 21775 15864 21824 15892
rect 21775 15861 21787 15864
rect 21729 15855 21787 15861
rect 21818 15852 21824 15864
rect 21876 15852 21882 15904
rect 22186 15852 22192 15904
rect 22244 15892 22250 15904
rect 22327 15895 22385 15901
rect 22327 15892 22339 15895
rect 22244 15864 22339 15892
rect 22244 15852 22250 15864
rect 22327 15861 22339 15864
rect 22373 15861 22385 15895
rect 25498 15892 25504 15904
rect 25459 15864 25504 15892
rect 22327 15855 22385 15861
rect 25498 15852 25504 15864
rect 25556 15852 25562 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1581 15691 1639 15697
rect 1581 15657 1593 15691
rect 1627 15688 1639 15691
rect 1670 15688 1676 15700
rect 1627 15660 1676 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 4246 15688 4252 15700
rect 4207 15660 4252 15688
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 5258 15688 5264 15700
rect 5219 15660 5264 15688
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 7469 15691 7527 15697
rect 7469 15657 7481 15691
rect 7515 15688 7527 15691
rect 7834 15688 7840 15700
rect 7515 15660 7840 15688
rect 7515 15657 7527 15660
rect 7469 15651 7527 15657
rect 7834 15648 7840 15660
rect 7892 15648 7898 15700
rect 8110 15688 8116 15700
rect 8071 15660 8116 15688
rect 8110 15648 8116 15660
rect 8168 15648 8174 15700
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 9582 15688 9588 15700
rect 9539 15660 9588 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 12250 15688 12256 15700
rect 11440 15660 12256 15688
rect 4890 15580 4896 15632
rect 4948 15620 4954 15632
rect 4948 15592 5488 15620
rect 4948 15580 4954 15592
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 2406 15552 2412 15564
rect 1443 15524 2412 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 2406 15512 2412 15524
rect 2464 15512 2470 15564
rect 2958 15552 2964 15564
rect 2919 15524 2964 15552
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 5166 15552 5172 15564
rect 5127 15524 5172 15552
rect 5166 15512 5172 15524
rect 5224 15512 5230 15564
rect 5258 15512 5264 15564
rect 5316 15552 5322 15564
rect 5460 15561 5488 15592
rect 6362 15580 6368 15632
rect 6420 15620 6426 15632
rect 6822 15620 6828 15632
rect 6420 15592 6828 15620
rect 6420 15580 6426 15592
rect 6822 15580 6828 15592
rect 6880 15629 6886 15632
rect 6880 15623 6928 15629
rect 6880 15589 6882 15623
rect 6916 15589 6928 15623
rect 6880 15583 6928 15589
rect 6880 15580 6886 15583
rect 5445 15555 5503 15561
rect 5445 15552 5457 15555
rect 5316 15524 5457 15552
rect 5316 15512 5322 15524
rect 5445 15521 5457 15524
rect 5491 15521 5503 15555
rect 6546 15552 6552 15564
rect 6507 15524 6552 15552
rect 5445 15515 5503 15521
rect 6546 15512 6552 15524
rect 6604 15552 6610 15564
rect 7006 15552 7012 15564
rect 6604 15524 7012 15552
rect 6604 15512 6610 15524
rect 7006 15512 7012 15524
rect 7064 15512 7070 15564
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 8608 15555 8666 15561
rect 8608 15552 8620 15555
rect 8536 15524 8620 15552
rect 8536 15512 8542 15524
rect 8608 15521 8620 15524
rect 8654 15521 8666 15555
rect 8608 15515 8666 15521
rect 8711 15555 8769 15561
rect 8711 15521 8723 15555
rect 8757 15552 8769 15555
rect 9582 15552 9588 15564
rect 8757 15524 9588 15552
rect 8757 15521 8769 15524
rect 8711 15515 8769 15521
rect 9582 15512 9588 15524
rect 9640 15512 9646 15564
rect 9766 15512 9772 15564
rect 9824 15552 9830 15564
rect 9861 15555 9919 15561
rect 9861 15552 9873 15555
rect 9824 15524 9873 15552
rect 9824 15512 9830 15524
rect 9861 15521 9873 15524
rect 9907 15521 9919 15555
rect 9861 15515 9919 15521
rect 9950 15512 9956 15564
rect 10008 15552 10014 15564
rect 10321 15555 10379 15561
rect 10321 15552 10333 15555
rect 10008 15524 10333 15552
rect 10008 15512 10014 15524
rect 10321 15521 10333 15524
rect 10367 15521 10379 15555
rect 10321 15515 10379 15521
rect 11330 15512 11336 15564
rect 11388 15552 11394 15564
rect 11440 15561 11468 15660
rect 12250 15648 12256 15660
rect 12308 15648 12314 15700
rect 12529 15691 12587 15697
rect 12529 15657 12541 15691
rect 12575 15688 12587 15691
rect 12621 15691 12679 15697
rect 12621 15688 12633 15691
rect 12575 15660 12633 15688
rect 12575 15657 12587 15660
rect 12529 15651 12587 15657
rect 12621 15657 12633 15660
rect 12667 15688 12679 15691
rect 13170 15688 13176 15700
rect 12667 15660 13176 15688
rect 12667 15657 12679 15660
rect 12621 15651 12679 15657
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 14826 15688 14832 15700
rect 14787 15660 14832 15688
rect 14826 15648 14832 15660
rect 14884 15648 14890 15700
rect 16482 15688 16488 15700
rect 16443 15660 16488 15688
rect 16482 15648 16488 15660
rect 16540 15648 16546 15700
rect 18230 15688 18236 15700
rect 18191 15660 18236 15688
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 18598 15688 18604 15700
rect 18559 15660 18604 15688
rect 18598 15648 18604 15660
rect 18656 15648 18662 15700
rect 19518 15648 19524 15700
rect 19576 15688 19582 15700
rect 19705 15691 19763 15697
rect 19705 15688 19717 15691
rect 19576 15660 19717 15688
rect 19576 15648 19582 15660
rect 19705 15657 19717 15660
rect 19751 15657 19763 15691
rect 19705 15651 19763 15657
rect 12161 15623 12219 15629
rect 12161 15589 12173 15623
rect 12207 15620 12219 15623
rect 13078 15620 13084 15632
rect 12207 15592 13084 15620
rect 12207 15589 12219 15592
rect 12161 15583 12219 15589
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 13262 15580 13268 15632
rect 13320 15629 13326 15632
rect 13320 15623 13368 15629
rect 13320 15589 13322 15623
rect 13356 15589 13368 15623
rect 13320 15583 13368 15589
rect 13320 15580 13326 15583
rect 14734 15580 14740 15632
rect 14792 15620 14798 15632
rect 15473 15623 15531 15629
rect 15473 15620 15485 15623
rect 14792 15592 15485 15620
rect 14792 15580 14798 15592
rect 15473 15589 15485 15592
rect 15519 15620 15531 15623
rect 16758 15620 16764 15632
rect 15519 15592 16764 15620
rect 15519 15589 15531 15592
rect 15473 15583 15531 15589
rect 16758 15580 16764 15592
rect 16816 15620 16822 15632
rect 17313 15623 17371 15629
rect 17313 15620 17325 15623
rect 16816 15592 17325 15620
rect 16816 15580 16822 15592
rect 17313 15589 17325 15592
rect 17359 15589 17371 15623
rect 17313 15583 17371 15589
rect 17678 15580 17684 15632
rect 17736 15620 17742 15632
rect 17865 15623 17923 15629
rect 17865 15620 17877 15623
rect 17736 15592 17877 15620
rect 17736 15580 17742 15592
rect 17865 15589 17877 15592
rect 17911 15620 17923 15623
rect 18782 15620 18788 15632
rect 17911 15592 18788 15620
rect 17911 15589 17923 15592
rect 17865 15583 17923 15589
rect 18782 15580 18788 15592
rect 18840 15580 18846 15632
rect 18874 15580 18880 15632
rect 18932 15620 18938 15632
rect 19426 15620 19432 15632
rect 18932 15592 18977 15620
rect 19387 15592 19432 15620
rect 18932 15580 18938 15592
rect 19426 15580 19432 15592
rect 19484 15580 19490 15632
rect 21174 15620 21180 15632
rect 21135 15592 21180 15620
rect 21174 15580 21180 15592
rect 21232 15580 21238 15632
rect 21269 15623 21327 15629
rect 21269 15589 21281 15623
rect 21315 15620 21327 15623
rect 21450 15620 21456 15632
rect 21315 15592 21456 15620
rect 21315 15589 21327 15592
rect 21269 15583 21327 15589
rect 21450 15580 21456 15592
rect 21508 15580 21514 15632
rect 11425 15555 11483 15561
rect 11425 15552 11437 15555
rect 11388 15524 11437 15552
rect 11388 15512 11394 15524
rect 11425 15521 11437 15524
rect 11471 15521 11483 15555
rect 11974 15552 11980 15564
rect 11887 15524 11980 15552
rect 11425 15515 11483 15521
rect 11974 15512 11980 15524
rect 12032 15552 12038 15564
rect 12342 15552 12348 15564
rect 12032 15524 12348 15552
rect 12032 15512 12038 15524
rect 12342 15512 12348 15524
rect 12400 15512 12406 15564
rect 22716 15555 22774 15561
rect 22716 15521 22728 15555
rect 22762 15552 22774 15555
rect 22922 15552 22928 15564
rect 22762 15524 22928 15552
rect 22762 15521 22774 15524
rect 22716 15515 22774 15521
rect 22922 15512 22928 15524
rect 22980 15512 22986 15564
rect 23750 15561 23756 15564
rect 23728 15555 23756 15561
rect 23728 15552 23740 15555
rect 23663 15524 23740 15552
rect 23728 15521 23740 15524
rect 23808 15552 23814 15564
rect 23934 15552 23940 15564
rect 23808 15524 23940 15552
rect 23728 15515 23756 15521
rect 23750 15512 23756 15515
rect 23808 15512 23814 15524
rect 23934 15512 23940 15524
rect 23992 15512 23998 15564
rect 24210 15512 24216 15564
rect 24268 15552 24274 15564
rect 24740 15555 24798 15561
rect 24740 15552 24752 15555
rect 24268 15524 24752 15552
rect 24268 15512 24274 15524
rect 24740 15521 24752 15524
rect 24786 15552 24798 15555
rect 25130 15552 25136 15564
rect 24786 15524 25136 15552
rect 24786 15521 24798 15524
rect 24740 15515 24798 15521
rect 25130 15512 25136 15524
rect 25188 15512 25194 15564
rect 3602 15484 3608 15496
rect 2700 15456 3608 15484
rect 1670 15376 1676 15428
rect 1728 15416 1734 15428
rect 2700 15425 2728 15456
rect 3602 15444 3608 15456
rect 3660 15444 3666 15496
rect 10594 15484 10600 15496
rect 10555 15456 10600 15484
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 12897 15487 12955 15493
rect 12897 15484 12909 15487
rect 12308 15456 12909 15484
rect 12308 15444 12314 15456
rect 12897 15453 12909 15456
rect 12943 15484 12955 15487
rect 12989 15487 13047 15493
rect 12989 15484 13001 15487
rect 12943 15456 13001 15484
rect 12943 15453 12955 15456
rect 12897 15447 12955 15453
rect 12989 15453 13001 15456
rect 13035 15453 13047 15487
rect 15381 15487 15439 15493
rect 15381 15484 15393 15487
rect 12989 15447 13047 15453
rect 15304 15456 15393 15484
rect 15304 15428 15332 15456
rect 15381 15453 15393 15456
rect 15427 15453 15439 15487
rect 15381 15447 15439 15453
rect 15470 15444 15476 15496
rect 15528 15484 15534 15496
rect 15657 15487 15715 15493
rect 15657 15484 15669 15487
rect 15528 15456 15669 15484
rect 15528 15444 15534 15456
rect 15657 15453 15669 15456
rect 15703 15453 15715 15487
rect 17218 15484 17224 15496
rect 17179 15456 17224 15484
rect 15657 15447 15715 15453
rect 17218 15444 17224 15456
rect 17276 15444 17282 15496
rect 18598 15444 18604 15496
rect 18656 15484 18662 15496
rect 18785 15487 18843 15493
rect 18785 15484 18797 15487
rect 18656 15456 18797 15484
rect 18656 15444 18662 15456
rect 18785 15453 18797 15456
rect 18831 15453 18843 15487
rect 18785 15447 18843 15453
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 22278 15484 22284 15496
rect 22152 15456 22284 15484
rect 22152 15444 22158 15456
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 2685 15419 2743 15425
rect 2685 15416 2697 15419
rect 1728 15388 2697 15416
rect 1728 15376 1734 15388
rect 2685 15385 2697 15388
rect 2731 15385 2743 15419
rect 2685 15379 2743 15385
rect 2866 15376 2872 15428
rect 2924 15416 2930 15428
rect 3145 15419 3203 15425
rect 3145 15416 3157 15419
rect 2924 15388 3157 15416
rect 2924 15376 2930 15388
rect 3145 15385 3157 15388
rect 3191 15416 3203 15419
rect 3694 15416 3700 15428
rect 3191 15388 3700 15416
rect 3191 15385 3203 15388
rect 3145 15379 3203 15385
rect 3694 15376 3700 15388
rect 3752 15376 3758 15428
rect 15286 15376 15292 15428
rect 15344 15376 15350 15428
rect 21726 15416 21732 15428
rect 21687 15388 21732 15416
rect 21726 15376 21732 15388
rect 21784 15376 21790 15428
rect 1302 15308 1308 15360
rect 1360 15348 1366 15360
rect 1949 15351 2007 15357
rect 1949 15348 1961 15351
rect 1360 15320 1961 15348
rect 1360 15308 1366 15320
rect 1949 15317 1961 15320
rect 1995 15348 2007 15351
rect 2130 15348 2136 15360
rect 1995 15320 2136 15348
rect 1995 15317 2007 15320
rect 1949 15311 2007 15317
rect 2130 15308 2136 15320
rect 2188 15308 2194 15360
rect 3602 15348 3608 15360
rect 3563 15320 3608 15348
rect 3602 15308 3608 15320
rect 3660 15308 3666 15360
rect 4338 15308 4344 15360
rect 4396 15348 4402 15360
rect 4617 15351 4675 15357
rect 4617 15348 4629 15351
rect 4396 15320 4629 15348
rect 4396 15308 4402 15320
rect 4617 15317 4629 15320
rect 4663 15317 4675 15351
rect 6362 15348 6368 15360
rect 6323 15320 6368 15348
rect 4617 15311 4675 15317
rect 6362 15308 6368 15320
rect 6420 15308 6426 15360
rect 7742 15308 7748 15360
rect 7800 15348 7806 15360
rect 7837 15351 7895 15357
rect 7837 15348 7849 15351
rect 7800 15320 7849 15348
rect 7800 15308 7806 15320
rect 7837 15317 7849 15320
rect 7883 15348 7895 15351
rect 8202 15348 8208 15360
rect 7883 15320 8208 15348
rect 7883 15317 7895 15320
rect 7837 15311 7895 15317
rect 8202 15308 8208 15320
rect 8260 15308 8266 15360
rect 12342 15308 12348 15360
rect 12400 15348 12406 15360
rect 12621 15351 12679 15357
rect 12621 15348 12633 15351
rect 12400 15320 12633 15348
rect 12400 15308 12406 15320
rect 12621 15317 12633 15320
rect 12667 15317 12679 15351
rect 12621 15311 12679 15317
rect 13909 15351 13967 15357
rect 13909 15317 13921 15351
rect 13955 15348 13967 15351
rect 14734 15348 14740 15360
rect 13955 15320 14740 15348
rect 13955 15317 13967 15320
rect 13909 15311 13967 15317
rect 14734 15308 14740 15320
rect 14792 15308 14798 15360
rect 22462 15308 22468 15360
rect 22520 15348 22526 15360
rect 22787 15351 22845 15357
rect 22787 15348 22799 15351
rect 22520 15320 22799 15348
rect 22520 15308 22526 15320
rect 22787 15317 22799 15320
rect 22833 15317 22845 15351
rect 22787 15311 22845 15317
rect 23474 15308 23480 15360
rect 23532 15348 23538 15360
rect 23799 15351 23857 15357
rect 23799 15348 23811 15351
rect 23532 15320 23811 15348
rect 23532 15308 23538 15320
rect 23799 15317 23811 15320
rect 23845 15317 23857 15351
rect 23799 15311 23857 15317
rect 24811 15351 24869 15357
rect 24811 15317 24823 15351
rect 24857 15348 24869 15351
rect 25222 15348 25228 15360
rect 24857 15320 25228 15348
rect 24857 15317 24869 15320
rect 24811 15311 24869 15317
rect 25222 15308 25228 15320
rect 25280 15308 25286 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1946 15144 1952 15156
rect 1907 15116 1952 15144
rect 1946 15104 1952 15116
rect 2004 15104 2010 15156
rect 2406 15144 2412 15156
rect 2367 15116 2412 15144
rect 2406 15104 2412 15116
rect 2464 15104 2470 15156
rect 4614 15144 4620 15156
rect 4575 15116 4620 15144
rect 4614 15104 4620 15116
rect 4672 15144 4678 15156
rect 4672 15116 5580 15144
rect 4672 15104 4678 15116
rect 1765 15079 1823 15085
rect 1765 15045 1777 15079
rect 1811 15045 1823 15079
rect 5074 15076 5080 15088
rect 1765 15039 1823 15045
rect 3896 15048 5080 15076
rect 1780 15008 1808 15039
rect 1780 14980 2360 15008
rect 2332 14952 2360 14980
rect 1581 14943 1639 14949
rect 1581 14909 1593 14943
rect 1627 14909 1639 14943
rect 1581 14903 1639 14909
rect 1596 14872 1624 14903
rect 2314 14900 2320 14952
rect 2372 14900 2378 14952
rect 2660 14943 2718 14949
rect 2660 14909 2672 14943
rect 2706 14940 2718 14943
rect 3142 14940 3148 14952
rect 2706 14912 3148 14940
rect 2706 14909 2718 14912
rect 2660 14903 2718 14909
rect 3142 14900 3148 14912
rect 3200 14900 3206 14952
rect 3694 14900 3700 14952
rect 3752 14940 3758 14952
rect 3896 14949 3924 15048
rect 5074 15036 5080 15048
rect 5132 15036 5138 15088
rect 4338 15008 4344 15020
rect 4299 14980 4344 15008
rect 4338 14968 4344 14980
rect 4396 14968 4402 15020
rect 3881 14943 3939 14949
rect 3881 14940 3893 14943
rect 3752 14912 3893 14940
rect 3752 14900 3758 14912
rect 3881 14909 3893 14912
rect 3927 14909 3939 14943
rect 4154 14940 4160 14952
rect 4115 14912 4160 14940
rect 3881 14903 3939 14909
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 5074 14900 5080 14952
rect 5132 14940 5138 14952
rect 5169 14943 5227 14949
rect 5169 14940 5181 14943
rect 5132 14912 5181 14940
rect 5132 14900 5138 14912
rect 5169 14909 5181 14912
rect 5215 14909 5227 14943
rect 5552 14940 5580 15116
rect 7006 15104 7012 15156
rect 7064 15144 7070 15156
rect 8021 15147 8079 15153
rect 8021 15144 8033 15147
rect 7064 15116 8033 15144
rect 7064 15104 7070 15116
rect 8021 15113 8033 15116
rect 8067 15113 8079 15147
rect 8021 15107 8079 15113
rect 9766 15104 9772 15156
rect 9824 15144 9830 15156
rect 9861 15147 9919 15153
rect 9861 15144 9873 15147
rect 9824 15116 9873 15144
rect 9824 15104 9830 15116
rect 9861 15113 9873 15116
rect 9907 15144 9919 15147
rect 10597 15147 10655 15153
rect 10597 15144 10609 15147
rect 9907 15116 10609 15144
rect 9907 15113 9919 15116
rect 9861 15107 9919 15113
rect 10597 15113 10609 15116
rect 10643 15144 10655 15147
rect 11422 15144 11428 15156
rect 10643 15116 11428 15144
rect 10643 15113 10655 15116
rect 10597 15107 10655 15113
rect 9950 15036 9956 15088
rect 10008 15076 10014 15088
rect 10229 15079 10287 15085
rect 10229 15076 10241 15079
rect 10008 15048 10241 15076
rect 10008 15036 10014 15048
rect 10229 15045 10241 15048
rect 10275 15045 10287 15079
rect 10229 15039 10287 15045
rect 5905 15011 5963 15017
rect 5905 14977 5917 15011
rect 5951 15008 5963 15011
rect 6362 15008 6368 15020
rect 5951 14980 6368 15008
rect 5951 14977 5963 14980
rect 5905 14971 5963 14977
rect 6362 14968 6368 14980
rect 6420 15008 6426 15020
rect 6825 15011 6883 15017
rect 6825 15008 6837 15011
rect 6420 14980 6837 15008
rect 6420 14968 6426 14980
rect 6825 14977 6837 14980
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 8662 14968 8668 15020
rect 8720 15008 8726 15020
rect 8941 15011 8999 15017
rect 8941 15008 8953 15011
rect 8720 14980 8953 15008
rect 8720 14968 8726 14980
rect 8941 14977 8953 14980
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 5629 14943 5687 14949
rect 5629 14940 5641 14943
rect 5552 14912 5641 14940
rect 5169 14903 5227 14909
rect 5629 14909 5641 14912
rect 5675 14940 5687 14943
rect 7006 14940 7012 14952
rect 5675 14912 7012 14940
rect 5675 14909 5687 14912
rect 5629 14903 5687 14909
rect 7006 14900 7012 14912
rect 7064 14900 7070 14952
rect 10612 14940 10640 15107
rect 11422 15104 11428 15116
rect 11480 15104 11486 15156
rect 11974 15104 11980 15156
rect 12032 15144 12038 15156
rect 12161 15147 12219 15153
rect 12161 15144 12173 15147
rect 12032 15116 12173 15144
rect 12032 15104 12038 15116
rect 12161 15113 12173 15116
rect 12207 15113 12219 15147
rect 12161 15107 12219 15113
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 12575 15147 12633 15153
rect 12575 15144 12587 15147
rect 12492 15116 12587 15144
rect 12492 15104 12498 15116
rect 12575 15113 12587 15116
rect 12621 15113 12633 15147
rect 12575 15107 12633 15113
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 12897 15147 12955 15153
rect 12897 15144 12909 15147
rect 12768 15116 12909 15144
rect 12768 15104 12774 15116
rect 12897 15113 12909 15116
rect 12943 15113 12955 15147
rect 14734 15144 14740 15156
rect 14695 15116 14740 15144
rect 12897 15107 12955 15113
rect 14734 15104 14740 15116
rect 14792 15104 14798 15156
rect 16758 15144 16764 15156
rect 16719 15116 16764 15144
rect 16758 15104 16764 15116
rect 16816 15144 16822 15156
rect 18874 15144 18880 15156
rect 16816 15116 18880 15144
rect 16816 15104 16822 15116
rect 18874 15104 18880 15116
rect 18932 15144 18938 15156
rect 19061 15147 19119 15153
rect 19061 15144 19073 15147
rect 18932 15116 19073 15144
rect 18932 15104 18938 15116
rect 19061 15113 19073 15116
rect 19107 15113 19119 15147
rect 19061 15107 19119 15113
rect 21174 15104 21180 15156
rect 21232 15144 21238 15156
rect 21729 15147 21787 15153
rect 21729 15144 21741 15147
rect 21232 15116 21741 15144
rect 21232 15104 21238 15116
rect 21729 15113 21741 15116
rect 21775 15113 21787 15147
rect 21729 15107 21787 15113
rect 22833 15147 22891 15153
rect 22833 15113 22845 15147
rect 22879 15144 22891 15147
rect 22922 15144 22928 15156
rect 22879 15116 22928 15144
rect 22879 15113 22891 15116
rect 22833 15107 22891 15113
rect 22922 15104 22928 15116
rect 22980 15104 22986 15156
rect 15930 15076 15936 15088
rect 15891 15048 15936 15076
rect 15930 15036 15936 15048
rect 15988 15036 15994 15088
rect 16574 15036 16580 15088
rect 16632 15076 16638 15088
rect 17681 15079 17739 15085
rect 17681 15076 17693 15079
rect 16632 15048 17693 15076
rect 16632 15036 16638 15048
rect 17681 15045 17693 15048
rect 17727 15076 17739 15079
rect 17773 15079 17831 15085
rect 17773 15076 17785 15079
rect 17727 15048 17785 15076
rect 17727 15045 17739 15048
rect 17681 15039 17739 15045
rect 17773 15045 17785 15048
rect 17819 15045 17831 15079
rect 17773 15039 17831 15045
rect 11517 15011 11575 15017
rect 11517 14977 11529 15011
rect 11563 15008 11575 15011
rect 12342 15008 12348 15020
rect 11563 14980 12348 15008
rect 11563 14977 11575 14980
rect 11517 14971 11575 14977
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 13817 15011 13875 15017
rect 13817 14977 13829 15011
rect 13863 15008 13875 15011
rect 13906 15008 13912 15020
rect 13863 14980 13912 15008
rect 13863 14977 13875 14980
rect 13817 14971 13875 14977
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 14090 15008 14096 15020
rect 14051 14980 14096 15008
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 15008 15439 15011
rect 16390 15008 16396 15020
rect 15427 14980 16396 15008
rect 15427 14977 15439 14980
rect 15381 14971 15439 14977
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 17126 14968 17132 15020
rect 17184 15008 17190 15020
rect 17405 15011 17463 15017
rect 17405 15008 17417 15011
rect 17184 14980 17417 15008
rect 17184 14968 17190 14980
rect 17405 14977 17417 14980
rect 17451 14977 17463 15011
rect 17405 14971 17463 14977
rect 18141 15011 18199 15017
rect 18141 14977 18153 15011
rect 18187 15008 18199 15011
rect 18230 15008 18236 15020
rect 18187 14980 18236 15008
rect 18187 14977 18199 14980
rect 18141 14971 18199 14977
rect 18230 14968 18236 14980
rect 18288 14968 18294 15020
rect 18782 15008 18788 15020
rect 18743 14980 18788 15008
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 22097 15011 22155 15017
rect 22097 15008 22109 15011
rect 21468 14980 22109 15008
rect 10781 14943 10839 14949
rect 10781 14940 10793 14943
rect 10612 14912 10793 14940
rect 10781 14909 10793 14912
rect 10827 14909 10839 14943
rect 11330 14940 11336 14952
rect 11243 14912 11336 14940
rect 10781 14903 10839 14909
rect 11330 14900 11336 14912
rect 11388 14940 11394 14952
rect 11974 14940 11980 14952
rect 11388 14912 11980 14940
rect 11388 14900 11394 14912
rect 11974 14900 11980 14912
rect 12032 14900 12038 14952
rect 12504 14943 12562 14949
rect 12504 14909 12516 14943
rect 12550 14940 12562 14943
rect 12710 14940 12716 14952
rect 12550 14912 12716 14940
rect 12550 14909 12562 14912
rect 12504 14903 12562 14909
rect 12710 14900 12716 14912
rect 12768 14900 12774 14952
rect 16298 14900 16304 14952
rect 16356 14940 16362 14952
rect 16996 14943 17054 14949
rect 16996 14940 17008 14943
rect 16356 14912 17008 14940
rect 16356 14900 16362 14912
rect 16996 14909 17008 14912
rect 17042 14940 17054 14943
rect 17144 14940 17172 14968
rect 21468 14952 21496 14980
rect 22097 14977 22109 14980
rect 22143 14977 22155 15011
rect 22097 14971 22155 14977
rect 20530 14940 20536 14952
rect 17042 14912 17172 14940
rect 20491 14912 20536 14940
rect 17042 14909 17054 14912
rect 16996 14903 17054 14909
rect 20530 14900 20536 14912
rect 20588 14900 20594 14952
rect 21450 14940 21456 14952
rect 21411 14912 21456 14940
rect 21450 14900 21456 14912
rect 21508 14900 21514 14952
rect 21634 14900 21640 14952
rect 21692 14940 21698 14952
rect 22332 14943 22390 14949
rect 22332 14940 22344 14943
rect 21692 14912 22344 14940
rect 21692 14900 21698 14912
rect 22332 14909 22344 14912
rect 22378 14940 22390 14943
rect 23109 14943 23167 14949
rect 23109 14940 23121 14943
rect 22378 14912 23121 14940
rect 22378 14909 22390 14912
rect 22332 14903 22390 14909
rect 23109 14909 23121 14912
rect 23155 14909 23167 14943
rect 23109 14903 23167 14909
rect 23728 14943 23786 14949
rect 23728 14909 23740 14943
rect 23774 14940 23786 14943
rect 24026 14940 24032 14952
rect 23774 14912 24032 14940
rect 23774 14909 23786 14912
rect 23728 14903 23786 14909
rect 24026 14900 24032 14912
rect 24084 14940 24090 14952
rect 24121 14943 24179 14949
rect 24121 14940 24133 14943
rect 24084 14912 24133 14940
rect 24084 14900 24090 14912
rect 24121 14909 24133 14912
rect 24167 14909 24179 14943
rect 24121 14903 24179 14909
rect 1949 14875 2007 14881
rect 1949 14872 1961 14875
rect 1596 14844 1961 14872
rect 1949 14841 1961 14844
rect 1995 14872 2007 14875
rect 2041 14875 2099 14881
rect 2041 14872 2053 14875
rect 1995 14844 2053 14872
rect 1995 14841 2007 14844
rect 1949 14835 2007 14841
rect 2041 14841 2053 14844
rect 2087 14872 2099 14875
rect 2087 14844 2912 14872
rect 2087 14841 2099 14844
rect 2041 14835 2099 14841
rect 2130 14764 2136 14816
rect 2188 14804 2194 14816
rect 2731 14807 2789 14813
rect 2731 14804 2743 14807
rect 2188 14776 2743 14804
rect 2188 14764 2194 14776
rect 2731 14773 2743 14776
rect 2777 14773 2789 14807
rect 2884 14804 2912 14844
rect 2958 14832 2964 14884
rect 3016 14872 3022 14884
rect 3513 14875 3571 14881
rect 3513 14872 3525 14875
rect 3016 14844 3525 14872
rect 3016 14832 3022 14844
rect 3513 14841 3525 14844
rect 3559 14872 3571 14875
rect 6822 14872 6828 14884
rect 3559 14844 5120 14872
rect 3559 14841 3571 14844
rect 3513 14835 3571 14841
rect 4338 14804 4344 14816
rect 2884 14776 4344 14804
rect 2731 14767 2789 14773
rect 4338 14764 4344 14776
rect 4396 14764 4402 14816
rect 5092 14813 5120 14844
rect 6564 14844 6828 14872
rect 6564 14816 6592 14844
rect 6822 14832 6828 14844
rect 6880 14872 6886 14884
rect 7146 14875 7204 14881
rect 7146 14872 7158 14875
rect 6880 14844 7158 14872
rect 6880 14832 6886 14844
rect 7146 14841 7158 14844
rect 7192 14841 7204 14875
rect 8662 14872 8668 14884
rect 8623 14844 8668 14872
rect 7146 14835 7204 14841
rect 8662 14832 8668 14844
rect 8720 14832 8726 14884
rect 8754 14832 8760 14884
rect 8812 14872 8818 14884
rect 8812 14844 8857 14872
rect 8812 14832 8818 14844
rect 11422 14832 11428 14884
rect 11480 14872 11486 14884
rect 11793 14875 11851 14881
rect 11793 14872 11805 14875
rect 11480 14844 11805 14872
rect 11480 14832 11486 14844
rect 11793 14841 11805 14844
rect 11839 14841 11851 14875
rect 11793 14835 11851 14841
rect 13906 14832 13912 14884
rect 13964 14872 13970 14884
rect 15197 14875 15255 14881
rect 13964 14844 14009 14872
rect 13964 14832 13970 14844
rect 15197 14841 15209 14875
rect 15243 14872 15255 14875
rect 15378 14872 15384 14884
rect 15243 14844 15384 14872
rect 15243 14841 15255 14844
rect 15197 14835 15255 14841
rect 15378 14832 15384 14844
rect 15436 14872 15442 14884
rect 15473 14875 15531 14881
rect 15473 14872 15485 14875
rect 15436 14844 15485 14872
rect 15436 14832 15442 14844
rect 15473 14841 15485 14844
rect 15519 14841 15531 14875
rect 15473 14835 15531 14841
rect 17083 14875 17141 14881
rect 17083 14841 17095 14875
rect 17129 14872 17141 14875
rect 17954 14872 17960 14884
rect 17129 14844 17960 14872
rect 17129 14841 17141 14844
rect 17083 14835 17141 14841
rect 17954 14832 17960 14844
rect 18012 14832 18018 14884
rect 18233 14875 18291 14881
rect 18233 14841 18245 14875
rect 18279 14872 18291 14875
rect 19242 14872 19248 14884
rect 18279 14844 19248 14872
rect 18279 14841 18291 14844
rect 18233 14835 18291 14841
rect 5077 14807 5135 14813
rect 5077 14773 5089 14807
rect 5123 14804 5135 14807
rect 5166 14804 5172 14816
rect 5123 14776 5172 14804
rect 5123 14773 5135 14776
rect 5077 14767 5135 14773
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 6273 14807 6331 14813
rect 6273 14773 6285 14807
rect 6319 14804 6331 14807
rect 6546 14804 6552 14816
rect 6319 14776 6552 14804
rect 6319 14773 6331 14776
rect 6273 14767 6331 14773
rect 6546 14764 6552 14776
rect 6604 14764 6610 14816
rect 7742 14804 7748 14816
rect 7703 14776 7748 14804
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 8478 14804 8484 14816
rect 8439 14776 8484 14804
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 12710 14764 12716 14816
rect 12768 14804 12774 14816
rect 12894 14804 12900 14816
rect 12768 14776 12900 14804
rect 12768 14764 12774 14776
rect 12894 14764 12900 14776
rect 12952 14764 12958 14816
rect 13078 14764 13084 14816
rect 13136 14804 13142 14816
rect 13262 14804 13268 14816
rect 13136 14776 13268 14804
rect 13136 14764 13142 14776
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 17681 14807 17739 14813
rect 17681 14773 17693 14807
rect 17727 14804 17739 14807
rect 18248 14804 18276 14835
rect 19242 14832 19248 14844
rect 19300 14832 19306 14884
rect 20854 14875 20912 14881
rect 20854 14872 20866 14875
rect 20364 14844 20866 14872
rect 17727 14776 18276 14804
rect 17727 14773 17739 14776
rect 17681 14767 17739 14773
rect 19334 14764 19340 14816
rect 19392 14804 19398 14816
rect 19429 14807 19487 14813
rect 19429 14804 19441 14807
rect 19392 14776 19441 14804
rect 19392 14764 19398 14776
rect 19429 14773 19441 14776
rect 19475 14773 19487 14807
rect 19429 14767 19487 14773
rect 19518 14764 19524 14816
rect 19576 14804 19582 14816
rect 20364 14813 20392 14844
rect 20854 14841 20866 14844
rect 20900 14841 20912 14875
rect 20854 14835 20912 14841
rect 23566 14832 23572 14884
rect 23624 14872 23630 14884
rect 24673 14875 24731 14881
rect 24673 14872 24685 14875
rect 23624 14844 24685 14872
rect 23624 14832 23630 14844
rect 24673 14841 24685 14844
rect 24719 14841 24731 14875
rect 24673 14835 24731 14841
rect 20349 14807 20407 14813
rect 20349 14804 20361 14807
rect 19576 14776 20361 14804
rect 19576 14764 19582 14776
rect 20349 14773 20361 14776
rect 20395 14773 20407 14807
rect 20349 14767 20407 14773
rect 20990 14764 20996 14816
rect 21048 14804 21054 14816
rect 22419 14807 22477 14813
rect 22419 14804 22431 14807
rect 21048 14776 22431 14804
rect 21048 14764 21054 14776
rect 22419 14773 22431 14776
rect 22465 14773 22477 14807
rect 22419 14767 22477 14773
rect 23474 14764 23480 14816
rect 23532 14804 23538 14816
rect 23799 14807 23857 14813
rect 23799 14804 23811 14807
rect 23532 14776 23811 14804
rect 23532 14764 23538 14776
rect 23799 14773 23811 14776
rect 23845 14773 23857 14807
rect 23799 14767 23857 14773
rect 23934 14764 23940 14816
rect 23992 14804 23998 14816
rect 24489 14807 24547 14813
rect 24489 14804 24501 14807
rect 23992 14776 24501 14804
rect 23992 14764 23998 14776
rect 24489 14773 24501 14776
rect 24535 14773 24547 14807
rect 25130 14804 25136 14816
rect 25091 14776 25136 14804
rect 24489 14767 24547 14773
rect 25130 14764 25136 14776
rect 25188 14764 25194 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 3142 14609 3148 14612
rect 3099 14603 3148 14609
rect 3099 14569 3111 14603
rect 3145 14569 3148 14603
rect 3099 14563 3148 14569
rect 3142 14560 3148 14563
rect 3200 14560 3206 14612
rect 3326 14560 3332 14612
rect 3384 14600 3390 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 3384 14572 4169 14600
rect 3384 14560 3390 14572
rect 4157 14569 4169 14572
rect 4203 14569 4215 14603
rect 4157 14563 4215 14569
rect 5074 14560 5080 14612
rect 5132 14600 5138 14612
rect 5169 14603 5227 14609
rect 5169 14600 5181 14603
rect 5132 14572 5181 14600
rect 5132 14560 5138 14572
rect 5169 14569 5181 14572
rect 5215 14569 5227 14603
rect 5169 14563 5227 14569
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 5537 14603 5595 14609
rect 5537 14600 5549 14603
rect 5316 14572 5549 14600
rect 5316 14560 5322 14572
rect 5537 14569 5549 14572
rect 5583 14569 5595 14603
rect 5537 14563 5595 14569
rect 8662 14560 8668 14612
rect 8720 14600 8726 14612
rect 8941 14603 8999 14609
rect 8941 14600 8953 14603
rect 8720 14572 8953 14600
rect 8720 14560 8726 14572
rect 8941 14569 8953 14572
rect 8987 14569 8999 14603
rect 9950 14600 9956 14612
rect 9911 14572 9956 14600
rect 8941 14563 8999 14569
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 10873 14603 10931 14609
rect 10873 14569 10885 14603
rect 10919 14600 10931 14603
rect 11330 14600 11336 14612
rect 10919 14572 11336 14600
rect 10919 14569 10931 14572
rect 10873 14563 10931 14569
rect 11330 14560 11336 14572
rect 11388 14560 11394 14612
rect 13814 14600 13820 14612
rect 13775 14572 13820 14600
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 17218 14600 17224 14612
rect 17179 14572 17224 14600
rect 17218 14560 17224 14572
rect 17276 14560 17282 14612
rect 17862 14600 17868 14612
rect 17604 14572 17868 14600
rect 3694 14532 3700 14544
rect 3655 14504 3700 14532
rect 3694 14492 3700 14504
rect 3752 14492 3758 14544
rect 4062 14492 4068 14544
rect 4120 14532 4126 14544
rect 7742 14532 7748 14544
rect 4120 14504 6316 14532
rect 7703 14504 7748 14532
rect 4120 14492 4126 14504
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 1578 14464 1584 14476
rect 1443 14436 1584 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 1578 14424 1584 14436
rect 1636 14424 1642 14476
rect 3028 14467 3086 14473
rect 3028 14433 3040 14467
rect 3074 14464 3086 14467
rect 3142 14464 3148 14476
rect 3074 14436 3148 14464
rect 3074 14433 3086 14436
rect 3028 14427 3086 14433
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 3602 14424 3608 14476
rect 3660 14464 3666 14476
rect 4154 14464 4160 14476
rect 3660 14436 4160 14464
rect 3660 14424 3666 14436
rect 4154 14424 4160 14436
rect 4212 14424 4218 14476
rect 4632 14473 4660 14504
rect 6288 14476 6316 14504
rect 7742 14492 7748 14504
rect 7800 14532 7806 14544
rect 8110 14532 8116 14544
rect 7800 14504 8116 14532
rect 7800 14492 7806 14504
rect 8110 14492 8116 14504
rect 8168 14532 8174 14544
rect 8573 14535 8631 14541
rect 8573 14532 8585 14535
rect 8168 14504 8585 14532
rect 8168 14492 8174 14504
rect 8573 14501 8585 14504
rect 8619 14532 8631 14535
rect 8754 14532 8760 14544
rect 8619 14504 8760 14532
rect 8619 14501 8631 14504
rect 8573 14495 8631 14501
rect 8754 14492 8760 14504
rect 8812 14492 8818 14544
rect 4617 14467 4675 14473
rect 4617 14433 4629 14467
rect 4663 14433 4675 14467
rect 4617 14427 4675 14433
rect 6089 14467 6147 14473
rect 6089 14433 6101 14467
rect 6135 14433 6147 14467
rect 6270 14464 6276 14476
rect 6231 14436 6276 14464
rect 6089 14427 6147 14433
rect 6104 14396 6132 14427
rect 6270 14424 6276 14436
rect 6328 14424 6334 14476
rect 9766 14464 9772 14476
rect 9727 14436 9772 14464
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 10137 14467 10195 14473
rect 10137 14433 10149 14467
rect 10183 14433 10195 14467
rect 10137 14427 10195 14433
rect 6178 14396 6184 14408
rect 6104 14368 6184 14396
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 6362 14396 6368 14408
rect 6323 14368 6368 14396
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 7653 14399 7711 14405
rect 7653 14365 7665 14399
rect 7699 14396 7711 14399
rect 7926 14396 7932 14408
rect 7699 14368 7932 14396
rect 7699 14365 7711 14368
rect 7653 14359 7711 14365
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 8018 14356 8024 14408
rect 8076 14396 8082 14408
rect 8076 14368 8121 14396
rect 8076 14356 8082 14368
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 10152 14396 10180 14427
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 11241 14467 11299 14473
rect 11241 14464 11253 14467
rect 11112 14436 11253 14464
rect 11112 14424 11118 14436
rect 11241 14433 11253 14436
rect 11287 14433 11299 14467
rect 11348 14464 11376 14560
rect 11977 14535 12035 14541
rect 11977 14501 11989 14535
rect 12023 14532 12035 14535
rect 12250 14532 12256 14544
rect 12023 14504 12256 14532
rect 12023 14501 12035 14504
rect 11977 14495 12035 14501
rect 12250 14492 12256 14504
rect 12308 14492 12314 14544
rect 12986 14532 12992 14544
rect 12947 14504 12992 14532
rect 12986 14492 12992 14504
rect 13044 14492 13050 14544
rect 13541 14535 13599 14541
rect 13541 14501 13553 14535
rect 13587 14532 13599 14535
rect 14090 14532 14096 14544
rect 13587 14504 14096 14532
rect 13587 14501 13599 14504
rect 13541 14495 13599 14501
rect 14090 14492 14096 14504
rect 14148 14492 14154 14544
rect 15473 14535 15531 14541
rect 15473 14532 15485 14535
rect 14200 14504 15485 14532
rect 11698 14464 11704 14476
rect 11348 14436 11704 14464
rect 11241 14427 11299 14433
rect 9640 14368 10180 14396
rect 11256 14396 11284 14427
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 11790 14396 11796 14408
rect 11256 14368 11796 14396
rect 9640 14356 9646 14368
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 12066 14356 12072 14408
rect 12124 14396 12130 14408
rect 12894 14396 12900 14408
rect 12124 14368 12900 14396
rect 12124 14356 12130 14368
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14200 14405 14228 14504
rect 15473 14501 15485 14504
rect 15519 14501 15531 14535
rect 15473 14495 15531 14501
rect 17402 14492 17408 14544
rect 17460 14532 17466 14544
rect 17604 14541 17632 14572
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 20530 14560 20536 14612
rect 20588 14600 20594 14612
rect 20625 14603 20683 14609
rect 20625 14600 20637 14603
rect 20588 14572 20637 14600
rect 20588 14560 20594 14572
rect 20625 14569 20637 14572
rect 20671 14600 20683 14603
rect 22557 14603 22615 14609
rect 22557 14600 22569 14603
rect 20671 14572 22569 14600
rect 20671 14569 20683 14572
rect 20625 14563 20683 14569
rect 22557 14569 22569 14572
rect 22603 14569 22615 14603
rect 24762 14600 24768 14612
rect 24723 14572 24768 14600
rect 22557 14563 22615 14569
rect 24762 14560 24768 14572
rect 24820 14560 24826 14612
rect 17589 14535 17647 14541
rect 17589 14532 17601 14535
rect 17460 14504 17601 14532
rect 17460 14492 17466 14504
rect 17589 14501 17601 14504
rect 17635 14501 17647 14535
rect 17589 14495 17647 14501
rect 17681 14535 17739 14541
rect 17681 14501 17693 14535
rect 17727 14532 17739 14535
rect 18046 14532 18052 14544
rect 17727 14504 18052 14532
rect 17727 14501 17739 14504
rect 17681 14495 17739 14501
rect 18046 14492 18052 14504
rect 18104 14492 18110 14544
rect 18966 14492 18972 14544
rect 19024 14532 19030 14544
rect 19382 14535 19440 14541
rect 19382 14532 19394 14535
rect 19024 14504 19394 14532
rect 19024 14492 19030 14504
rect 19382 14501 19394 14504
rect 19428 14532 19440 14535
rect 19518 14532 19524 14544
rect 19428 14504 19524 14532
rect 19428 14501 19440 14504
rect 19382 14495 19440 14501
rect 19518 14492 19524 14504
rect 19576 14492 19582 14544
rect 20162 14532 20168 14544
rect 19996 14504 20168 14532
rect 19996 14473 20024 14504
rect 20162 14492 20168 14504
rect 20220 14532 20226 14544
rect 21082 14532 21088 14544
rect 20220 14504 21088 14532
rect 20220 14492 20226 14504
rect 21082 14492 21088 14504
rect 21140 14492 21146 14544
rect 19981 14467 20039 14473
rect 19981 14433 19993 14467
rect 20027 14433 20039 14467
rect 22738 14464 22744 14476
rect 22699 14436 22744 14464
rect 19981 14427 20039 14433
rect 22738 14424 22744 14436
rect 22796 14424 22802 14476
rect 22922 14464 22928 14476
rect 22883 14436 22928 14464
rect 22922 14424 22928 14436
rect 22980 14424 22986 14476
rect 24581 14467 24639 14473
rect 24581 14433 24593 14467
rect 24627 14464 24639 14467
rect 24670 14464 24676 14476
rect 24627 14436 24676 14464
rect 24627 14433 24639 14436
rect 24581 14427 24639 14433
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 14185 14399 14243 14405
rect 14185 14396 14197 14399
rect 13872 14368 14197 14396
rect 13872 14356 13878 14368
rect 14185 14365 14197 14368
rect 14231 14365 14243 14399
rect 14185 14359 14243 14365
rect 14826 14356 14832 14408
rect 14884 14396 14890 14408
rect 15381 14399 15439 14405
rect 15381 14396 15393 14399
rect 14884 14368 15393 14396
rect 14884 14356 14890 14368
rect 15381 14365 15393 14368
rect 15427 14396 15439 14399
rect 15470 14396 15476 14408
rect 15427 14368 15476 14396
rect 15427 14365 15439 14368
rect 15381 14359 15439 14365
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 16022 14396 16028 14408
rect 15983 14368 16028 14396
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 18233 14399 18291 14405
rect 18233 14365 18245 14399
rect 18279 14396 18291 14399
rect 18782 14396 18788 14408
rect 18279 14368 18788 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 18782 14356 18788 14368
rect 18840 14356 18846 14408
rect 19061 14399 19119 14405
rect 19061 14365 19073 14399
rect 19107 14396 19119 14399
rect 19242 14396 19248 14408
rect 19107 14368 19248 14396
rect 19107 14365 19119 14368
rect 19061 14359 19119 14365
rect 19242 14356 19248 14368
rect 19300 14356 19306 14408
rect 20990 14396 20996 14408
rect 20951 14368 20996 14396
rect 20990 14356 20996 14368
rect 21048 14356 21054 14408
rect 21450 14396 21456 14408
rect 21411 14368 21456 14396
rect 21450 14356 21456 14368
rect 21508 14356 21514 14408
rect 3050 14288 3056 14340
rect 3108 14328 3114 14340
rect 3694 14328 3700 14340
rect 3108 14300 3700 14328
rect 3108 14288 3114 14300
rect 3694 14288 3700 14300
rect 3752 14288 3758 14340
rect 13538 14288 13544 14340
rect 13596 14328 13602 14340
rect 15013 14331 15071 14337
rect 15013 14328 15025 14331
rect 13596 14300 15025 14328
rect 13596 14288 13602 14300
rect 15013 14297 15025 14300
rect 15059 14328 15071 14331
rect 15286 14328 15292 14340
rect 15059 14300 15292 14328
rect 15059 14297 15071 14300
rect 15013 14291 15071 14297
rect 15286 14288 15292 14300
rect 15344 14288 15350 14340
rect 7193 14263 7251 14269
rect 7193 14229 7205 14263
rect 7239 14260 7251 14263
rect 7282 14260 7288 14272
rect 7239 14232 7288 14260
rect 7239 14229 7251 14232
rect 7193 14223 7251 14229
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 9493 14263 9551 14269
rect 9493 14229 9505 14263
rect 9539 14260 9551 14263
rect 10134 14260 10140 14272
rect 9539 14232 10140 14260
rect 9539 14229 9551 14232
rect 9493 14223 9551 14229
rect 10134 14220 10140 14232
rect 10192 14220 10198 14272
rect 21634 14220 21640 14272
rect 21692 14260 21698 14272
rect 21913 14263 21971 14269
rect 21913 14260 21925 14263
rect 21692 14232 21925 14260
rect 21692 14220 21698 14232
rect 21913 14229 21925 14232
rect 21959 14229 21971 14263
rect 22278 14260 22284 14272
rect 22239 14232 22284 14260
rect 21913 14223 21971 14229
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 23750 14260 23756 14272
rect 23711 14232 23756 14260
rect 23750 14220 23756 14232
rect 23808 14220 23814 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1486 14016 1492 14068
rect 1544 14056 1550 14068
rect 1673 14059 1731 14065
rect 1673 14056 1685 14059
rect 1544 14028 1685 14056
rect 1544 14016 1550 14028
rect 1673 14025 1685 14028
rect 1719 14025 1731 14059
rect 1673 14019 1731 14025
rect 2041 14059 2099 14065
rect 2041 14025 2053 14059
rect 2087 14056 2099 14059
rect 2774 14056 2780 14068
rect 2087 14028 2780 14056
rect 2087 14025 2099 14028
rect 2041 14019 2099 14025
rect 1688 13852 1716 14019
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 5629 14059 5687 14065
rect 5629 14056 5641 14059
rect 4212 14028 5641 14056
rect 4212 14016 4218 14028
rect 5629 14025 5641 14028
rect 5675 14025 5687 14059
rect 5629 14019 5687 14025
rect 6089 14059 6147 14065
rect 6089 14025 6101 14059
rect 6135 14056 6147 14059
rect 6178 14056 6184 14068
rect 6135 14028 6184 14056
rect 6135 14025 6147 14028
rect 6089 14019 6147 14025
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 6270 14016 6276 14068
rect 6328 14056 6334 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 6328 14028 6377 14056
rect 6328 14016 6334 14028
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 8110 14056 8116 14068
rect 8071 14028 8116 14056
rect 6365 14019 6423 14025
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 8294 14016 8300 14068
rect 8352 14056 8358 14068
rect 8803 14059 8861 14065
rect 8803 14056 8815 14059
rect 8352 14028 8815 14056
rect 8352 14016 8358 14028
rect 8803 14025 8815 14028
rect 8849 14025 8861 14059
rect 9766 14056 9772 14068
rect 9727 14028 9772 14056
rect 8803 14019 8861 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11241 14059 11299 14065
rect 11241 14056 11253 14059
rect 11112 14028 11253 14056
rect 11112 14016 11118 14028
rect 11241 14025 11253 14028
rect 11287 14025 11299 14059
rect 11698 14056 11704 14068
rect 11659 14028 11704 14056
rect 11241 14019 11299 14025
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 12894 14016 12900 14068
rect 12952 14056 12958 14068
rect 14001 14059 14059 14065
rect 14001 14056 14013 14059
rect 12952 14028 14013 14056
rect 12952 14016 12958 14028
rect 14001 14025 14013 14028
rect 14047 14025 14059 14059
rect 14001 14019 14059 14025
rect 18966 14016 18972 14068
rect 19024 14056 19030 14068
rect 19061 14059 19119 14065
rect 19061 14056 19073 14059
rect 19024 14028 19073 14056
rect 19024 14016 19030 14028
rect 19061 14025 19073 14028
rect 19107 14025 19119 14059
rect 19061 14019 19119 14025
rect 20993 14059 21051 14065
rect 20993 14025 21005 14059
rect 21039 14056 21051 14059
rect 21082 14056 21088 14068
rect 21039 14028 21088 14056
rect 21039 14025 21051 14028
rect 20993 14019 21051 14025
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 24670 14056 24676 14068
rect 24631 14028 24676 14056
rect 24670 14016 24676 14028
rect 24728 14016 24734 14068
rect 24854 14016 24860 14068
rect 24912 14056 24918 14068
rect 25363 14059 25421 14065
rect 25363 14056 25375 14059
rect 24912 14028 25375 14056
rect 24912 14016 24918 14028
rect 25363 14025 25375 14028
rect 25409 14025 25421 14059
rect 25363 14019 25421 14025
rect 2682 13948 2688 14000
rect 2740 13988 2746 14000
rect 3789 13991 3847 13997
rect 3789 13988 3801 13991
rect 2740 13960 3801 13988
rect 2740 13948 2746 13960
rect 3789 13957 3801 13960
rect 3835 13957 3847 13991
rect 7466 13988 7472 14000
rect 3789 13951 3847 13957
rect 7208 13960 7472 13988
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13920 2835 13923
rect 3142 13920 3148 13932
rect 2823 13892 3148 13920
rect 2823 13889 2835 13892
rect 2777 13883 2835 13889
rect 3142 13880 3148 13892
rect 3200 13880 3206 13932
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13920 4215 13923
rect 4203 13892 5212 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 5184 13864 5212 13892
rect 5534 13880 5540 13932
rect 5592 13920 5598 13932
rect 6270 13920 6276 13932
rect 5592 13892 6276 13920
rect 5592 13880 5598 13892
rect 6270 13880 6276 13892
rect 6328 13880 6334 13932
rect 7208 13929 7236 13960
rect 7466 13948 7472 13960
rect 7524 13988 7530 14000
rect 8662 13988 8668 14000
rect 7524 13960 8668 13988
rect 7524 13948 7530 13960
rect 8662 13948 8668 13960
rect 8720 13988 8726 14000
rect 8720 13960 10732 13988
rect 8720 13948 8726 13960
rect 7193 13923 7251 13929
rect 7193 13889 7205 13923
rect 7239 13889 7251 13923
rect 10045 13923 10103 13929
rect 10045 13920 10057 13923
rect 7193 13883 7251 13889
rect 9692 13892 10057 13920
rect 1857 13855 1915 13861
rect 1857 13852 1869 13855
rect 1688 13824 1869 13852
rect 1857 13821 1869 13824
rect 1903 13821 1915 13855
rect 1857 13815 1915 13821
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13852 2927 13855
rect 3326 13852 3332 13864
rect 2915 13824 3332 13852
rect 2915 13821 2927 13824
rect 2869 13815 2927 13821
rect 1872 13716 1900 13815
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 4525 13855 4583 13861
rect 4525 13821 4537 13855
rect 4571 13852 4583 13855
rect 4706 13852 4712 13864
rect 4571 13824 4712 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 4706 13812 4712 13824
rect 4764 13812 4770 13864
rect 5166 13852 5172 13864
rect 5127 13824 5172 13852
rect 5166 13812 5172 13824
rect 5224 13812 5230 13864
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 8202 13852 8208 13864
rect 7883 13824 8208 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 8732 13855 8790 13861
rect 8732 13852 8744 13855
rect 8444 13824 8744 13852
rect 8444 13812 8450 13824
rect 8732 13821 8744 13824
rect 8778 13852 8790 13855
rect 9214 13852 9220 13864
rect 8778 13824 9220 13852
rect 8778 13821 8790 13824
rect 8732 13815 8790 13821
rect 9214 13812 9220 13824
rect 9272 13812 9278 13864
rect 9692 13852 9720 13892
rect 10045 13889 10057 13892
rect 10091 13889 10103 13923
rect 10045 13883 10103 13889
rect 10704 13861 10732 13960
rect 12986 13948 12992 14000
rect 13044 13988 13050 14000
rect 13357 13991 13415 13997
rect 13357 13988 13369 13991
rect 13044 13960 13369 13988
rect 13044 13948 13050 13960
rect 13357 13957 13369 13960
rect 13403 13988 13415 13991
rect 13630 13988 13636 14000
rect 13403 13960 13636 13988
rect 13403 13957 13415 13960
rect 13357 13951 13415 13957
rect 13630 13948 13636 13960
rect 13688 13948 13694 14000
rect 13814 13948 13820 14000
rect 13872 13988 13878 14000
rect 14829 13991 14887 13997
rect 14829 13988 14841 13991
rect 13872 13960 14841 13988
rect 13872 13948 13878 13960
rect 14829 13957 14841 13960
rect 14875 13988 14887 13991
rect 14921 13991 14979 13997
rect 14921 13988 14933 13991
rect 14875 13960 14933 13988
rect 14875 13957 14887 13960
rect 14829 13951 14887 13957
rect 14921 13957 14933 13960
rect 14967 13988 14979 13991
rect 16117 13991 16175 13997
rect 16117 13988 16129 13991
rect 14967 13960 16129 13988
rect 14967 13957 14979 13960
rect 14921 13951 14979 13957
rect 16117 13957 16129 13960
rect 16163 13957 16175 13991
rect 16117 13951 16175 13957
rect 16853 13991 16911 13997
rect 16853 13957 16865 13991
rect 16899 13988 16911 13991
rect 17865 13991 17923 13997
rect 17865 13988 17877 13991
rect 16899 13960 17877 13988
rect 16899 13957 16911 13960
rect 16853 13951 16911 13957
rect 17865 13957 17877 13960
rect 17911 13988 17923 13991
rect 18046 13988 18052 14000
rect 17911 13960 18052 13988
rect 17911 13957 17923 13960
rect 17865 13951 17923 13957
rect 18046 13948 18052 13960
rect 18104 13948 18110 14000
rect 18782 13948 18788 14000
rect 18840 13988 18846 14000
rect 20441 13991 20499 13997
rect 20441 13988 20453 13991
rect 18840 13960 20453 13988
rect 18840 13948 18846 13960
rect 20441 13957 20453 13960
rect 20487 13988 20499 13991
rect 22278 13988 22284 14000
rect 20487 13960 22284 13988
rect 20487 13957 20499 13960
rect 20441 13951 20499 13957
rect 12434 13880 12440 13932
rect 12492 13920 12498 13932
rect 14645 13923 14703 13929
rect 12492 13892 12537 13920
rect 12492 13880 12498 13892
rect 14645 13889 14657 13923
rect 14691 13920 14703 13923
rect 15194 13920 15200 13932
rect 14691 13892 15200 13920
rect 14691 13889 14703 13892
rect 14645 13883 14703 13889
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 15841 13923 15899 13929
rect 15841 13889 15853 13923
rect 15887 13920 15899 13923
rect 15930 13920 15936 13932
rect 15887 13892 15936 13920
rect 15887 13889 15899 13892
rect 15841 13883 15899 13889
rect 15930 13880 15936 13892
rect 15988 13880 15994 13932
rect 17083 13923 17141 13929
rect 17083 13889 17095 13923
rect 17129 13920 17141 13923
rect 18141 13923 18199 13929
rect 18141 13920 18153 13923
rect 17129 13892 18153 13920
rect 17129 13889 17141 13892
rect 17083 13883 17141 13889
rect 18141 13889 18153 13892
rect 18187 13920 18199 13923
rect 18230 13920 18236 13932
rect 18187 13892 18236 13920
rect 18187 13889 18199 13892
rect 18141 13883 18199 13889
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 20070 13920 20076 13932
rect 19935 13892 20076 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 20070 13880 20076 13892
rect 20128 13920 20134 13932
rect 20622 13920 20628 13932
rect 20128 13892 20628 13920
rect 20128 13880 20134 13892
rect 20622 13880 20628 13892
rect 20680 13880 20686 13932
rect 21468 13929 21496 13960
rect 22278 13948 22284 13960
rect 22336 13988 22342 14000
rect 23014 13988 23020 14000
rect 22336 13960 23020 13988
rect 22336 13948 22342 13960
rect 23014 13948 23020 13960
rect 23072 13948 23078 14000
rect 21453 13923 21511 13929
rect 21453 13889 21465 13923
rect 21499 13889 21511 13923
rect 21726 13920 21732 13932
rect 21687 13892 21732 13920
rect 21453 13883 21511 13889
rect 21726 13880 21732 13892
rect 21784 13880 21790 13932
rect 9508 13824 9720 13852
rect 10689 13855 10747 13861
rect 2409 13787 2467 13793
rect 2409 13753 2421 13787
rect 2455 13784 2467 13787
rect 3231 13787 3289 13793
rect 3231 13784 3243 13787
rect 2455 13756 3243 13784
rect 2455 13753 2467 13756
rect 2409 13747 2467 13753
rect 3231 13753 3243 13756
rect 3277 13784 3289 13787
rect 3970 13784 3976 13796
rect 3277 13756 3976 13784
rect 3277 13753 3289 13756
rect 3231 13747 3289 13753
rect 3970 13744 3976 13756
rect 4028 13744 4034 13796
rect 5350 13784 5356 13796
rect 5311 13756 5356 13784
rect 5350 13744 5356 13756
rect 5408 13744 5414 13796
rect 7282 13744 7288 13796
rect 7340 13784 7346 13796
rect 7340 13756 7385 13784
rect 7340 13744 7346 13756
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 9508 13784 9536 13824
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 10962 13852 10968 13864
rect 10735 13824 10968 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 10962 13812 10968 13824
rect 11020 13812 11026 13864
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13852 14887 13855
rect 15948 13852 15976 13880
rect 14875 13824 15056 13852
rect 15948 13824 16528 13852
rect 14875 13821 14887 13824
rect 14829 13815 14887 13821
rect 9180 13756 9536 13784
rect 9180 13744 9186 13756
rect 10134 13744 10140 13796
rect 10192 13784 10198 13796
rect 12758 13787 12816 13793
rect 12758 13784 12770 13787
rect 10192 13756 10237 13784
rect 12176 13756 12770 13784
rect 10192 13744 10198 13756
rect 5534 13716 5540 13728
rect 1872 13688 5540 13716
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 9214 13716 9220 13728
rect 9175 13688 9220 13716
rect 9214 13676 9220 13688
rect 9272 13676 9278 13728
rect 9306 13676 9312 13728
rect 9364 13716 9370 13728
rect 11330 13716 11336 13728
rect 9364 13688 11336 13716
rect 9364 13676 9370 13688
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 12066 13676 12072 13728
rect 12124 13716 12130 13728
rect 12176 13725 12204 13756
rect 12758 13753 12770 13756
rect 12804 13753 12816 13787
rect 15028 13784 15056 13824
rect 15289 13787 15347 13793
rect 15289 13784 15301 13787
rect 15028 13756 15301 13784
rect 12758 13747 12816 13753
rect 15289 13753 15301 13756
rect 15335 13753 15347 13787
rect 16500 13784 16528 13824
rect 16850 13812 16856 13864
rect 16908 13852 16914 13864
rect 16980 13855 17038 13861
rect 16980 13852 16992 13855
rect 16908 13824 16992 13852
rect 16908 13812 16914 13824
rect 16980 13821 16992 13824
rect 17026 13852 17038 13855
rect 17218 13852 17224 13864
rect 17026 13824 17224 13852
rect 17026 13821 17038 13824
rect 16980 13815 17038 13821
rect 17218 13812 17224 13824
rect 17276 13852 17282 13864
rect 17405 13855 17463 13861
rect 17405 13852 17417 13855
rect 17276 13824 17417 13852
rect 17276 13812 17282 13824
rect 17405 13821 17417 13824
rect 17451 13821 17463 13855
rect 17405 13815 17463 13821
rect 22557 13855 22615 13861
rect 22557 13821 22569 13855
rect 22603 13852 22615 13855
rect 22738 13852 22744 13864
rect 22603 13824 22744 13852
rect 22603 13821 22615 13824
rect 22557 13815 22615 13821
rect 22738 13812 22744 13824
rect 22796 13812 22802 13864
rect 23750 13852 23756 13864
rect 23711 13824 23756 13852
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 24121 13855 24179 13861
rect 24121 13821 24133 13855
rect 24167 13821 24179 13855
rect 24121 13815 24179 13821
rect 17310 13784 17316 13796
rect 16500 13756 17316 13784
rect 15289 13747 15347 13753
rect 17310 13744 17316 13756
rect 17368 13744 17374 13796
rect 18138 13744 18144 13796
rect 18196 13784 18202 13796
rect 18233 13787 18291 13793
rect 18233 13784 18245 13787
rect 18196 13756 18245 13784
rect 18196 13744 18202 13756
rect 18233 13753 18245 13756
rect 18279 13753 18291 13787
rect 18233 13747 18291 13753
rect 18785 13787 18843 13793
rect 18785 13753 18797 13787
rect 18831 13784 18843 13787
rect 18874 13784 18880 13796
rect 18831 13756 18880 13784
rect 18831 13753 18843 13756
rect 18785 13747 18843 13753
rect 18874 13744 18880 13756
rect 18932 13744 18938 13796
rect 19705 13787 19763 13793
rect 19705 13753 19717 13787
rect 19751 13784 19763 13787
rect 19981 13787 20039 13793
rect 19981 13784 19993 13787
rect 19751 13756 19993 13784
rect 19751 13753 19763 13756
rect 19705 13747 19763 13753
rect 19981 13753 19993 13756
rect 20027 13784 20039 13787
rect 20162 13784 20168 13796
rect 20027 13756 20168 13784
rect 20027 13753 20039 13756
rect 19981 13747 20039 13753
rect 20162 13744 20168 13756
rect 20220 13744 20226 13796
rect 21545 13787 21603 13793
rect 21545 13753 21557 13787
rect 21591 13784 21603 13787
rect 21634 13784 21640 13796
rect 21591 13756 21640 13784
rect 21591 13753 21603 13756
rect 21545 13747 21603 13753
rect 21634 13744 21640 13756
rect 21692 13784 21698 13796
rect 22186 13784 22192 13796
rect 21692 13756 22192 13784
rect 21692 13744 21698 13756
rect 22186 13744 22192 13756
rect 22244 13744 22250 13796
rect 22922 13784 22928 13796
rect 22835 13756 22928 13784
rect 22922 13744 22928 13756
rect 22980 13784 22986 13796
rect 23385 13787 23443 13793
rect 23385 13784 23397 13787
rect 22980 13756 23397 13784
rect 22980 13744 22986 13756
rect 23385 13753 23397 13756
rect 23431 13784 23443 13787
rect 23842 13784 23848 13796
rect 23431 13756 23848 13784
rect 23431 13753 23443 13756
rect 23385 13747 23443 13753
rect 23842 13744 23848 13756
rect 23900 13784 23906 13796
rect 24136 13784 24164 13815
rect 24946 13812 24952 13864
rect 25004 13852 25010 13864
rect 25292 13855 25350 13861
rect 25292 13852 25304 13855
rect 25004 13824 25304 13852
rect 25004 13812 25010 13824
rect 25292 13821 25304 13824
rect 25338 13852 25350 13855
rect 25685 13855 25743 13861
rect 25685 13852 25697 13855
rect 25338 13824 25697 13852
rect 25338 13821 25350 13824
rect 25292 13815 25350 13821
rect 25685 13821 25697 13824
rect 25731 13821 25743 13855
rect 25685 13815 25743 13821
rect 23900 13756 24164 13784
rect 23900 13744 23906 13756
rect 12161 13719 12219 13725
rect 12161 13716 12173 13719
rect 12124 13688 12173 13716
rect 12124 13676 12130 13688
rect 12161 13685 12173 13688
rect 12207 13685 12219 13719
rect 12161 13679 12219 13685
rect 23474 13676 23480 13728
rect 23532 13716 23538 13728
rect 23753 13719 23811 13725
rect 23753 13716 23765 13719
rect 23532 13688 23765 13716
rect 23532 13676 23538 13688
rect 23753 13685 23765 13688
rect 23799 13685 23811 13719
rect 23753 13679 23811 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 3326 13512 3332 13524
rect 3287 13484 3332 13512
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 3881 13515 3939 13521
rect 3881 13481 3893 13515
rect 3927 13512 3939 13515
rect 4062 13512 4068 13524
rect 3927 13484 4068 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 2409 13447 2467 13453
rect 2409 13413 2421 13447
rect 2455 13444 2467 13447
rect 2682 13444 2688 13456
rect 2455 13416 2688 13444
rect 2455 13413 2467 13416
rect 2409 13407 2467 13413
rect 2682 13404 2688 13416
rect 2740 13404 2746 13456
rect 2774 13404 2780 13456
rect 2832 13444 2838 13456
rect 3896 13444 3924 13475
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 6181 13515 6239 13521
rect 6181 13481 6193 13515
rect 6227 13512 6239 13515
rect 6362 13512 6368 13524
rect 6227 13484 6368 13512
rect 6227 13481 6239 13484
rect 6181 13475 6239 13481
rect 2832 13416 3924 13444
rect 2832 13404 2838 13416
rect 3970 13404 3976 13456
rect 4028 13444 4034 13456
rect 4427 13447 4485 13453
rect 4427 13444 4439 13447
rect 4028 13416 4439 13444
rect 4028 13404 4034 13416
rect 4427 13413 4439 13416
rect 4473 13444 4485 13447
rect 4890 13444 4896 13456
rect 4473 13416 4896 13444
rect 4473 13413 4485 13416
rect 4427 13407 4485 13413
rect 4890 13404 4896 13416
rect 4948 13404 4954 13456
rect 6288 13385 6316 13484
rect 6362 13472 6368 13484
rect 6420 13472 6426 13524
rect 7193 13515 7251 13521
rect 7193 13481 7205 13515
rect 7239 13512 7251 13515
rect 7282 13512 7288 13524
rect 7239 13484 7288 13512
rect 7239 13481 7251 13484
rect 7193 13475 7251 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7466 13512 7472 13524
rect 7427 13484 7472 13512
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 9122 13512 9128 13524
rect 9083 13484 9128 13512
rect 9122 13472 9128 13484
rect 9180 13472 9186 13524
rect 9493 13515 9551 13521
rect 9493 13481 9505 13515
rect 9539 13512 9551 13515
rect 9582 13512 9588 13524
rect 9539 13484 9588 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 10597 13515 10655 13521
rect 10597 13512 10609 13515
rect 10192 13484 10609 13512
rect 10192 13472 10198 13484
rect 10597 13481 10609 13484
rect 10643 13481 10655 13515
rect 10597 13475 10655 13481
rect 11054 13472 11060 13524
rect 11112 13512 11118 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 11112 13484 11621 13512
rect 11112 13472 11118 13484
rect 11609 13481 11621 13484
rect 11655 13481 11667 13515
rect 11609 13475 11667 13481
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 13541 13515 13599 13521
rect 12492 13484 12537 13512
rect 12492 13472 12498 13484
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 13722 13512 13728 13524
rect 13587 13484 13728 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 14826 13472 14832 13524
rect 14884 13512 14890 13524
rect 15013 13515 15071 13521
rect 15013 13512 15025 13515
rect 14884 13484 15025 13512
rect 14884 13472 14890 13484
rect 15013 13481 15025 13484
rect 15059 13481 15071 13515
rect 15013 13475 15071 13481
rect 17862 13472 17868 13524
rect 17920 13512 17926 13524
rect 17957 13515 18015 13521
rect 17957 13512 17969 13515
rect 17920 13484 17969 13512
rect 17920 13472 17926 13484
rect 17957 13481 17969 13484
rect 18003 13481 18015 13515
rect 18230 13512 18236 13524
rect 18191 13484 18236 13512
rect 17957 13475 18015 13481
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 19889 13515 19947 13521
rect 19889 13481 19901 13515
rect 19935 13512 19947 13515
rect 20070 13512 20076 13524
rect 19935 13484 20076 13512
rect 19935 13481 19947 13484
rect 19889 13475 19947 13481
rect 20070 13472 20076 13484
rect 20128 13472 20134 13524
rect 20717 13515 20775 13521
rect 20717 13481 20729 13515
rect 20763 13512 20775 13515
rect 20990 13512 20996 13524
rect 20763 13484 20996 13512
rect 20763 13481 20775 13484
rect 20717 13475 20775 13481
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 6546 13404 6552 13456
rect 6604 13453 6610 13456
rect 6604 13447 6652 13453
rect 6604 13413 6606 13447
rect 6640 13413 6652 13447
rect 8202 13444 8208 13456
rect 8163 13416 8208 13444
rect 6604 13407 6652 13413
rect 6604 13404 6610 13407
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 9858 13404 9864 13456
rect 9916 13444 9922 13456
rect 9998 13447 10056 13453
rect 9998 13444 10010 13447
rect 9916 13416 10010 13444
rect 9916 13404 9922 13416
rect 9998 13413 10010 13416
rect 10044 13444 10056 13447
rect 12066 13444 12072 13456
rect 10044 13416 12072 13444
rect 10044 13413 10056 13416
rect 9998 13407 10056 13413
rect 12066 13404 12072 13416
rect 12124 13444 12130 13456
rect 12986 13453 12992 13456
rect 12942 13447 12992 13453
rect 12942 13444 12954 13447
rect 12124 13416 12954 13444
rect 12124 13404 12130 13416
rect 12942 13413 12954 13416
rect 12988 13413 12992 13447
rect 12942 13407 12992 13413
rect 12986 13404 12992 13407
rect 13044 13444 13050 13456
rect 13044 13416 13090 13444
rect 13044 13404 13050 13416
rect 15378 13404 15384 13456
rect 15436 13444 15442 13456
rect 15473 13447 15531 13453
rect 15473 13444 15485 13447
rect 15436 13416 15485 13444
rect 15436 13404 15442 13416
rect 15473 13413 15485 13416
rect 15519 13413 15531 13447
rect 16022 13444 16028 13456
rect 15983 13416 16028 13444
rect 15473 13407 15531 13413
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 17034 13444 17040 13456
rect 16995 13416 17040 13444
rect 17034 13404 17040 13416
rect 17092 13404 17098 13456
rect 18598 13444 18604 13456
rect 18559 13416 18604 13444
rect 18598 13404 18604 13416
rect 18656 13404 18662 13456
rect 19242 13404 19248 13456
rect 19300 13444 19306 13456
rect 19521 13447 19579 13453
rect 19521 13444 19533 13447
rect 19300 13416 19533 13444
rect 19300 13404 19306 13416
rect 19521 13413 19533 13416
rect 19567 13444 19579 13447
rect 20162 13444 20168 13456
rect 19567 13416 20168 13444
rect 19567 13413 19579 13416
rect 19521 13407 19579 13413
rect 20162 13404 20168 13416
rect 20220 13404 20226 13456
rect 21542 13444 21548 13456
rect 21503 13416 21548 13444
rect 21542 13404 21548 13416
rect 21600 13404 21606 13456
rect 23109 13447 23167 13453
rect 23109 13413 23121 13447
rect 23155 13444 23167 13447
rect 23382 13444 23388 13456
rect 23155 13416 23388 13444
rect 23155 13413 23167 13416
rect 23109 13407 23167 13413
rect 23382 13404 23388 13416
rect 23440 13404 23446 13456
rect 6273 13379 6331 13385
rect 6273 13345 6285 13379
rect 6319 13345 6331 13379
rect 11422 13376 11428 13388
rect 11383 13348 11428 13376
rect 6273 13339 6331 13345
rect 11422 13336 11428 13348
rect 11480 13336 11486 13388
rect 12618 13376 12624 13388
rect 12579 13348 12624 13376
rect 12618 13336 12624 13348
rect 12676 13336 12682 13388
rect 24210 13336 24216 13388
rect 24268 13376 24274 13388
rect 24524 13379 24582 13385
rect 24524 13376 24536 13379
rect 24268 13348 24536 13376
rect 24268 13336 24274 13348
rect 24524 13345 24536 13348
rect 24570 13345 24582 13379
rect 24524 13339 24582 13345
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13308 2375 13311
rect 2498 13308 2504 13320
rect 2363 13280 2504 13308
rect 2363 13277 2375 13280
rect 2317 13271 2375 13277
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 4062 13308 4068 13320
rect 4023 13280 4068 13308
rect 4062 13268 4068 13280
rect 4120 13268 4126 13320
rect 8110 13308 8116 13320
rect 8071 13280 8116 13308
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 8294 13268 8300 13320
rect 8352 13308 8358 13320
rect 8389 13311 8447 13317
rect 8389 13308 8401 13311
rect 8352 13280 8401 13308
rect 8352 13268 8358 13280
rect 8389 13277 8401 13280
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13308 9735 13311
rect 9766 13308 9772 13320
rect 9723 13280 9772 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 9766 13268 9772 13280
rect 9824 13308 9830 13320
rect 10778 13308 10784 13320
rect 9824 13280 10784 13308
rect 9824 13268 9830 13280
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 14550 13268 14556 13320
rect 14608 13308 14614 13320
rect 15381 13311 15439 13317
rect 15381 13308 15393 13311
rect 14608 13280 15393 13308
rect 14608 13268 14614 13280
rect 15381 13277 15393 13280
rect 15427 13277 15439 13311
rect 15381 13271 15439 13277
rect 16945 13311 17003 13317
rect 16945 13277 16957 13311
rect 16991 13308 17003 13311
rect 17218 13308 17224 13320
rect 16991 13280 17224 13308
rect 16991 13277 17003 13280
rect 16945 13271 17003 13277
rect 17218 13268 17224 13280
rect 17276 13268 17282 13320
rect 17310 13268 17316 13320
rect 17368 13308 17374 13320
rect 18506 13308 18512 13320
rect 17368 13280 17413 13308
rect 18467 13280 18512 13308
rect 17368 13268 17374 13280
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 18782 13308 18788 13320
rect 18743 13280 18788 13308
rect 18782 13268 18788 13280
rect 18840 13268 18846 13320
rect 21450 13308 21456 13320
rect 21411 13280 21456 13308
rect 21450 13268 21456 13280
rect 21508 13308 21514 13320
rect 21508 13280 22140 13308
rect 21508 13268 21514 13280
rect 22112 13252 22140 13280
rect 22462 13268 22468 13320
rect 22520 13308 22526 13320
rect 23017 13311 23075 13317
rect 23017 13308 23029 13311
rect 22520 13280 23029 13308
rect 22520 13268 22526 13280
rect 23017 13277 23029 13280
rect 23063 13308 23075 13311
rect 24627 13311 24685 13317
rect 24627 13308 24639 13311
rect 23063 13280 24639 13308
rect 23063 13277 23075 13280
rect 23017 13271 23075 13277
rect 24627 13277 24639 13280
rect 24673 13277 24685 13311
rect 24627 13271 24685 13277
rect 2866 13240 2872 13252
rect 2779 13212 2872 13240
rect 2866 13200 2872 13212
rect 2924 13240 2930 13252
rect 4614 13240 4620 13252
rect 2924 13212 4620 13240
rect 2924 13200 2930 13212
rect 4614 13200 4620 13212
rect 4672 13200 4678 13252
rect 9398 13200 9404 13252
rect 9456 13240 9462 13252
rect 11054 13240 11060 13252
rect 9456 13212 11060 13240
rect 9456 13200 9462 13212
rect 11054 13200 11060 13212
rect 11112 13200 11118 13252
rect 20714 13200 20720 13252
rect 20772 13240 20778 13252
rect 21726 13240 21732 13252
rect 20772 13212 21732 13240
rect 20772 13200 20778 13212
rect 21726 13200 21732 13212
rect 21784 13240 21790 13252
rect 22005 13243 22063 13249
rect 22005 13240 22017 13243
rect 21784 13212 22017 13240
rect 21784 13200 21790 13212
rect 22005 13209 22017 13212
rect 22051 13209 22063 13243
rect 22005 13203 22063 13209
rect 22094 13200 22100 13252
rect 22152 13240 22158 13252
rect 23569 13243 23627 13249
rect 23569 13240 23581 13243
rect 22152 13212 23581 13240
rect 22152 13200 22158 13212
rect 23569 13209 23581 13212
rect 23615 13209 23627 13243
rect 23569 13203 23627 13209
rect 1670 13172 1676 13184
rect 1631 13144 1676 13172
rect 1670 13132 1676 13144
rect 1728 13132 1734 13184
rect 3970 13132 3976 13184
rect 4028 13172 4034 13184
rect 4985 13175 5043 13181
rect 4985 13172 4997 13175
rect 4028 13144 4997 13172
rect 4028 13132 4034 13144
rect 4985 13141 4997 13144
rect 5031 13141 5043 13175
rect 7926 13172 7932 13184
rect 7887 13144 7932 13172
rect 4985 13135 5043 13141
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 9674 13132 9680 13184
rect 9732 13172 9738 13184
rect 11790 13172 11796 13184
rect 9732 13144 11796 13172
rect 9732 13132 9738 13144
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 13814 13172 13820 13184
rect 13775 13144 13820 13172
rect 13814 13132 13820 13144
rect 13872 13132 13878 13184
rect 21082 13172 21088 13184
rect 21043 13144 21088 13172
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1673 12971 1731 12977
rect 1673 12937 1685 12971
rect 1719 12968 1731 12971
rect 2498 12968 2504 12980
rect 1719 12940 2504 12968
rect 1719 12937 1731 12940
rect 1673 12931 1731 12937
rect 2498 12928 2504 12940
rect 2556 12928 2562 12980
rect 2682 12968 2688 12980
rect 2643 12940 2688 12968
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 4062 12928 4068 12980
rect 4120 12968 4126 12980
rect 5169 12971 5227 12977
rect 5169 12968 5181 12971
rect 4120 12940 5181 12968
rect 4120 12928 4126 12940
rect 5169 12937 5181 12940
rect 5215 12937 5227 12971
rect 5169 12931 5227 12937
rect 8110 12928 8116 12980
rect 8168 12968 8174 12980
rect 8389 12971 8447 12977
rect 8389 12968 8401 12971
rect 8168 12940 8401 12968
rect 8168 12928 8174 12940
rect 8389 12937 8401 12940
rect 8435 12968 8447 12971
rect 8478 12968 8484 12980
rect 8435 12940 8484 12968
rect 8435 12937 8447 12940
rect 8389 12931 8447 12937
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 8754 12968 8760 12980
rect 8715 12940 8760 12968
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 10778 12968 10784 12980
rect 10739 12940 10784 12968
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 11974 12968 11980 12980
rect 11480 12940 11980 12968
rect 11480 12928 11486 12940
rect 11974 12928 11980 12940
rect 12032 12968 12038 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 12032 12940 12173 12968
rect 12032 12928 12038 12940
rect 12161 12937 12173 12940
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 12667 12971 12725 12977
rect 12667 12937 12679 12971
rect 12713 12968 12725 12971
rect 13538 12968 13544 12980
rect 12713 12940 13544 12968
rect 12713 12937 12725 12940
rect 12667 12931 12725 12937
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 15378 12968 15384 12980
rect 15339 12940 15384 12968
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 21542 12928 21548 12980
rect 21600 12968 21606 12980
rect 22005 12971 22063 12977
rect 22005 12968 22017 12971
rect 21600 12940 22017 12968
rect 21600 12928 21606 12940
rect 22005 12937 22017 12940
rect 22051 12937 22063 12971
rect 22462 12968 22468 12980
rect 22423 12940 22468 12968
rect 22005 12931 22063 12937
rect 22462 12928 22468 12940
rect 22520 12928 22526 12980
rect 23382 12968 23388 12980
rect 23343 12940 23388 12968
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 24305 12971 24363 12977
rect 24305 12937 24317 12971
rect 24351 12968 24363 12971
rect 24762 12968 24768 12980
rect 24351 12940 24768 12968
rect 24351 12937 24363 12940
rect 24305 12931 24363 12937
rect 24762 12928 24768 12940
rect 24820 12968 24826 12980
rect 24857 12971 24915 12977
rect 24857 12968 24869 12971
rect 24820 12940 24869 12968
rect 24820 12928 24826 12940
rect 24857 12937 24869 12940
rect 24903 12937 24915 12971
rect 25590 12968 25596 12980
rect 25551 12940 25596 12968
rect 24857 12931 24915 12937
rect 25590 12928 25596 12940
rect 25648 12928 25654 12980
rect 1762 12860 1768 12912
rect 1820 12900 1826 12912
rect 1949 12903 2007 12909
rect 1949 12900 1961 12903
rect 1820 12872 1961 12900
rect 1820 12860 1826 12872
rect 1949 12869 1961 12872
rect 1995 12869 2007 12903
rect 1949 12863 2007 12869
rect 5905 12903 5963 12909
rect 5905 12869 5917 12903
rect 5951 12900 5963 12903
rect 6638 12900 6644 12912
rect 5951 12872 6644 12900
rect 5951 12869 5963 12872
rect 5905 12863 5963 12869
rect 6638 12860 6644 12872
rect 6696 12860 6702 12912
rect 7745 12903 7803 12909
rect 7745 12869 7757 12903
rect 7791 12869 7803 12903
rect 11149 12903 11207 12909
rect 11149 12900 11161 12903
rect 7745 12863 7803 12869
rect 10336 12872 11161 12900
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 2792 12804 3341 12832
rect 2792 12773 2820 12804
rect 3329 12801 3341 12804
rect 3375 12832 3387 12835
rect 4062 12832 4068 12844
rect 3375 12804 4068 12832
rect 3375 12801 3387 12804
rect 3329 12795 3387 12801
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12832 4583 12835
rect 4614 12832 4620 12844
rect 4571 12804 4620 12832
rect 4571 12801 4583 12804
rect 4525 12795 4583 12801
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 7760 12832 7788 12863
rect 10336 12844 10364 12872
rect 11149 12869 11161 12872
rect 11195 12869 11207 12903
rect 11149 12863 11207 12869
rect 12986 12860 12992 12912
rect 13044 12900 13050 12912
rect 13357 12903 13415 12909
rect 13357 12900 13369 12903
rect 13044 12872 13369 12900
rect 13044 12860 13050 12872
rect 13357 12869 13369 12872
rect 13403 12869 13415 12903
rect 15930 12900 15936 12912
rect 13357 12863 13415 12869
rect 14936 12872 15936 12900
rect 8113 12835 8171 12841
rect 8113 12832 8125 12835
rect 7760 12804 8125 12832
rect 8113 12801 8125 12804
rect 8159 12832 8171 12835
rect 8202 12832 8208 12844
rect 8159 12804 8208 12832
rect 8159 12801 8171 12804
rect 8113 12795 8171 12801
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 9861 12835 9919 12841
rect 9861 12801 9873 12835
rect 9907 12832 9919 12835
rect 10318 12832 10324 12844
rect 9907 12804 10324 12832
rect 9907 12801 9919 12804
rect 9861 12795 9919 12801
rect 10318 12792 10324 12804
rect 10376 12792 10382 12844
rect 11054 12792 11060 12844
rect 11112 12832 11118 12844
rect 11471 12835 11529 12841
rect 11471 12832 11483 12835
rect 11112 12804 11483 12832
rect 11112 12792 11118 12804
rect 11471 12801 11483 12804
rect 11517 12801 11529 12835
rect 11471 12795 11529 12801
rect 12434 12792 12440 12844
rect 12492 12832 12498 12844
rect 13633 12835 13691 12841
rect 13633 12832 13645 12835
rect 12492 12804 13645 12832
rect 12492 12792 12498 12804
rect 13633 12801 13645 12804
rect 13679 12832 13691 12835
rect 13814 12832 13820 12844
rect 13679 12804 13820 12832
rect 13679 12801 13691 12804
rect 13633 12795 13691 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14090 12832 14096 12844
rect 14051 12804 14096 12832
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 1765 12767 1823 12773
rect 1765 12733 1777 12767
rect 1811 12764 1823 12767
rect 2317 12767 2375 12773
rect 2317 12764 2329 12767
rect 1811 12736 2329 12764
rect 1811 12733 1823 12736
rect 1765 12727 1823 12733
rect 2317 12733 2329 12736
rect 2363 12764 2375 12767
rect 2777 12767 2835 12773
rect 2777 12764 2789 12767
rect 2363 12736 2789 12764
rect 2363 12733 2375 12736
rect 2317 12727 2375 12733
rect 2777 12733 2789 12736
rect 2823 12733 2835 12767
rect 2777 12727 2835 12733
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12764 5779 12767
rect 6822 12764 6828 12776
rect 5767 12736 5801 12764
rect 6783 12736 6828 12764
rect 5767 12733 5779 12736
rect 5721 12727 5779 12733
rect 3697 12699 3755 12705
rect 3697 12665 3709 12699
rect 3743 12696 3755 12699
rect 3878 12696 3884 12708
rect 3743 12668 3884 12696
rect 3743 12665 3755 12668
rect 3697 12659 3755 12665
rect 3878 12656 3884 12668
rect 3936 12656 3942 12708
rect 3970 12656 3976 12708
rect 4028 12696 4034 12708
rect 5629 12699 5687 12705
rect 4028 12668 4073 12696
rect 4028 12656 4034 12668
rect 5629 12665 5641 12699
rect 5675 12696 5687 12699
rect 5736 12696 5764 12727
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 7282 12724 7288 12776
rect 7340 12764 7346 12776
rect 8573 12767 8631 12773
rect 8573 12764 8585 12767
rect 7340 12736 8585 12764
rect 7340 12724 7346 12736
rect 8573 12733 8585 12736
rect 8619 12764 8631 12767
rect 9033 12767 9091 12773
rect 9033 12764 9045 12767
rect 8619 12736 9045 12764
rect 8619 12733 8631 12736
rect 8573 12727 8631 12733
rect 9033 12733 9045 12736
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 11238 12724 11244 12776
rect 11296 12764 11302 12776
rect 11368 12767 11426 12773
rect 11368 12764 11380 12767
rect 11296 12736 11380 12764
rect 11296 12724 11302 12736
rect 11368 12733 11380 12736
rect 11414 12764 11426 12767
rect 11793 12767 11851 12773
rect 11793 12764 11805 12767
rect 11414 12736 11805 12764
rect 11414 12733 11426 12736
rect 11368 12727 11426 12733
rect 11793 12733 11805 12736
rect 11839 12764 11851 12767
rect 12066 12764 12072 12776
rect 11839 12736 12072 12764
rect 11839 12733 11851 12736
rect 11793 12727 11851 12733
rect 12066 12724 12072 12736
rect 12124 12724 12130 12776
rect 12596 12767 12654 12773
rect 12596 12733 12608 12767
rect 12642 12764 12654 12767
rect 12710 12764 12716 12776
rect 12642 12736 12716 12764
rect 12642 12733 12654 12736
rect 12596 12727 12654 12733
rect 12710 12724 12716 12736
rect 12768 12764 12774 12776
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12768 12736 13001 12764
rect 12768 12724 12774 12736
rect 12989 12733 13001 12736
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 5994 12696 6000 12708
rect 5675 12668 6000 12696
rect 5675 12665 5687 12668
rect 5629 12659 5687 12665
rect 5994 12656 6000 12668
rect 6052 12656 6058 12708
rect 6365 12699 6423 12705
rect 6365 12665 6377 12699
rect 6411 12696 6423 12699
rect 6546 12696 6552 12708
rect 6411 12668 6552 12696
rect 6411 12665 6423 12668
rect 6365 12659 6423 12665
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 2961 12631 3019 12637
rect 2961 12628 2973 12631
rect 2832 12600 2973 12628
rect 2832 12588 2838 12600
rect 2961 12597 2973 12600
rect 3007 12597 3019 12631
rect 4890 12628 4896 12640
rect 4803 12600 4896 12628
rect 2961 12591 3019 12597
rect 4890 12588 4896 12600
rect 4948 12628 4954 12640
rect 6380 12628 6408 12659
rect 6546 12656 6552 12668
rect 6604 12696 6610 12708
rect 7098 12696 7104 12708
rect 6604 12668 7104 12696
rect 6604 12656 6610 12668
rect 7098 12656 7104 12668
rect 7156 12705 7162 12708
rect 7156 12699 7204 12705
rect 7156 12665 7158 12699
rect 7192 12665 7204 12699
rect 7156 12659 7204 12665
rect 9677 12699 9735 12705
rect 9677 12665 9689 12699
rect 9723 12696 9735 12699
rect 9858 12696 9864 12708
rect 9723 12668 9864 12696
rect 9723 12665 9735 12668
rect 9677 12659 9735 12665
rect 7156 12656 7162 12659
rect 9858 12656 9864 12668
rect 9916 12656 9922 12708
rect 9953 12699 10011 12705
rect 9953 12665 9965 12699
rect 9999 12696 10011 12699
rect 10134 12696 10140 12708
rect 9999 12668 10140 12696
rect 9999 12665 10011 12668
rect 9953 12659 10011 12665
rect 10134 12656 10140 12668
rect 10192 12656 10198 12708
rect 10505 12699 10563 12705
rect 10505 12665 10517 12699
rect 10551 12696 10563 12699
rect 11054 12696 11060 12708
rect 10551 12668 11060 12696
rect 10551 12665 10563 12668
rect 10505 12659 10563 12665
rect 11054 12656 11060 12668
rect 11112 12656 11118 12708
rect 13722 12696 13728 12708
rect 13683 12668 13728 12696
rect 13722 12656 13728 12668
rect 13780 12696 13786 12708
rect 14936 12705 14964 12872
rect 15930 12860 15936 12872
rect 15988 12860 15994 12912
rect 18874 12900 18880 12912
rect 18835 12872 18880 12900
rect 18874 12860 18880 12872
rect 18932 12860 18938 12912
rect 22278 12860 22284 12912
rect 22336 12900 22342 12912
rect 23400 12900 23428 12928
rect 22336 12872 23428 12900
rect 22336 12860 22342 12872
rect 24210 12860 24216 12912
rect 24268 12900 24274 12912
rect 24489 12903 24547 12909
rect 24489 12900 24501 12903
rect 24268 12872 24501 12900
rect 24268 12860 24274 12872
rect 24489 12869 24501 12872
rect 24535 12869 24547 12903
rect 24489 12863 24547 12869
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 16022 12832 16028 12844
rect 15620 12804 16028 12832
rect 15620 12792 15626 12804
rect 16022 12792 16028 12804
rect 16080 12832 16086 12844
rect 16117 12835 16175 12841
rect 16117 12832 16129 12835
rect 16080 12804 16129 12832
rect 16080 12792 16086 12804
rect 16117 12801 16129 12804
rect 16163 12801 16175 12835
rect 16117 12795 16175 12801
rect 17954 12792 17960 12844
rect 18012 12832 18018 12844
rect 18138 12832 18144 12844
rect 18012 12804 18144 12832
rect 18012 12792 18018 12804
rect 18138 12792 18144 12804
rect 18196 12832 18202 12844
rect 18325 12835 18383 12841
rect 18325 12832 18337 12835
rect 18196 12804 18337 12832
rect 18196 12792 18202 12804
rect 18325 12801 18337 12804
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 20622 12792 20628 12844
rect 20680 12832 20686 12844
rect 20809 12835 20867 12841
rect 20809 12832 20821 12835
rect 20680 12804 20821 12832
rect 20680 12792 20686 12804
rect 20809 12801 20821 12804
rect 20855 12832 20867 12835
rect 21082 12832 21088 12844
rect 20855 12804 21088 12832
rect 20855 12801 20867 12804
rect 20809 12795 20867 12801
rect 21082 12792 21088 12804
rect 21140 12792 21146 12844
rect 21450 12792 21456 12844
rect 21508 12832 21514 12844
rect 22002 12832 22008 12844
rect 21508 12804 22008 12832
rect 21508 12792 21514 12804
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 22462 12792 22468 12844
rect 22520 12832 22526 12844
rect 22738 12832 22744 12844
rect 22520 12804 22744 12832
rect 22520 12792 22526 12804
rect 22738 12792 22744 12804
rect 22796 12792 22802 12844
rect 23109 12835 23167 12841
rect 23109 12801 23121 12835
rect 23155 12832 23167 12835
rect 23155 12804 24808 12832
rect 23155 12801 23167 12804
rect 23109 12795 23167 12801
rect 19794 12724 19800 12776
rect 19852 12773 19858 12776
rect 19852 12767 19890 12773
rect 19878 12764 19890 12767
rect 20257 12767 20315 12773
rect 20257 12764 20269 12767
rect 19878 12736 20269 12764
rect 19878 12733 19890 12736
rect 19852 12727 19890 12733
rect 20257 12733 20269 12736
rect 20303 12733 20315 12767
rect 20257 12727 20315 12733
rect 22624 12767 22682 12773
rect 22624 12733 22636 12767
rect 22670 12764 22682 12767
rect 23124 12764 23152 12795
rect 22670 12736 23152 12764
rect 24096 12767 24154 12773
rect 22670 12733 22682 12736
rect 22624 12727 22682 12733
rect 24096 12733 24108 12767
rect 24142 12764 24154 12767
rect 24305 12767 24363 12773
rect 24305 12764 24317 12767
rect 24142 12736 24317 12764
rect 24142 12733 24154 12736
rect 24096 12727 24154 12733
rect 24305 12733 24317 12736
rect 24351 12733 24363 12767
rect 24780 12764 24808 12804
rect 24854 12792 24860 12844
rect 24912 12832 24918 12844
rect 25222 12832 25228 12844
rect 24912 12804 25228 12832
rect 24912 12792 24918 12804
rect 25222 12792 25228 12804
rect 25280 12792 25286 12844
rect 25092 12767 25150 12773
rect 25092 12764 25104 12767
rect 24780 12736 25104 12764
rect 24305 12727 24363 12733
rect 25092 12733 25104 12736
rect 25138 12764 25150 12767
rect 25590 12764 25596 12776
rect 25138 12736 25596 12764
rect 25138 12733 25150 12736
rect 25092 12727 25150 12733
rect 19852 12724 19858 12727
rect 25590 12724 25596 12736
rect 25648 12724 25654 12776
rect 14921 12699 14979 12705
rect 14921 12696 14933 12699
rect 13780 12668 14933 12696
rect 13780 12656 13786 12668
rect 14921 12665 14933 12668
rect 14967 12665 14979 12699
rect 15841 12699 15899 12705
rect 15841 12696 15853 12699
rect 14921 12659 14979 12665
rect 15764 12668 15853 12696
rect 4948 12600 6408 12628
rect 4948 12588 4954 12600
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 10042 12628 10048 12640
rect 9824 12600 10048 12628
rect 9824 12588 9830 12600
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 14550 12628 14556 12640
rect 14511 12600 14556 12628
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 15764 12628 15792 12668
rect 15841 12665 15853 12668
rect 15887 12665 15899 12699
rect 15841 12659 15899 12665
rect 15930 12656 15936 12708
rect 15988 12696 15994 12708
rect 16853 12699 16911 12705
rect 16853 12696 16865 12699
rect 15988 12668 16865 12696
rect 15988 12656 15994 12668
rect 16853 12665 16865 12668
rect 16899 12696 16911 12699
rect 17034 12696 17040 12708
rect 16899 12668 17040 12696
rect 16899 12665 16911 12668
rect 16853 12659 16911 12665
rect 17034 12656 17040 12668
rect 17092 12656 17098 12708
rect 17865 12699 17923 12705
rect 17865 12665 17877 12699
rect 17911 12696 17923 12699
rect 18414 12696 18420 12708
rect 17911 12668 18420 12696
rect 17911 12665 17923 12668
rect 17865 12659 17923 12665
rect 18414 12656 18420 12668
rect 18472 12696 18478 12708
rect 18598 12696 18604 12708
rect 18472 12668 18604 12696
rect 18472 12656 18478 12668
rect 18598 12656 18604 12668
rect 18656 12696 18662 12708
rect 21174 12705 21180 12708
rect 19245 12699 19303 12705
rect 19245 12696 19257 12699
rect 18656 12668 19257 12696
rect 18656 12656 18662 12668
rect 19245 12665 19257 12668
rect 19291 12665 19303 12699
rect 19245 12659 19303 12665
rect 20717 12699 20775 12705
rect 20717 12665 20729 12699
rect 20763 12696 20775 12699
rect 21130 12699 21180 12705
rect 21130 12696 21142 12699
rect 20763 12668 21142 12696
rect 20763 12665 20775 12668
rect 20717 12659 20775 12665
rect 21130 12665 21142 12668
rect 21176 12665 21180 12699
rect 21130 12659 21180 12665
rect 21174 12656 21180 12659
rect 21232 12696 21238 12708
rect 21232 12668 21278 12696
rect 21232 12656 21238 12668
rect 22002 12656 22008 12708
rect 22060 12696 22066 12708
rect 22186 12696 22192 12708
rect 22060 12668 22192 12696
rect 22060 12656 22066 12668
rect 22186 12656 22192 12668
rect 22244 12656 22250 12708
rect 24946 12656 24952 12708
rect 25004 12696 25010 12708
rect 25179 12699 25237 12705
rect 25179 12696 25191 12699
rect 25004 12668 25191 12696
rect 25004 12656 25010 12668
rect 25179 12665 25191 12668
rect 25225 12665 25237 12699
rect 25179 12659 25237 12665
rect 16390 12628 16396 12640
rect 15764 12600 16396 12628
rect 16390 12588 16396 12600
rect 16448 12588 16454 12640
rect 17218 12628 17224 12640
rect 17179 12600 17224 12628
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 18506 12588 18512 12640
rect 18564 12628 18570 12640
rect 19935 12631 19993 12637
rect 19935 12628 19947 12631
rect 18564 12600 19947 12628
rect 18564 12588 18570 12600
rect 19935 12597 19947 12600
rect 19981 12597 19993 12631
rect 19935 12591 19993 12597
rect 21729 12631 21787 12637
rect 21729 12597 21741 12631
rect 21775 12628 21787 12631
rect 22278 12628 22284 12640
rect 21775 12600 22284 12628
rect 21775 12597 21787 12600
rect 21729 12591 21787 12597
rect 22278 12588 22284 12600
rect 22336 12588 22342 12640
rect 22738 12637 22744 12640
rect 22695 12631 22744 12637
rect 22695 12597 22707 12631
rect 22741 12597 22744 12631
rect 22695 12591 22744 12597
rect 22738 12588 22744 12591
rect 22796 12588 22802 12640
rect 23290 12588 23296 12640
rect 23348 12628 23354 12640
rect 24167 12631 24225 12637
rect 24167 12628 24179 12631
rect 23348 12600 24179 12628
rect 23348 12588 23354 12600
rect 24167 12597 24179 12600
rect 24213 12597 24225 12631
rect 24167 12591 24225 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 3881 12427 3939 12433
rect 3881 12393 3893 12427
rect 3927 12424 3939 12427
rect 3970 12424 3976 12436
rect 3927 12396 3976 12424
rect 3927 12393 3939 12396
rect 3881 12387 3939 12393
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4154 12424 4160 12436
rect 4115 12396 4160 12424
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 4338 12384 4344 12436
rect 4396 12424 4402 12436
rect 9030 12424 9036 12436
rect 4396 12396 9036 12424
rect 4396 12384 4402 12396
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9950 12424 9956 12436
rect 9911 12396 9956 12424
rect 9950 12384 9956 12396
rect 10008 12384 10014 12436
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 10192 12396 10241 12424
rect 10192 12384 10198 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 10229 12387 10287 12393
rect 12437 12427 12495 12433
rect 12437 12393 12449 12427
rect 12483 12424 12495 12427
rect 12618 12424 12624 12436
rect 12483 12396 12624 12424
rect 12483 12393 12495 12396
rect 12437 12387 12495 12393
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 13449 12427 13507 12433
rect 13449 12393 13461 12427
rect 13495 12424 13507 12427
rect 13722 12424 13728 12436
rect 13495 12396 13728 12424
rect 13495 12393 13507 12396
rect 13449 12387 13507 12393
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 16390 12424 16396 12436
rect 16351 12396 16396 12424
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 18046 12384 18052 12436
rect 18104 12424 18110 12436
rect 18141 12427 18199 12433
rect 18141 12424 18153 12427
rect 18104 12396 18153 12424
rect 18104 12384 18110 12396
rect 18141 12393 18153 12396
rect 18187 12393 18199 12427
rect 18506 12424 18512 12436
rect 18467 12396 18512 12424
rect 18141 12387 18199 12393
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 21821 12427 21879 12433
rect 21821 12393 21833 12427
rect 21867 12424 21879 12427
rect 22002 12424 22008 12436
rect 21867 12396 22008 12424
rect 21867 12393 21879 12396
rect 21821 12387 21879 12393
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 22186 12384 22192 12436
rect 22244 12424 22250 12436
rect 22462 12424 22468 12436
rect 22244 12396 22468 12424
rect 22244 12384 22250 12396
rect 22462 12384 22468 12396
rect 22520 12384 22526 12436
rect 24118 12384 24124 12436
rect 24176 12424 24182 12436
rect 24305 12427 24363 12433
rect 24305 12424 24317 12427
rect 24176 12396 24317 12424
rect 24176 12384 24182 12396
rect 24305 12393 24317 12396
rect 24351 12393 24363 12427
rect 24305 12387 24363 12393
rect 3145 12359 3203 12365
rect 3145 12325 3157 12359
rect 3191 12356 3203 12359
rect 3326 12356 3332 12368
rect 3191 12328 3332 12356
rect 3191 12325 3203 12328
rect 3145 12319 3203 12325
rect 3326 12316 3332 12328
rect 3384 12316 3390 12368
rect 6270 12356 6276 12368
rect 5920 12328 6276 12356
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 1486 12288 1492 12300
rect 1443 12260 1492 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 1486 12248 1492 12260
rect 1544 12248 1550 12300
rect 2314 12248 2320 12300
rect 2372 12288 2378 12300
rect 2409 12291 2467 12297
rect 2409 12288 2421 12291
rect 2372 12260 2421 12288
rect 2372 12248 2378 12260
rect 2409 12257 2421 12260
rect 2455 12257 2467 12291
rect 2866 12288 2872 12300
rect 2827 12260 2872 12288
rect 2409 12251 2467 12257
rect 2866 12248 2872 12260
rect 2924 12248 2930 12300
rect 2958 12248 2964 12300
rect 3016 12288 3022 12300
rect 3878 12288 3884 12300
rect 3016 12260 3884 12288
rect 3016 12248 3022 12260
rect 3878 12248 3884 12260
rect 3936 12288 3942 12300
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 3936 12260 4077 12288
rect 3936 12248 3942 12260
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 4065 12251 4123 12257
rect 4246 12248 4252 12300
rect 4304 12288 4310 12300
rect 5920 12297 5948 12328
rect 6270 12316 6276 12328
rect 6328 12316 6334 12368
rect 8757 12359 8815 12365
rect 8757 12325 8769 12359
rect 8803 12356 8815 12359
rect 9674 12356 9680 12368
rect 8803 12328 9680 12356
rect 8803 12325 8815 12328
rect 8757 12319 8815 12325
rect 9674 12316 9680 12328
rect 9732 12316 9738 12368
rect 9766 12316 9772 12368
rect 9824 12356 9830 12368
rect 10594 12356 10600 12368
rect 9824 12328 10600 12356
rect 9824 12316 9830 12328
rect 10594 12316 10600 12328
rect 10652 12316 10658 12368
rect 10689 12359 10747 12365
rect 10689 12325 10701 12359
rect 10735 12356 10747 12359
rect 10870 12356 10876 12368
rect 10735 12328 10876 12356
rect 10735 12325 10747 12328
rect 10689 12319 10747 12325
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 12891 12359 12949 12365
rect 12891 12325 12903 12359
rect 12937 12356 12949 12359
rect 12986 12356 12992 12368
rect 12937 12328 12992 12356
rect 12937 12325 12949 12328
rect 12891 12319 12949 12325
rect 12986 12316 12992 12328
rect 13044 12316 13050 12368
rect 15378 12316 15384 12368
rect 15436 12356 15442 12368
rect 15473 12359 15531 12365
rect 15473 12356 15485 12359
rect 15436 12328 15485 12356
rect 15436 12316 15442 12328
rect 15473 12325 15485 12328
rect 15519 12325 15531 12359
rect 16022 12356 16028 12368
rect 15983 12328 16028 12356
rect 15473 12319 15531 12325
rect 16022 12316 16028 12328
rect 16080 12316 16086 12368
rect 16206 12316 16212 12368
rect 16264 12356 16270 12368
rect 16850 12356 16856 12368
rect 16264 12328 16856 12356
rect 16264 12316 16270 12328
rect 16850 12316 16856 12328
rect 16908 12316 16914 12368
rect 17402 12316 17408 12368
rect 17460 12356 17466 12368
rect 17583 12359 17641 12365
rect 17583 12356 17595 12359
rect 17460 12328 17595 12356
rect 17460 12316 17466 12328
rect 17583 12325 17595 12328
rect 17629 12356 17641 12359
rect 18874 12356 18880 12368
rect 17629 12328 18880 12356
rect 17629 12325 17641 12328
rect 17583 12319 17641 12325
rect 18874 12316 18880 12328
rect 18932 12316 18938 12368
rect 19429 12359 19487 12365
rect 19429 12325 19441 12359
rect 19475 12356 19487 12359
rect 19610 12356 19616 12368
rect 19475 12328 19616 12356
rect 19475 12325 19487 12328
rect 19429 12319 19487 12325
rect 19610 12316 19616 12328
rect 19668 12316 19674 12368
rect 19981 12359 20039 12365
rect 19981 12325 19993 12359
rect 20027 12356 20039 12359
rect 20530 12356 20536 12368
rect 20027 12328 20536 12356
rect 20027 12325 20039 12328
rect 19981 12319 20039 12325
rect 20530 12316 20536 12328
rect 20588 12316 20594 12368
rect 21174 12316 21180 12368
rect 21232 12365 21238 12368
rect 21232 12359 21280 12365
rect 21232 12325 21234 12359
rect 21268 12325 21280 12359
rect 21232 12319 21280 12325
rect 21232 12316 21238 12319
rect 22278 12316 22284 12368
rect 22336 12356 22342 12368
rect 22833 12359 22891 12365
rect 22833 12356 22845 12359
rect 22336 12328 22845 12356
rect 22336 12316 22342 12328
rect 22833 12325 22845 12328
rect 22879 12356 22891 12359
rect 23198 12356 23204 12368
rect 22879 12328 23204 12356
rect 22879 12325 22891 12328
rect 22833 12319 22891 12325
rect 23198 12316 23204 12328
rect 23256 12316 23262 12368
rect 4617 12291 4675 12297
rect 4617 12288 4629 12291
rect 4304 12260 4629 12288
rect 4304 12248 4310 12260
rect 4617 12257 4629 12260
rect 4663 12257 4675 12291
rect 4617 12251 4675 12257
rect 5905 12291 5963 12297
rect 5905 12257 5917 12291
rect 5951 12257 5963 12291
rect 6086 12288 6092 12300
rect 6047 12260 6092 12288
rect 5905 12251 5963 12257
rect 4632 12220 4660 12251
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 8297 12291 8355 12297
rect 8297 12288 8309 12291
rect 7064 12260 8309 12288
rect 7064 12248 7070 12260
rect 8297 12257 8309 12260
rect 8343 12257 8355 12291
rect 8570 12288 8576 12300
rect 8483 12260 8576 12288
rect 8297 12251 8355 12257
rect 6104 12220 6132 12248
rect 4632 12192 6132 12220
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 6822 12220 6828 12232
rect 6411 12192 6828 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 6822 12180 6828 12192
rect 6880 12220 6886 12232
rect 7193 12223 7251 12229
rect 7193 12220 7205 12223
rect 6880 12192 7205 12220
rect 6880 12180 6886 12192
rect 7193 12189 7205 12192
rect 7239 12189 7251 12223
rect 8312 12220 8340 12251
rect 8570 12248 8576 12260
rect 8628 12288 8634 12300
rect 9582 12288 9588 12300
rect 8628 12260 9588 12288
rect 8628 12248 8634 12260
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 18138 12248 18144 12300
rect 18196 12288 18202 12300
rect 18785 12291 18843 12297
rect 18785 12288 18797 12291
rect 18196 12260 18797 12288
rect 18196 12248 18202 12260
rect 18785 12257 18797 12260
rect 18831 12257 18843 12291
rect 18785 12251 18843 12257
rect 22094 12248 22100 12300
rect 22152 12288 22158 12300
rect 24489 12291 24547 12297
rect 22152 12260 22197 12288
rect 22152 12248 22158 12260
rect 24489 12257 24501 12291
rect 24535 12288 24547 12291
rect 24578 12288 24584 12300
rect 24535 12260 24584 12288
rect 24535 12257 24547 12260
rect 24489 12251 24547 12257
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 24765 12291 24823 12297
rect 24765 12257 24777 12291
rect 24811 12288 24823 12291
rect 25130 12288 25136 12300
rect 24811 12260 25136 12288
rect 24811 12257 24823 12260
rect 24765 12251 24823 12257
rect 25130 12248 25136 12260
rect 25188 12248 25194 12300
rect 8938 12220 8944 12232
rect 8312 12192 8944 12220
rect 7193 12183 7251 12189
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 12492 12192 12541 12220
rect 12492 12180 12498 12192
rect 12529 12189 12541 12192
rect 12575 12220 12587 12223
rect 13078 12220 13084 12232
rect 12575 12192 13084 12220
rect 12575 12189 12587 12192
rect 12529 12183 12587 12189
rect 13078 12180 13084 12192
rect 13136 12180 13142 12232
rect 14090 12180 14096 12232
rect 14148 12220 14154 12232
rect 14734 12220 14740 12232
rect 14148 12192 14740 12220
rect 14148 12180 14154 12192
rect 14734 12180 14740 12192
rect 14792 12220 14798 12232
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 14792 12192 15393 12220
rect 14792 12180 14798 12192
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 17221 12223 17279 12229
rect 17221 12189 17233 12223
rect 17267 12220 17279 12223
rect 17678 12220 17684 12232
rect 17267 12192 17684 12220
rect 17267 12189 17279 12192
rect 17221 12183 17279 12189
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 19334 12220 19340 12232
rect 19295 12192 19340 12220
rect 19334 12180 19340 12192
rect 19392 12180 19398 12232
rect 20901 12223 20959 12229
rect 20901 12189 20913 12223
rect 20947 12220 20959 12223
rect 20990 12220 20996 12232
rect 20947 12192 20996 12220
rect 20947 12189 20959 12192
rect 20901 12183 20959 12189
rect 20990 12180 20996 12192
rect 21048 12180 21054 12232
rect 22738 12220 22744 12232
rect 22699 12192 22744 12220
rect 22738 12180 22744 12192
rect 22796 12180 22802 12232
rect 23014 12220 23020 12232
rect 22975 12192 23020 12220
rect 23014 12180 23020 12192
rect 23072 12180 23078 12232
rect 23750 12180 23756 12232
rect 23808 12180 23814 12232
rect 1581 12155 1639 12161
rect 1581 12121 1593 12155
rect 1627 12152 1639 12155
rect 4706 12152 4712 12164
rect 1627 12124 4712 12152
rect 1627 12121 1639 12124
rect 1581 12115 1639 12121
rect 4706 12112 4712 12124
rect 4764 12112 4770 12164
rect 10778 12112 10784 12164
rect 10836 12152 10842 12164
rect 11054 12152 11060 12164
rect 10836 12124 11060 12152
rect 10836 12112 10842 12124
rect 11054 12112 11060 12124
rect 11112 12152 11118 12164
rect 11149 12155 11207 12161
rect 11149 12152 11161 12155
rect 11112 12124 11161 12152
rect 11112 12112 11118 12124
rect 11149 12121 11161 12124
rect 11195 12121 11207 12155
rect 11149 12115 11207 12121
rect 20530 12112 20536 12164
rect 20588 12152 20594 12164
rect 21174 12152 21180 12164
rect 20588 12124 21180 12152
rect 20588 12112 20594 12124
rect 21174 12112 21180 12124
rect 21232 12112 21238 12164
rect 23768 12152 23796 12180
rect 23032 12124 23796 12152
rect 23032 12096 23060 12124
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 2317 12087 2375 12093
rect 2317 12053 2329 12087
rect 2363 12084 2375 12087
rect 2406 12084 2412 12096
rect 2363 12056 2412 12084
rect 2363 12053 2375 12056
rect 2317 12047 2375 12053
rect 2406 12044 2412 12056
rect 2464 12044 2470 12096
rect 4614 12044 4620 12096
rect 4672 12084 4678 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 4672 12056 5089 12084
rect 4672 12044 4678 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 5077 12047 5135 12053
rect 6917 12087 6975 12093
rect 6917 12053 6929 12087
rect 6963 12084 6975 12087
rect 7098 12084 7104 12096
rect 6963 12056 7104 12084
rect 6963 12053 6975 12056
rect 6917 12047 6975 12053
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 7929 12087 7987 12093
rect 7929 12053 7941 12087
rect 7975 12084 7987 12087
rect 8018 12084 8024 12096
rect 7975 12056 8024 12084
rect 7975 12053 7987 12056
rect 7929 12047 7987 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 14090 12084 14096 12096
rect 14051 12056 14096 12084
rect 14090 12044 14096 12056
rect 14148 12044 14154 12096
rect 19150 12044 19156 12096
rect 19208 12084 19214 12096
rect 20254 12084 20260 12096
rect 19208 12056 20260 12084
rect 19208 12044 19214 12056
rect 20254 12044 20260 12056
rect 20312 12044 20318 12096
rect 20714 12084 20720 12096
rect 20627 12056 20720 12084
rect 20714 12044 20720 12056
rect 20772 12084 20778 12096
rect 22094 12084 22100 12096
rect 20772 12056 22100 12084
rect 20772 12044 20778 12056
rect 22094 12044 22100 12056
rect 22152 12044 22158 12096
rect 23014 12044 23020 12096
rect 23072 12044 23078 12096
rect 23658 12084 23664 12096
rect 23619 12056 23664 12084
rect 23658 12044 23664 12056
rect 23716 12044 23722 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1486 11840 1492 11892
rect 1544 11880 1550 11892
rect 1673 11883 1731 11889
rect 1673 11880 1685 11883
rect 1544 11852 1685 11880
rect 1544 11840 1550 11852
rect 1673 11849 1685 11852
rect 1719 11880 1731 11883
rect 2958 11880 2964 11892
rect 1719 11852 2964 11880
rect 1719 11849 1731 11852
rect 1673 11843 1731 11849
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 3237 11883 3295 11889
rect 3237 11849 3249 11883
rect 3283 11880 3295 11883
rect 3602 11880 3608 11892
rect 3283 11852 3608 11880
rect 3283 11849 3295 11852
rect 3237 11843 3295 11849
rect 2038 11772 2044 11824
rect 2096 11812 2102 11824
rect 2501 11815 2559 11821
rect 2501 11812 2513 11815
rect 2096 11784 2513 11812
rect 2096 11772 2102 11784
rect 2501 11781 2513 11784
rect 2547 11781 2559 11815
rect 2501 11775 2559 11781
rect 1302 11704 1308 11756
rect 1360 11744 1366 11756
rect 1486 11744 1492 11756
rect 1360 11716 1492 11744
rect 1360 11704 1366 11716
rect 1486 11704 1492 11716
rect 1544 11704 1550 11756
rect 1578 11704 1584 11756
rect 1636 11744 1642 11756
rect 3344 11744 3372 11852
rect 3602 11840 3608 11852
rect 3660 11840 3666 11892
rect 3878 11880 3884 11892
rect 3839 11852 3884 11880
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 5721 11883 5779 11889
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 6270 11880 6276 11892
rect 5767 11852 6276 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 7745 11883 7803 11889
rect 7745 11849 7757 11883
rect 7791 11880 7803 11883
rect 8570 11880 8576 11892
rect 7791 11852 8576 11880
rect 7791 11849 7803 11852
rect 7745 11843 7803 11849
rect 6086 11812 6092 11824
rect 5999 11784 6092 11812
rect 6086 11772 6092 11784
rect 6144 11812 6150 11824
rect 7760 11812 7788 11843
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 11149 11883 11207 11889
rect 11149 11880 11161 11883
rect 10652 11852 11161 11880
rect 10652 11840 10658 11852
rect 11149 11849 11161 11852
rect 11195 11849 11207 11883
rect 11149 11843 11207 11849
rect 16945 11883 17003 11889
rect 16945 11849 16957 11883
rect 16991 11880 17003 11883
rect 17310 11880 17316 11892
rect 16991 11852 17316 11880
rect 16991 11849 17003 11852
rect 16945 11843 17003 11849
rect 8938 11812 8944 11824
rect 6144 11784 7788 11812
rect 8899 11784 8944 11812
rect 6144 11772 6150 11784
rect 8938 11772 8944 11784
rect 8996 11772 9002 11824
rect 16960 11812 16988 11843
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 18785 11883 18843 11889
rect 18785 11849 18797 11883
rect 18831 11880 18843 11883
rect 18874 11880 18880 11892
rect 18831 11852 18880 11880
rect 18831 11849 18843 11852
rect 18785 11843 18843 11849
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 21542 11840 21548 11892
rect 21600 11880 21606 11892
rect 21637 11883 21695 11889
rect 21637 11880 21649 11883
rect 21600 11852 21649 11880
rect 21600 11840 21606 11852
rect 21637 11849 21649 11852
rect 21683 11849 21695 11883
rect 21637 11843 21695 11849
rect 22278 11840 22284 11892
rect 22336 11880 22342 11892
rect 22603 11883 22661 11889
rect 22603 11880 22615 11883
rect 22336 11852 22615 11880
rect 22336 11840 22342 11852
rect 22603 11849 22615 11852
rect 22649 11849 22661 11883
rect 25406 11880 25412 11892
rect 25367 11852 25412 11880
rect 22603 11843 22661 11849
rect 25406 11840 25412 11852
rect 25464 11840 25470 11892
rect 15948 11784 16988 11812
rect 18417 11815 18475 11821
rect 1636 11716 3372 11744
rect 1636 11704 1642 11716
rect 3344 11685 3372 11716
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11744 4307 11747
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 4295 11716 4445 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 4433 11713 4445 11716
rect 4479 11744 4491 11747
rect 4522 11744 4528 11756
rect 4479 11716 4528 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 4522 11704 4528 11716
rect 4580 11704 4586 11756
rect 7190 11704 7196 11756
rect 7248 11744 7254 11756
rect 7929 11747 7987 11753
rect 7929 11744 7941 11747
rect 7248 11716 7941 11744
rect 7248 11704 7254 11716
rect 7929 11713 7941 11716
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 8573 11747 8631 11753
rect 8573 11713 8585 11747
rect 8619 11744 8631 11747
rect 8662 11744 8668 11756
rect 8619 11716 8668 11744
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11744 9643 11747
rect 9950 11744 9956 11756
rect 9631 11716 9956 11744
rect 9631 11713 9643 11716
rect 9585 11707 9643 11713
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 15378 11744 15384 11756
rect 13556 11716 15384 11744
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11676 2375 11679
rect 3329 11679 3387 11685
rect 2363 11648 2636 11676
rect 2363 11645 2375 11648
rect 2317 11639 2375 11645
rect 2225 11543 2283 11549
rect 2225 11509 2237 11543
rect 2271 11540 2283 11543
rect 2314 11540 2320 11552
rect 2271 11512 2320 11540
rect 2271 11509 2283 11512
rect 2225 11503 2283 11509
rect 2314 11500 2320 11512
rect 2372 11500 2378 11552
rect 2608 11540 2636 11648
rect 3329 11645 3341 11679
rect 3375 11645 3387 11679
rect 3329 11639 3387 11645
rect 4062 11636 4068 11688
rect 4120 11676 4126 11688
rect 4341 11679 4399 11685
rect 4341 11676 4353 11679
rect 4120 11648 4353 11676
rect 4120 11636 4126 11648
rect 4341 11645 4353 11648
rect 4387 11645 4399 11679
rect 4614 11676 4620 11688
rect 4575 11648 4620 11676
rect 4341 11639 4399 11645
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 6822 11676 6828 11688
rect 6783 11648 6828 11676
rect 6822 11636 6828 11648
rect 6880 11676 6886 11688
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 6880 11648 7297 11676
rect 6880 11636 6886 11648
rect 7285 11645 7297 11648
rect 7331 11645 7343 11679
rect 7285 11639 7343 11645
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11333 11679 11391 11685
rect 11333 11676 11345 11679
rect 11112 11648 11345 11676
rect 11112 11636 11118 11648
rect 11333 11645 11345 11648
rect 11379 11676 11391 11679
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 11379 11648 11805 11676
rect 11379 11645 11391 11648
rect 11333 11639 11391 11645
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 12526 11676 12532 11688
rect 12487 11648 12532 11676
rect 11793 11639 11851 11645
rect 12526 11636 12532 11648
rect 12584 11636 12590 11688
rect 12986 11676 12992 11688
rect 12947 11648 12992 11676
rect 12986 11636 12992 11648
rect 13044 11676 13050 11688
rect 13556 11685 13584 11716
rect 15378 11704 15384 11716
rect 15436 11704 15442 11756
rect 15948 11753 15976 11784
rect 18417 11781 18429 11815
rect 18463 11812 18475 11815
rect 19610 11812 19616 11824
rect 18463 11784 19616 11812
rect 18463 11781 18475 11784
rect 18417 11775 18475 11781
rect 19610 11772 19616 11784
rect 19668 11812 19674 11824
rect 19797 11815 19855 11821
rect 19797 11812 19809 11815
rect 19668 11784 19809 11812
rect 19668 11772 19674 11784
rect 19797 11781 19809 11784
rect 19843 11781 19855 11815
rect 19797 11775 19855 11781
rect 22373 11815 22431 11821
rect 22373 11781 22385 11815
rect 22419 11812 22431 11815
rect 23198 11812 23204 11824
rect 22419 11784 23204 11812
rect 22419 11781 22431 11784
rect 22373 11775 22431 11781
rect 23198 11772 23204 11784
rect 23256 11772 23262 11824
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16022 11704 16028 11756
rect 16080 11744 16086 11756
rect 16209 11747 16267 11753
rect 16209 11744 16221 11747
rect 16080 11716 16221 11744
rect 16080 11704 16086 11716
rect 16209 11713 16221 11716
rect 16255 11713 16267 11747
rect 16209 11707 16267 11713
rect 17313 11747 17371 11753
rect 17313 11713 17325 11747
rect 17359 11744 17371 11747
rect 17402 11744 17408 11756
rect 17359 11716 17408 11744
rect 17359 11713 17371 11716
rect 17313 11707 17371 11713
rect 17402 11704 17408 11716
rect 17460 11704 17466 11756
rect 20714 11704 20720 11756
rect 20772 11744 20778 11756
rect 20772 11716 20817 11744
rect 20772 11704 20778 11716
rect 20990 11704 20996 11756
rect 21048 11744 21054 11756
rect 21913 11747 21971 11753
rect 21913 11744 21925 11747
rect 21048 11716 21925 11744
rect 21048 11704 21054 11716
rect 21913 11713 21925 11716
rect 21959 11713 21971 11747
rect 21913 11707 21971 11713
rect 13541 11679 13599 11685
rect 13541 11676 13553 11679
rect 13044 11648 13553 11676
rect 13044 11636 13050 11648
rect 13541 11645 13553 11648
rect 13587 11645 13599 11679
rect 14090 11676 14096 11688
rect 14051 11648 14096 11676
rect 13541 11639 13599 11645
rect 14090 11636 14096 11648
rect 14148 11636 14154 11688
rect 15013 11679 15071 11685
rect 15013 11645 15025 11679
rect 15059 11676 15071 11679
rect 15657 11679 15715 11685
rect 15657 11676 15669 11679
rect 15059 11648 15669 11676
rect 15059 11645 15071 11648
rect 15013 11639 15071 11645
rect 15657 11645 15669 11648
rect 15703 11645 15715 11679
rect 18874 11676 18880 11688
rect 18835 11648 18880 11676
rect 15657 11639 15715 11645
rect 5074 11608 5080 11620
rect 3436 11580 5080 11608
rect 2869 11543 2927 11549
rect 2869 11540 2881 11543
rect 2608 11512 2881 11540
rect 2869 11509 2881 11512
rect 2915 11540 2927 11543
rect 3436 11540 3464 11580
rect 5074 11568 5080 11580
rect 5132 11568 5138 11620
rect 8018 11568 8024 11620
rect 8076 11608 8082 11620
rect 9858 11608 9864 11620
rect 8076 11580 8121 11608
rect 9816 11580 9864 11608
rect 8076 11568 8082 11580
rect 9858 11568 9864 11580
rect 9916 11617 9922 11620
rect 9916 11611 9964 11617
rect 9916 11577 9918 11611
rect 9952 11608 9964 11611
rect 12161 11611 12219 11617
rect 12161 11608 12173 11611
rect 9952 11580 12173 11608
rect 9952 11577 9964 11580
rect 9916 11571 9964 11577
rect 12161 11577 12173 11580
rect 12207 11577 12219 11611
rect 13262 11608 13268 11620
rect 13223 11580 13268 11608
rect 12161 11571 12219 11577
rect 9916 11568 9949 11571
rect 2915 11512 3464 11540
rect 3513 11543 3571 11549
rect 2915 11509 2927 11512
rect 2869 11503 2927 11509
rect 3513 11509 3525 11543
rect 3559 11540 3571 11543
rect 3970 11540 3976 11552
rect 3559 11512 3976 11540
rect 3559 11509 3571 11512
rect 3513 11503 3571 11509
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 7006 11540 7012 11552
rect 6967 11512 7012 11540
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 7742 11540 7748 11552
rect 7616 11512 7748 11540
rect 7616 11500 7622 11512
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 9398 11540 9404 11552
rect 9359 11512 9404 11540
rect 9398 11500 9404 11512
rect 9456 11540 9462 11552
rect 9921 11540 9949 11568
rect 9456 11512 9949 11540
rect 10505 11543 10563 11549
rect 9456 11500 9462 11512
rect 10505 11509 10517 11543
rect 10551 11540 10563 11543
rect 10870 11540 10876 11552
rect 10551 11512 10876 11540
rect 10551 11509 10563 11512
rect 10505 11503 10563 11509
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 11514 11540 11520 11552
rect 11475 11512 11520 11540
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 12176 11540 12204 11571
rect 13262 11568 13268 11580
rect 13320 11568 13326 11620
rect 14414 11611 14472 11617
rect 14414 11577 14426 11611
rect 14460 11577 14472 11611
rect 14414 11571 14472 11577
rect 13722 11540 13728 11552
rect 12176 11512 13728 11540
rect 13722 11500 13728 11512
rect 13780 11540 13786 11552
rect 13909 11543 13967 11549
rect 13909 11540 13921 11543
rect 13780 11512 13921 11540
rect 13780 11500 13786 11512
rect 13909 11509 13921 11512
rect 13955 11540 13967 11543
rect 14429 11540 14457 11571
rect 15286 11540 15292 11552
rect 13955 11512 14457 11540
rect 15247 11512 15292 11540
rect 13955 11509 13967 11512
rect 13909 11503 13967 11509
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 15672 11540 15700 11639
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 22462 11636 22468 11688
rect 22520 11685 22526 11688
rect 22520 11679 22558 11685
rect 22546 11676 22558 11679
rect 22925 11679 22983 11685
rect 22925 11676 22937 11679
rect 22546 11648 22937 11676
rect 22546 11645 22558 11648
rect 22520 11639 22558 11645
rect 22925 11645 22937 11648
rect 22971 11645 22983 11679
rect 22925 11639 22983 11645
rect 22520 11636 22526 11639
rect 23658 11636 23664 11688
rect 23716 11676 23722 11688
rect 23753 11679 23811 11685
rect 23753 11676 23765 11679
rect 23716 11648 23765 11676
rect 23716 11636 23722 11648
rect 23753 11645 23765 11648
rect 23799 11645 23811 11679
rect 23753 11639 23811 11645
rect 23842 11636 23848 11688
rect 23900 11676 23906 11688
rect 24121 11679 24179 11685
rect 24121 11676 24133 11679
rect 23900 11648 24133 11676
rect 23900 11636 23906 11648
rect 24121 11645 24133 11648
rect 24167 11645 24179 11679
rect 24121 11639 24179 11645
rect 25225 11679 25283 11685
rect 25225 11645 25237 11679
rect 25271 11676 25283 11679
rect 25314 11676 25320 11688
rect 25271 11648 25320 11676
rect 25271 11645 25283 11648
rect 25225 11639 25283 11645
rect 25314 11636 25320 11648
rect 25372 11676 25378 11688
rect 25777 11679 25835 11685
rect 25777 11676 25789 11679
rect 25372 11648 25789 11676
rect 25372 11636 25378 11648
rect 25777 11645 25789 11648
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 16025 11611 16083 11617
rect 16025 11577 16037 11611
rect 16071 11577 16083 11611
rect 16025 11571 16083 11577
rect 16040 11540 16068 11571
rect 18966 11568 18972 11620
rect 19024 11608 19030 11620
rect 19198 11611 19256 11617
rect 19198 11608 19210 11611
rect 19024 11580 19210 11608
rect 19024 11568 19030 11580
rect 19198 11577 19210 11580
rect 19244 11608 19256 11611
rect 20165 11611 20223 11617
rect 20165 11608 20177 11611
rect 19244 11580 20177 11608
rect 19244 11577 19256 11580
rect 19198 11571 19256 11577
rect 20165 11577 20177 11580
rect 20211 11608 20223 11611
rect 20530 11608 20536 11620
rect 20211 11580 20536 11608
rect 20211 11577 20223 11580
rect 20165 11571 20223 11577
rect 20530 11568 20536 11580
rect 20588 11608 20594 11620
rect 21038 11611 21096 11617
rect 21038 11608 21050 11611
rect 20588 11580 21050 11608
rect 20588 11568 20594 11580
rect 21038 11577 21050 11580
rect 21084 11608 21096 11611
rect 21084 11580 22048 11608
rect 21084 11577 21096 11580
rect 21038 11571 21096 11577
rect 22020 11552 22048 11580
rect 23290 11568 23296 11620
rect 23348 11608 23354 11620
rect 24670 11608 24676 11620
rect 23348 11580 24676 11608
rect 23348 11568 23354 11580
rect 24670 11568 24676 11580
rect 24728 11568 24734 11620
rect 17678 11540 17684 11552
rect 15672 11512 16068 11540
rect 17639 11512 17684 11540
rect 17678 11500 17684 11512
rect 17736 11500 17742 11552
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 21358 11540 21364 11552
rect 20864 11512 21364 11540
rect 20864 11500 20870 11512
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 22002 11500 22008 11552
rect 22060 11500 22066 11552
rect 23198 11500 23204 11552
rect 23256 11540 23262 11552
rect 23385 11543 23443 11549
rect 23385 11540 23397 11543
rect 23256 11512 23397 11540
rect 23256 11500 23262 11512
rect 23385 11509 23397 11512
rect 23431 11509 23443 11543
rect 23750 11540 23756 11552
rect 23711 11512 23756 11540
rect 23385 11503 23443 11509
rect 23750 11500 23756 11512
rect 23808 11500 23814 11552
rect 25130 11540 25136 11552
rect 25043 11512 25136 11540
rect 25130 11500 25136 11512
rect 25188 11540 25194 11552
rect 25866 11540 25872 11552
rect 25188 11512 25872 11540
rect 25188 11500 25194 11512
rect 25866 11500 25872 11512
rect 25924 11500 25930 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2866 11336 2872 11348
rect 2363 11308 2872 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 4893 11339 4951 11345
rect 4893 11336 4905 11339
rect 4212 11308 4905 11336
rect 4212 11296 4218 11308
rect 4893 11305 4905 11308
rect 4939 11305 4951 11339
rect 4893 11299 4951 11305
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 7248 11308 7389 11336
rect 7248 11296 7254 11308
rect 7377 11305 7389 11308
rect 7423 11305 7435 11339
rect 7377 11299 7435 11305
rect 8018 11296 8024 11348
rect 8076 11336 8082 11348
rect 8481 11339 8539 11345
rect 8481 11336 8493 11339
rect 8076 11308 8493 11336
rect 8076 11296 8082 11308
rect 8481 11305 8493 11308
rect 8527 11305 8539 11339
rect 8481 11299 8539 11305
rect 12437 11339 12495 11345
rect 12437 11305 12449 11339
rect 12483 11305 12495 11339
rect 12437 11299 12495 11305
rect 2498 11228 2504 11280
rect 2556 11268 2562 11280
rect 3789 11271 3847 11277
rect 3789 11268 3801 11271
rect 2556 11240 3801 11268
rect 2556 11228 2562 11240
rect 3789 11237 3801 11240
rect 3835 11268 3847 11271
rect 4062 11268 4068 11280
rect 3835 11240 4068 11268
rect 3835 11237 3847 11240
rect 3789 11231 3847 11237
rect 4062 11228 4068 11240
rect 4120 11228 4126 11280
rect 4246 11268 4252 11280
rect 4207 11240 4252 11268
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 4356 11240 4660 11268
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 1578 11200 1584 11212
rect 1443 11172 1584 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 1578 11160 1584 11172
rect 1636 11200 1642 11212
rect 1762 11200 1768 11212
rect 1636 11172 1768 11200
rect 1636 11160 1642 11172
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 2409 11203 2467 11209
rect 2409 11169 2421 11203
rect 2455 11200 2467 11203
rect 2590 11200 2596 11212
rect 2455 11172 2596 11200
rect 2455 11169 2467 11172
rect 2409 11163 2467 11169
rect 2590 11160 2596 11172
rect 2648 11160 2654 11212
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 4356 11200 4384 11240
rect 4632 11212 4660 11240
rect 7098 11228 7104 11280
rect 7156 11268 7162 11280
rect 7650 11268 7656 11280
rect 7156 11240 7656 11268
rect 7156 11228 7162 11240
rect 7650 11228 7656 11240
rect 7708 11268 7714 11280
rect 7923 11271 7981 11277
rect 7923 11268 7935 11271
rect 7708 11240 7935 11268
rect 7708 11228 7714 11240
rect 7923 11237 7935 11240
rect 7969 11268 7981 11271
rect 9398 11268 9404 11280
rect 7969 11240 9404 11268
rect 7969 11237 7981 11240
rect 7923 11231 7981 11237
rect 9398 11228 9404 11240
rect 9456 11228 9462 11280
rect 10870 11268 10876 11280
rect 10831 11240 10876 11268
rect 10870 11228 10876 11240
rect 10928 11228 10934 11280
rect 12452 11268 12480 11299
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 12713 11339 12771 11345
rect 12713 11336 12725 11339
rect 12584 11308 12725 11336
rect 12584 11296 12590 11308
rect 12713 11305 12725 11308
rect 12759 11305 12771 11339
rect 13078 11336 13084 11348
rect 13039 11308 13084 11336
rect 12713 11299 12771 11305
rect 13078 11296 13084 11308
rect 13136 11296 13142 11348
rect 14277 11339 14335 11345
rect 14277 11305 14289 11339
rect 14323 11336 14335 11339
rect 15286 11336 15292 11348
rect 14323 11308 15292 11336
rect 14323 11305 14335 11308
rect 14277 11299 14335 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 18233 11339 18291 11345
rect 18233 11305 18245 11339
rect 18279 11336 18291 11339
rect 18414 11336 18420 11348
rect 18279 11308 18420 11336
rect 18279 11305 18291 11308
rect 18233 11299 18291 11305
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 18874 11336 18880 11348
rect 18835 11308 18880 11336
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 20990 11336 20996 11348
rect 20951 11308 20996 11336
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 22738 11336 22744 11348
rect 22699 11308 22744 11336
rect 22738 11296 22744 11308
rect 22796 11296 22802 11348
rect 23198 11296 23204 11348
rect 23256 11336 23262 11348
rect 23842 11336 23848 11348
rect 23256 11308 23848 11336
rect 23256 11296 23262 11308
rect 23842 11296 23848 11308
rect 23900 11296 23906 11348
rect 24946 11336 24952 11348
rect 24907 11308 24952 11336
rect 24946 11296 24952 11308
rect 25004 11296 25010 11348
rect 12802 11268 12808 11280
rect 12452 11240 12808 11268
rect 12802 11228 12808 11240
rect 12860 11228 12866 11280
rect 13722 11277 13728 11280
rect 13719 11268 13728 11277
rect 13683 11240 13728 11268
rect 13719 11231 13728 11240
rect 13722 11228 13728 11231
rect 13780 11228 13786 11280
rect 14826 11228 14832 11280
rect 14884 11268 14890 11280
rect 15562 11268 15568 11280
rect 14884 11240 15568 11268
rect 14884 11228 14890 11240
rect 15562 11228 15568 11240
rect 15620 11228 15626 11280
rect 15654 11228 15660 11280
rect 15712 11268 15718 11280
rect 15712 11240 15757 11268
rect 15712 11228 15718 11240
rect 17402 11228 17408 11280
rect 17460 11268 17466 11280
rect 17634 11271 17692 11277
rect 17634 11268 17646 11271
rect 17460 11240 17646 11268
rect 17460 11228 17466 11240
rect 17634 11237 17646 11240
rect 17680 11237 17692 11271
rect 17634 11231 17692 11237
rect 18601 11271 18659 11277
rect 18601 11237 18613 11271
rect 18647 11268 18659 11271
rect 19334 11268 19340 11280
rect 18647 11240 19340 11268
rect 18647 11237 18659 11240
rect 18601 11231 18659 11237
rect 19334 11228 19340 11240
rect 19392 11228 19398 11280
rect 19981 11271 20039 11277
rect 19981 11237 19993 11271
rect 20027 11268 20039 11271
rect 20622 11268 20628 11280
rect 20027 11240 20628 11268
rect 20027 11237 20039 11240
rect 19981 11231 20039 11237
rect 20622 11228 20628 11240
rect 20680 11228 20686 11280
rect 23382 11268 23388 11280
rect 23343 11240 23388 11268
rect 23382 11228 23388 11240
rect 23440 11228 23446 11280
rect 23474 11228 23480 11280
rect 23532 11268 23538 11280
rect 23532 11240 23577 11268
rect 23532 11228 23538 11240
rect 2731 11172 4384 11200
rect 4433 11203 4491 11209
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 4433 11169 4445 11203
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 2314 11092 2320 11144
rect 2372 11132 2378 11144
rect 2501 11135 2559 11141
rect 2501 11132 2513 11135
rect 2372 11104 2513 11132
rect 2372 11092 2378 11104
rect 2501 11101 2513 11104
rect 2547 11132 2559 11135
rect 2866 11132 2872 11144
rect 2547 11104 2703 11132
rect 2827 11104 2872 11132
rect 2547 11101 2559 11104
rect 2501 11095 2559 11101
rect 1578 11024 1584 11076
rect 1636 11064 1642 11076
rect 1857 11067 1915 11073
rect 1857 11064 1869 11067
rect 1636 11036 1869 11064
rect 1636 11024 1642 11036
rect 1857 11033 1869 11036
rect 1903 11033 1915 11067
rect 1857 11027 1915 11033
rect 2675 10996 2703 11104
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 3694 11092 3700 11144
rect 3752 11132 3758 11144
rect 4062 11132 4068 11144
rect 3752 11104 4068 11132
rect 3752 11092 3758 11104
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 4448 11132 4476 11163
rect 4614 11160 4620 11212
rect 4672 11200 4678 11212
rect 4709 11203 4767 11209
rect 4709 11200 4721 11203
rect 4672 11172 4721 11200
rect 4672 11160 4678 11172
rect 4709 11169 4721 11172
rect 4755 11169 4767 11203
rect 4709 11163 4767 11169
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 5997 11203 6055 11209
rect 5997 11200 6009 11203
rect 5316 11172 6009 11200
rect 5316 11160 5322 11172
rect 5997 11169 6009 11172
rect 6043 11200 6055 11203
rect 6362 11200 6368 11212
rect 6043 11172 6368 11200
rect 6043 11169 6055 11172
rect 5997 11163 6055 11169
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11200 6515 11203
rect 8386 11200 8392 11212
rect 6503 11172 8392 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 4798 11132 4804 11144
rect 4448 11104 4804 11132
rect 4798 11092 4804 11104
rect 4856 11092 4862 11144
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 6472 11132 6500 11163
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 9674 11200 9680 11212
rect 9635 11172 9680 11200
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 12253 11203 12311 11209
rect 12253 11200 12265 11203
rect 12124 11172 12265 11200
rect 12124 11160 12130 11172
rect 12253 11169 12265 11172
rect 12299 11169 12311 11203
rect 12253 11163 12311 11169
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 13357 11203 13415 11209
rect 13357 11200 13369 11203
rect 13320 11172 13369 11200
rect 13320 11160 13326 11172
rect 13357 11169 13369 11172
rect 13403 11169 13415 11203
rect 13357 11163 13415 11169
rect 14734 11160 14740 11212
rect 14792 11200 14798 11212
rect 15013 11203 15071 11209
rect 15013 11200 15025 11203
rect 14792 11172 15025 11200
rect 14792 11160 14798 11172
rect 15013 11169 15025 11172
rect 15059 11169 15071 11203
rect 17310 11200 17316 11212
rect 17271 11172 17316 11200
rect 15013 11163 15071 11169
rect 17310 11160 17316 11172
rect 17368 11160 17374 11212
rect 19426 11200 19432 11212
rect 19387 11172 19432 11200
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 19705 11203 19763 11209
rect 19705 11169 19717 11203
rect 19751 11169 19763 11203
rect 19705 11163 19763 11169
rect 5592 11104 6500 11132
rect 6733 11135 6791 11141
rect 5592 11092 5598 11104
rect 6733 11101 6745 11135
rect 6779 11132 6791 11135
rect 7190 11132 7196 11144
rect 6779 11104 7196 11132
rect 6779 11101 6791 11104
rect 6733 11095 6791 11101
rect 7190 11092 7196 11104
rect 7248 11132 7254 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7248 11104 7573 11132
rect 7248 11092 7254 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11101 10839 11135
rect 11054 11132 11060 11144
rect 11015 11104 11060 11132
rect 10781 11095 10839 11101
rect 4522 11064 4528 11076
rect 4483 11036 4528 11064
rect 4522 11024 4528 11036
rect 4580 11024 4586 11076
rect 9861 11067 9919 11073
rect 9861 11033 9873 11067
rect 9907 11064 9919 11067
rect 9950 11064 9956 11076
rect 9907 11036 9956 11064
rect 9907 11033 9919 11036
rect 9861 11027 9919 11033
rect 9950 11024 9956 11036
rect 10008 11024 10014 11076
rect 10796 11064 10824 11095
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 11238 11092 11244 11144
rect 11296 11132 11302 11144
rect 11422 11132 11428 11144
rect 11296 11104 11428 11132
rect 11296 11092 11302 11104
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12526 11132 12532 11144
rect 12207 11104 12532 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12526 11092 12532 11104
rect 12584 11092 12590 11144
rect 16022 11132 16028 11144
rect 15983 11104 16028 11132
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 19334 11092 19340 11144
rect 19392 11132 19398 11144
rect 19720 11132 19748 11163
rect 20530 11160 20536 11212
rect 20588 11200 20594 11212
rect 20901 11203 20959 11209
rect 20901 11200 20913 11203
rect 20588 11172 20913 11200
rect 20588 11160 20594 11172
rect 20901 11169 20913 11172
rect 20947 11169 20959 11203
rect 20901 11163 20959 11169
rect 21315 11203 21373 11209
rect 21315 11169 21327 11203
rect 21361 11169 21373 11203
rect 21315 11163 21373 11169
rect 24857 11203 24915 11209
rect 24857 11169 24869 11203
rect 24903 11169 24915 11203
rect 25317 11203 25375 11209
rect 25317 11200 25329 11203
rect 24857 11163 24915 11169
rect 24964 11172 25329 11200
rect 21330 11132 21358 11163
rect 23658 11132 23664 11144
rect 19392 11104 21358 11132
rect 23619 11104 23664 11132
rect 19392 11092 19398 11104
rect 21330 11064 21358 11104
rect 23658 11092 23664 11104
rect 23716 11092 23722 11144
rect 21542 11064 21548 11076
rect 10796 11036 11008 11064
rect 21330 11036 21548 11064
rect 3513 10999 3571 11005
rect 3513 10996 3525 10999
rect 2675 10968 3525 10996
rect 3513 10965 3525 10968
rect 3559 10996 3571 10999
rect 3694 10996 3700 11008
rect 3559 10968 3700 10996
rect 3559 10965 3571 10968
rect 3513 10959 3571 10965
rect 3694 10956 3700 10968
rect 3752 10956 3758 11008
rect 10980 10996 11008 11036
rect 21542 11024 21548 11036
rect 21600 11024 21606 11076
rect 21910 11024 21916 11076
rect 21968 11064 21974 11076
rect 23842 11064 23848 11076
rect 21968 11036 23848 11064
rect 21968 11024 21974 11036
rect 23842 11024 23848 11036
rect 23900 11024 23906 11076
rect 24872 11064 24900 11163
rect 24964 11144 24992 11172
rect 25317 11169 25329 11172
rect 25363 11169 25375 11203
rect 25317 11163 25375 11169
rect 24946 11092 24952 11144
rect 25004 11092 25010 11144
rect 25590 11064 25596 11076
rect 24872 11036 25596 11064
rect 25590 11024 25596 11036
rect 25648 11024 25654 11076
rect 11238 10996 11244 11008
rect 10980 10968 11244 10996
rect 11238 10956 11244 10968
rect 11296 10996 11302 11008
rect 11882 10996 11888 11008
rect 11296 10968 11888 10996
rect 11296 10956 11302 10968
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 20438 10956 20444 11008
rect 20496 10996 20502 11008
rect 20533 10999 20591 11005
rect 20533 10996 20545 10999
rect 20496 10968 20545 10996
rect 20496 10956 20502 10968
rect 20533 10965 20545 10968
rect 20579 10996 20591 10999
rect 20990 10996 20996 11008
rect 20579 10968 20996 10996
rect 20579 10965 20591 10968
rect 20533 10959 20591 10965
rect 20990 10956 20996 10968
rect 21048 10956 21054 11008
rect 22097 10999 22155 11005
rect 22097 10965 22109 10999
rect 22143 10996 22155 10999
rect 22278 10996 22284 11008
rect 22143 10968 22284 10996
rect 22143 10965 22155 10968
rect 22097 10959 22155 10965
rect 22278 10956 22284 10968
rect 22336 10956 22342 11008
rect 23750 10956 23756 11008
rect 23808 10996 23814 11008
rect 24305 10999 24363 11005
rect 24305 10996 24317 10999
rect 23808 10968 24317 10996
rect 23808 10956 23814 10968
rect 24305 10965 24317 10968
rect 24351 10965 24363 10999
rect 24305 10959 24363 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1673 10795 1731 10801
rect 1673 10761 1685 10795
rect 1719 10792 1731 10795
rect 1762 10792 1768 10804
rect 1719 10764 1768 10792
rect 1719 10761 1731 10764
rect 1673 10755 1731 10761
rect 1762 10752 1768 10764
rect 1820 10752 1826 10804
rect 2590 10752 2596 10804
rect 2648 10792 2654 10804
rect 2866 10792 2872 10804
rect 2648 10764 2872 10792
rect 2648 10752 2654 10764
rect 2866 10752 2872 10764
rect 2924 10792 2930 10804
rect 3237 10795 3295 10801
rect 3237 10792 3249 10795
rect 2924 10764 3249 10792
rect 2924 10752 2930 10764
rect 3237 10761 3249 10764
rect 3283 10761 3295 10795
rect 4798 10792 4804 10804
rect 4759 10764 4804 10792
rect 3237 10755 3295 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 5534 10792 5540 10804
rect 5495 10764 5540 10792
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 6420 10764 6561 10792
rect 6420 10752 6426 10764
rect 6549 10761 6561 10764
rect 6595 10761 6607 10795
rect 7190 10792 7196 10804
rect 7151 10764 7196 10792
rect 6549 10755 6607 10761
rect 7190 10752 7196 10764
rect 7248 10752 7254 10804
rect 7650 10792 7656 10804
rect 7611 10764 7656 10792
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 10870 10792 10876 10804
rect 10831 10764 10876 10792
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11241 10795 11299 10801
rect 11241 10761 11253 10795
rect 11287 10792 11299 10795
rect 11330 10792 11336 10804
rect 11287 10764 11336 10792
rect 11287 10761 11299 10764
rect 11241 10755 11299 10761
rect 11330 10752 11336 10764
rect 11388 10752 11394 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 13541 10795 13599 10801
rect 13541 10792 13553 10795
rect 12860 10764 13553 10792
rect 12860 10752 12866 10764
rect 13541 10761 13553 10764
rect 13587 10792 13599 10795
rect 13722 10792 13728 10804
rect 13587 10764 13728 10792
rect 13587 10761 13599 10764
rect 13541 10755 13599 10761
rect 13722 10752 13728 10764
rect 13780 10792 13786 10804
rect 14093 10795 14151 10801
rect 14093 10792 14105 10795
rect 13780 10764 14105 10792
rect 13780 10752 13786 10764
rect 14093 10761 14105 10764
rect 14139 10761 14151 10795
rect 14093 10755 14151 10761
rect 2314 10724 2320 10736
rect 2275 10696 2320 10724
rect 2314 10684 2320 10696
rect 2372 10684 2378 10736
rect 2406 10656 2412 10668
rect 2240 10628 2412 10656
rect 2240 10597 2268 10628
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 6181 10659 6239 10665
rect 6181 10656 6193 10659
rect 3007 10628 6193 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10557 2283 10591
rect 2498 10588 2504 10600
rect 2459 10560 2504 10588
rect 2225 10551 2283 10557
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 3605 10591 3663 10597
rect 3605 10557 3617 10591
rect 3651 10588 3663 10591
rect 4433 10591 4491 10597
rect 4433 10588 4445 10591
rect 3651 10560 4445 10588
rect 3651 10557 3663 10560
rect 3605 10551 3663 10557
rect 4433 10557 4445 10560
rect 4479 10588 4491 10591
rect 4522 10588 4528 10600
rect 4479 10560 4528 10588
rect 4479 10557 4491 10560
rect 4433 10551 4491 10557
rect 4522 10548 4528 10560
rect 4580 10588 4586 10600
rect 5736 10597 5764 10628
rect 6181 10625 6193 10628
rect 6227 10656 6239 10659
rect 7282 10656 7288 10668
rect 6227 10628 7288 10656
rect 6227 10625 6239 10628
rect 6181 10619 6239 10625
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7834 10656 7840 10668
rect 7795 10628 7840 10656
rect 7834 10616 7840 10628
rect 7892 10656 7898 10668
rect 8757 10659 8815 10665
rect 8757 10656 8769 10659
rect 7892 10628 8769 10656
rect 7892 10616 7898 10628
rect 8757 10625 8769 10628
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 10505 10659 10563 10665
rect 10505 10656 10517 10659
rect 9732 10628 10517 10656
rect 9732 10616 9738 10628
rect 10505 10625 10517 10628
rect 10551 10656 10563 10659
rect 12526 10656 12532 10668
rect 10551 10628 11100 10656
rect 12487 10628 12532 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 5721 10591 5779 10597
rect 4580 10560 4936 10588
rect 4580 10548 4586 10560
rect 2133 10523 2191 10529
rect 2133 10489 2145 10523
rect 2179 10520 2191 10523
rect 2516 10520 2544 10548
rect 2179 10492 2544 10520
rect 2179 10489 2191 10492
rect 2133 10483 2191 10489
rect 4908 10464 4936 10560
rect 5721 10557 5733 10591
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 8478 10548 8484 10600
rect 8536 10588 8542 10600
rect 9306 10588 9312 10600
rect 8536 10560 8581 10588
rect 9267 10560 9312 10588
rect 8536 10548 8542 10560
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 11072 10597 11100 10628
rect 12526 10616 12532 10628
rect 12584 10616 12590 10668
rect 13354 10616 13360 10668
rect 13412 10656 13418 10668
rect 13538 10656 13544 10668
rect 13412 10628 13544 10656
rect 13412 10616 13418 10628
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10588 11115 10591
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 11103 10560 11529 10588
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 7929 10523 7987 10529
rect 7929 10489 7941 10523
rect 7975 10520 7987 10523
rect 8018 10520 8024 10532
rect 7975 10492 8024 10520
rect 7975 10489 7987 10492
rect 7929 10483 7987 10489
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 9217 10523 9275 10529
rect 9217 10489 9229 10523
rect 9263 10520 9275 10523
rect 9398 10520 9404 10532
rect 9263 10492 9404 10520
rect 9263 10489 9275 10492
rect 9217 10483 9275 10489
rect 9398 10480 9404 10492
rect 9456 10520 9462 10532
rect 9630 10523 9688 10529
rect 9630 10520 9642 10523
rect 9456 10492 9642 10520
rect 9456 10480 9462 10492
rect 9630 10489 9642 10492
rect 9676 10489 9688 10523
rect 9630 10483 9688 10489
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 13173 10523 13231 10529
rect 12676 10492 12721 10520
rect 12676 10480 12682 10492
rect 13173 10489 13185 10523
rect 13219 10520 13231 10523
rect 13354 10520 13360 10532
rect 13219 10492 13360 10520
rect 13219 10489 13231 10492
rect 13173 10483 13231 10489
rect 13354 10480 13360 10492
rect 13412 10480 13418 10532
rect 14108 10520 14136 10755
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 15473 10795 15531 10801
rect 15473 10792 15485 10795
rect 15436 10764 15485 10792
rect 15436 10752 15442 10764
rect 15473 10761 15485 10764
rect 15519 10761 15531 10795
rect 15838 10792 15844 10804
rect 15799 10764 15844 10792
rect 15473 10755 15531 10761
rect 15488 10656 15516 10755
rect 15838 10752 15844 10764
rect 15896 10752 15902 10804
rect 17034 10752 17040 10804
rect 17092 10792 17098 10804
rect 17773 10795 17831 10801
rect 17773 10792 17785 10795
rect 17092 10764 17785 10792
rect 17092 10752 17098 10764
rect 17773 10761 17785 10764
rect 17819 10792 17831 10795
rect 18046 10792 18052 10804
rect 17819 10764 18052 10792
rect 17819 10761 17831 10764
rect 17773 10755 17831 10761
rect 18046 10752 18052 10764
rect 18104 10792 18110 10804
rect 18690 10792 18696 10804
rect 18104 10764 18696 10792
rect 18104 10752 18110 10764
rect 18690 10752 18696 10764
rect 18748 10752 18754 10804
rect 21542 10752 21548 10804
rect 21600 10792 21606 10804
rect 21600 10764 21645 10792
rect 21600 10752 21606 10764
rect 25314 10752 25320 10804
rect 25372 10801 25378 10804
rect 25372 10795 25421 10801
rect 25372 10761 25375 10795
rect 25409 10761 25421 10795
rect 25372 10755 25421 10761
rect 25372 10752 25378 10755
rect 17402 10724 17408 10736
rect 17363 10696 17408 10724
rect 17402 10684 17408 10696
rect 17460 10724 17466 10736
rect 17954 10724 17960 10736
rect 17460 10696 17960 10724
rect 17460 10684 17466 10696
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 21560 10724 21588 10752
rect 21821 10727 21879 10733
rect 21821 10724 21833 10727
rect 21560 10696 21833 10724
rect 21821 10693 21833 10696
rect 21867 10693 21879 10727
rect 21821 10687 21879 10693
rect 18322 10656 18328 10668
rect 15488 10628 18328 10656
rect 14277 10591 14335 10597
rect 14277 10557 14289 10591
rect 14323 10588 14335 10591
rect 14366 10588 14372 10600
rect 14323 10560 14372 10588
rect 14323 10557 14335 10560
rect 14277 10551 14335 10557
rect 14366 10548 14372 10560
rect 14424 10588 14430 10600
rect 14424 10560 14964 10588
rect 14424 10548 14430 10560
rect 14598 10523 14656 10529
rect 14598 10520 14610 10523
rect 14108 10492 14610 10520
rect 14598 10489 14610 10492
rect 14644 10489 14656 10523
rect 14936 10520 14964 10560
rect 15838 10548 15844 10600
rect 15896 10588 15902 10600
rect 16500 10597 16528 10628
rect 18322 10616 18328 10628
rect 18380 10656 18386 10668
rect 18380 10628 18552 10656
rect 18380 10616 18386 10628
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15896 10560 16037 10588
rect 15896 10548 15902 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 16485 10591 16543 10597
rect 16485 10557 16497 10591
rect 16531 10557 16543 10591
rect 18046 10588 18052 10600
rect 18007 10560 18052 10588
rect 16485 10551 16543 10557
rect 18046 10548 18052 10560
rect 18104 10548 18110 10600
rect 18524 10597 18552 10628
rect 21174 10616 21180 10668
rect 21232 10656 21238 10668
rect 21358 10656 21364 10668
rect 21232 10628 21364 10656
rect 21232 10616 21238 10628
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 18509 10591 18567 10597
rect 18509 10557 18521 10591
rect 18555 10557 18567 10591
rect 18509 10551 18567 10557
rect 20441 10591 20499 10597
rect 20441 10557 20453 10591
rect 20487 10588 20499 10591
rect 20990 10588 20996 10600
rect 20487 10560 20521 10588
rect 20951 10560 20996 10588
rect 20487 10557 20499 10560
rect 20441 10551 20499 10557
rect 14936 10492 16160 10520
rect 14598 10483 14656 10489
rect 4246 10452 4252 10464
rect 4207 10424 4252 10452
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 5169 10455 5227 10461
rect 5169 10452 5181 10455
rect 4948 10424 5181 10452
rect 4948 10412 4954 10424
rect 5169 10421 5181 10424
rect 5215 10421 5227 10455
rect 5169 10415 5227 10421
rect 5905 10455 5963 10461
rect 5905 10421 5917 10455
rect 5951 10452 5963 10455
rect 6086 10452 6092 10464
rect 5951 10424 6092 10452
rect 5951 10421 5963 10424
rect 5905 10415 5963 10421
rect 6086 10412 6092 10424
rect 6144 10412 6150 10464
rect 10134 10412 10140 10464
rect 10192 10452 10198 10464
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 10192 10424 10241 10452
rect 10192 10412 10198 10424
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 10229 10415 10287 10421
rect 12066 10412 12072 10464
rect 12124 10452 12130 10464
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 12124 10424 12173 10452
rect 12124 10412 12130 10424
rect 12161 10421 12173 10424
rect 12207 10421 12219 10455
rect 15194 10452 15200 10464
rect 15155 10424 15200 10452
rect 12161 10415 12219 10421
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 16132 10461 16160 10492
rect 19426 10480 19432 10532
rect 19484 10520 19490 10532
rect 19705 10523 19763 10529
rect 19705 10520 19717 10523
rect 19484 10492 19717 10520
rect 19484 10480 19490 10492
rect 19705 10489 19717 10492
rect 19751 10520 19763 10523
rect 20456 10520 20484 10551
rect 20990 10548 20996 10560
rect 21048 10548 21054 10600
rect 20622 10520 20628 10532
rect 19751 10492 20628 10520
rect 19751 10489 19763 10492
rect 19705 10483 19763 10489
rect 20622 10480 20628 10492
rect 20680 10480 20686 10532
rect 21174 10520 21180 10532
rect 21135 10492 21180 10520
rect 21174 10480 21180 10492
rect 21232 10480 21238 10532
rect 21836 10520 21864 10687
rect 22278 10588 22284 10600
rect 22239 10560 22284 10588
rect 22278 10548 22284 10560
rect 22336 10548 22342 10600
rect 22465 10591 22523 10597
rect 22465 10557 22477 10591
rect 22511 10557 22523 10591
rect 22465 10551 22523 10557
rect 22480 10520 22508 10551
rect 24486 10548 24492 10600
rect 24544 10588 24550 10600
rect 25292 10591 25350 10597
rect 25292 10588 25304 10591
rect 24544 10560 25304 10588
rect 24544 10548 24550 10560
rect 25292 10557 25304 10560
rect 25338 10588 25350 10591
rect 26053 10591 26111 10597
rect 26053 10588 26065 10591
rect 25338 10560 26065 10588
rect 25338 10557 25350 10560
rect 25292 10551 25350 10557
rect 26053 10557 26065 10560
rect 26099 10557 26111 10591
rect 26053 10551 26111 10557
rect 23198 10520 23204 10532
rect 21836 10492 23204 10520
rect 23198 10480 23204 10492
rect 23256 10480 23262 10532
rect 23750 10520 23756 10532
rect 23711 10492 23756 10520
rect 23750 10480 23756 10492
rect 23808 10480 23814 10532
rect 23845 10523 23903 10529
rect 23845 10489 23857 10523
rect 23891 10489 23903 10523
rect 23845 10483 23903 10489
rect 24397 10523 24455 10529
rect 24397 10489 24409 10523
rect 24443 10489 24455 10523
rect 24397 10483 24455 10489
rect 16117 10455 16175 10461
rect 16117 10421 16129 10455
rect 16163 10421 16175 10455
rect 18138 10452 18144 10464
rect 18099 10424 18144 10452
rect 16117 10415 16175 10421
rect 18138 10412 18144 10424
rect 18196 10412 18202 10464
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 20349 10455 20407 10461
rect 19392 10424 19437 10452
rect 19392 10412 19398 10424
rect 20349 10421 20361 10455
rect 20395 10452 20407 10455
rect 20438 10452 20444 10464
rect 20395 10424 20444 10452
rect 20395 10421 20407 10424
rect 20349 10415 20407 10421
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 22094 10452 22100 10464
rect 22055 10424 22100 10452
rect 22094 10412 22100 10424
rect 22152 10412 22158 10464
rect 22738 10412 22744 10464
rect 22796 10452 22802 10464
rect 23017 10455 23075 10461
rect 23017 10452 23029 10455
rect 22796 10424 23029 10452
rect 22796 10412 22802 10424
rect 23017 10421 23029 10424
rect 23063 10452 23075 10455
rect 23385 10455 23443 10461
rect 23385 10452 23397 10455
rect 23063 10424 23397 10452
rect 23063 10421 23075 10424
rect 23017 10415 23075 10421
rect 23385 10421 23397 10424
rect 23431 10452 23443 10455
rect 23474 10452 23480 10464
rect 23431 10424 23480 10452
rect 23431 10421 23443 10424
rect 23385 10415 23443 10421
rect 23474 10412 23480 10424
rect 23532 10452 23538 10464
rect 23860 10452 23888 10483
rect 23532 10424 23888 10452
rect 23532 10412 23538 10424
rect 24302 10412 24308 10464
rect 24360 10452 24366 10464
rect 24412 10452 24440 10483
rect 24670 10480 24676 10532
rect 24728 10520 24734 10532
rect 24854 10520 24860 10532
rect 24728 10492 24860 10520
rect 24728 10480 24734 10492
rect 24854 10480 24860 10492
rect 24912 10480 24918 10532
rect 24946 10452 24952 10464
rect 24360 10424 24440 10452
rect 24907 10424 24952 10452
rect 24360 10412 24366 10424
rect 24946 10412 24952 10424
rect 25004 10412 25010 10464
rect 25590 10412 25596 10464
rect 25648 10452 25654 10464
rect 25685 10455 25743 10461
rect 25685 10452 25697 10455
rect 25648 10424 25697 10452
rect 25648 10412 25654 10424
rect 25685 10421 25697 10424
rect 25731 10421 25743 10455
rect 25685 10415 25743 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 4614 10208 4620 10260
rect 4672 10208 4678 10260
rect 5258 10248 5264 10260
rect 5219 10220 5264 10248
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 7837 10251 7895 10257
rect 7837 10217 7849 10251
rect 7883 10248 7895 10251
rect 8018 10248 8024 10260
rect 7883 10220 8024 10248
rect 7883 10217 7895 10220
rect 7837 10211 7895 10217
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 11238 10248 11244 10260
rect 11199 10220 11244 10248
rect 11238 10208 11244 10220
rect 11296 10208 11302 10260
rect 12115 10251 12173 10257
rect 12115 10217 12127 10251
rect 12161 10248 12173 10251
rect 12342 10248 12348 10260
rect 12161 10220 12348 10248
rect 12161 10217 12173 10220
rect 12115 10211 12173 10217
rect 12342 10208 12348 10220
rect 12400 10208 12406 10260
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 12529 10251 12587 10257
rect 12529 10248 12541 10251
rect 12492 10220 12541 10248
rect 12492 10208 12498 10220
rect 12529 10217 12541 10220
rect 12575 10248 12587 10251
rect 12618 10248 12624 10260
rect 12575 10220 12624 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 12897 10251 12955 10257
rect 12897 10217 12909 10251
rect 12943 10248 12955 10251
rect 13262 10248 13268 10260
rect 12943 10220 13268 10248
rect 12943 10217 12955 10220
rect 12897 10211 12955 10217
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 14366 10248 14372 10260
rect 14327 10220 14372 10248
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 15013 10251 15071 10257
rect 15013 10248 15025 10251
rect 14884 10220 15025 10248
rect 14884 10208 14890 10220
rect 15013 10217 15025 10220
rect 15059 10217 15071 10251
rect 15013 10211 15071 10217
rect 15194 10208 15200 10260
rect 15252 10248 15258 10260
rect 15654 10248 15660 10260
rect 15252 10220 15660 10248
rect 15252 10208 15258 10220
rect 15654 10208 15660 10220
rect 15712 10248 15718 10260
rect 16301 10251 16359 10257
rect 16301 10248 16313 10251
rect 15712 10220 16313 10248
rect 15712 10208 15718 10220
rect 16301 10217 16313 10220
rect 16347 10217 16359 10251
rect 16301 10211 16359 10217
rect 17221 10251 17279 10257
rect 17221 10217 17233 10251
rect 17267 10248 17279 10251
rect 17310 10248 17316 10260
rect 17267 10220 17316 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 18322 10248 18328 10260
rect 18283 10220 18328 10248
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 21082 10257 21088 10260
rect 21039 10251 21088 10257
rect 21039 10217 21051 10251
rect 21085 10217 21088 10251
rect 21039 10211 21088 10217
rect 21082 10208 21088 10211
rect 21140 10208 21146 10260
rect 21174 10208 21180 10260
rect 21232 10248 21238 10260
rect 21729 10251 21787 10257
rect 21729 10248 21741 10251
rect 21232 10220 21741 10248
rect 21232 10208 21238 10220
rect 21729 10217 21741 10220
rect 21775 10248 21787 10251
rect 21818 10248 21824 10260
rect 21775 10220 21824 10248
rect 21775 10217 21787 10220
rect 21729 10211 21787 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 22833 10251 22891 10257
rect 22833 10217 22845 10251
rect 22879 10217 22891 10251
rect 23382 10248 23388 10260
rect 23343 10220 23388 10248
rect 22833 10211 22891 10217
rect 1762 10140 1768 10192
rect 1820 10180 1826 10192
rect 2225 10183 2283 10189
rect 2225 10180 2237 10183
rect 1820 10152 2237 10180
rect 1820 10140 1826 10152
rect 2225 10149 2237 10152
rect 2271 10149 2283 10183
rect 2225 10143 2283 10149
rect 2590 10140 2596 10192
rect 2648 10180 2654 10192
rect 3145 10183 3203 10189
rect 3145 10180 3157 10183
rect 2648 10152 3157 10180
rect 2648 10140 2654 10152
rect 3145 10149 3157 10152
rect 3191 10149 3203 10183
rect 3145 10143 3203 10149
rect 4341 10183 4399 10189
rect 4341 10149 4353 10183
rect 4387 10180 4399 10183
rect 4632 10180 4660 10208
rect 8757 10183 8815 10189
rect 4387 10152 4660 10180
rect 5092 10152 6684 10180
rect 4387 10149 4399 10152
rect 4341 10143 4399 10149
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 2314 10112 2320 10124
rect 1443 10084 2320 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 2314 10072 2320 10084
rect 2372 10072 2378 10124
rect 2406 10072 2412 10124
rect 2464 10112 2470 10124
rect 2685 10115 2743 10121
rect 2464 10084 2636 10112
rect 2464 10072 2470 10084
rect 2608 10056 2636 10084
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 3513 10115 3571 10121
rect 3513 10112 3525 10115
rect 2731 10084 3525 10112
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 3513 10081 3525 10084
rect 3559 10112 3571 10115
rect 3878 10112 3884 10124
rect 3559 10084 3884 10112
rect 3559 10081 3571 10084
rect 3513 10075 3571 10081
rect 3878 10072 3884 10084
rect 3936 10112 3942 10124
rect 4356 10112 4384 10143
rect 5092 10124 5120 10152
rect 3936 10084 4384 10112
rect 3936 10072 3942 10084
rect 4614 10072 4620 10124
rect 4672 10112 4678 10124
rect 4798 10112 4804 10124
rect 4672 10084 4804 10112
rect 4672 10072 4678 10084
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 5074 10112 5080 10124
rect 5035 10084 5080 10112
rect 5074 10072 5080 10084
rect 5132 10072 5138 10124
rect 6362 10072 6368 10124
rect 6420 10121 6426 10124
rect 6656 10121 6684 10152
rect 8757 10149 8769 10183
rect 8803 10180 8815 10183
rect 9306 10180 9312 10192
rect 8803 10152 9312 10180
rect 8803 10149 8815 10152
rect 8757 10143 8815 10149
rect 9306 10140 9312 10152
rect 9364 10140 9370 10192
rect 10134 10140 10140 10192
rect 10192 10180 10198 10192
rect 10413 10183 10471 10189
rect 10413 10180 10425 10183
rect 10192 10152 10425 10180
rect 10192 10140 10198 10152
rect 10413 10149 10425 10152
rect 10459 10149 10471 10183
rect 10962 10180 10968 10192
rect 10923 10152 10968 10180
rect 10413 10143 10471 10149
rect 10962 10140 10968 10152
rect 11020 10140 11026 10192
rect 13170 10180 13176 10192
rect 13131 10152 13176 10180
rect 13170 10140 13176 10152
rect 13228 10140 13234 10192
rect 17494 10180 17500 10192
rect 17455 10152 17500 10180
rect 17494 10140 17500 10152
rect 17552 10140 17558 10192
rect 22002 10140 22008 10192
rect 22060 10180 22066 10192
rect 22094 10180 22100 10192
rect 22060 10152 22100 10180
rect 22060 10140 22066 10152
rect 22094 10140 22100 10152
rect 22152 10180 22158 10192
rect 22234 10183 22292 10189
rect 22234 10180 22246 10183
rect 22152 10152 22246 10180
rect 22152 10140 22158 10152
rect 22234 10149 22246 10152
rect 22280 10149 22292 10183
rect 22848 10180 22876 10211
rect 23382 10208 23388 10220
rect 23440 10208 23446 10260
rect 24854 10248 24860 10260
rect 23860 10220 24860 10248
rect 23860 10189 23888 10220
rect 24854 10208 24860 10220
rect 24912 10208 24918 10260
rect 23845 10183 23903 10189
rect 23845 10180 23857 10183
rect 22848 10152 23857 10180
rect 22234 10143 22292 10149
rect 23845 10149 23857 10152
rect 23891 10149 23903 10183
rect 23845 10143 23903 10149
rect 24210 10140 24216 10192
rect 24268 10180 24274 10192
rect 24397 10183 24455 10189
rect 24397 10180 24409 10183
rect 24268 10152 24409 10180
rect 24268 10140 24274 10152
rect 24397 10149 24409 10152
rect 24443 10180 24455 10183
rect 24486 10180 24492 10192
rect 24443 10152 24492 10180
rect 24443 10149 24455 10152
rect 24397 10143 24455 10149
rect 24486 10140 24492 10152
rect 24544 10140 24550 10192
rect 6420 10112 6428 10121
rect 6641 10115 6699 10121
rect 6420 10084 6465 10112
rect 6420 10075 6428 10084
rect 6641 10081 6653 10115
rect 6687 10081 6699 10115
rect 6641 10075 6699 10081
rect 6420 10072 6426 10075
rect 7006 10072 7012 10124
rect 7064 10112 7070 10124
rect 8018 10112 8024 10124
rect 7064 10084 8024 10112
rect 7064 10072 7070 10084
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 8481 10115 8539 10121
rect 8481 10112 8493 10115
rect 8444 10084 8493 10112
rect 8444 10072 8450 10084
rect 8481 10081 8493 10084
rect 8527 10081 8539 10115
rect 8481 10075 8539 10081
rect 11790 10072 11796 10124
rect 11848 10112 11854 10124
rect 12012 10115 12070 10121
rect 12012 10112 12024 10115
rect 11848 10084 12024 10112
rect 11848 10072 11854 10084
rect 12012 10081 12024 10084
rect 12058 10112 12070 10115
rect 12710 10112 12716 10124
rect 12058 10084 12716 10112
rect 12058 10081 12070 10084
rect 12012 10075 12070 10081
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 15565 10115 15623 10121
rect 15565 10081 15577 10115
rect 15611 10081 15623 10115
rect 15746 10112 15752 10124
rect 15707 10084 15752 10112
rect 15565 10075 15623 10081
rect 1302 10004 1308 10056
rect 1360 10044 1366 10056
rect 1578 10044 1584 10056
rect 1360 10016 1584 10044
rect 1360 10004 1366 10016
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 1946 10004 1952 10056
rect 2004 10004 2010 10056
rect 2590 10004 2596 10056
rect 2648 10004 2654 10056
rect 6914 10044 6920 10056
rect 6875 10016 6920 10044
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 10042 10004 10048 10056
rect 10100 10044 10106 10056
rect 10321 10047 10379 10053
rect 10321 10044 10333 10047
rect 10100 10016 10333 10044
rect 10100 10004 10106 10016
rect 10321 10013 10333 10016
rect 10367 10013 10379 10047
rect 10321 10007 10379 10013
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10013 13139 10047
rect 13354 10044 13360 10056
rect 13315 10016 13360 10044
rect 13081 10007 13139 10013
rect 1964 9976 1992 10004
rect 2406 9976 2412 9988
rect 1964 9948 2412 9976
rect 2406 9936 2412 9948
rect 2464 9936 2470 9988
rect 2501 9979 2559 9985
rect 2501 9945 2513 9979
rect 2547 9945 2559 9979
rect 2501 9939 2559 9945
rect 4709 9979 4767 9985
rect 4709 9945 4721 9979
rect 4755 9976 4767 9979
rect 4890 9976 4896 9988
rect 4755 9948 4896 9976
rect 4755 9945 4767 9948
rect 4709 9939 4767 9945
rect 1578 9908 1584 9920
rect 1539 9880 1584 9908
rect 1578 9868 1584 9880
rect 1636 9868 1642 9920
rect 1946 9908 1952 9920
rect 1907 9880 1952 9908
rect 1946 9868 1952 9880
rect 2004 9868 2010 9920
rect 2516 9908 2544 9939
rect 4890 9936 4896 9948
rect 4948 9936 4954 9988
rect 6273 9979 6331 9985
rect 6273 9945 6285 9979
rect 6319 9976 6331 9979
rect 6457 9979 6515 9985
rect 6457 9976 6469 9979
rect 6319 9948 6469 9976
rect 6319 9945 6331 9948
rect 6273 9939 6331 9945
rect 6457 9945 6469 9948
rect 6503 9945 6515 9979
rect 13096 9976 13124 10007
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 15580 10044 15608 10075
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 18874 10112 18880 10124
rect 18835 10084 18880 10112
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 19337 10115 19395 10121
rect 19337 10081 19349 10115
rect 19383 10112 19395 10115
rect 20254 10112 20260 10124
rect 19383 10084 20260 10112
rect 19383 10081 19395 10084
rect 19337 10075 19395 10081
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 20968 10115 21026 10121
rect 20968 10081 20980 10115
rect 21014 10112 21026 10115
rect 21450 10112 21456 10124
rect 21014 10084 21456 10112
rect 21014 10081 21026 10084
rect 20968 10075 21026 10081
rect 21450 10072 21456 10084
rect 21508 10112 21514 10124
rect 21634 10112 21640 10124
rect 21508 10084 21640 10112
rect 21508 10072 21514 10084
rect 21634 10072 21640 10084
rect 21692 10072 21698 10124
rect 25222 10112 25228 10124
rect 25183 10084 25228 10112
rect 25222 10072 25228 10084
rect 25280 10072 25286 10124
rect 15654 10044 15660 10056
rect 15580 10016 15660 10044
rect 15654 10004 15660 10016
rect 15712 10004 15718 10056
rect 15838 10044 15844 10056
rect 15799 10016 15844 10044
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 17405 10047 17463 10053
rect 17405 10013 17417 10047
rect 17451 10044 17463 10047
rect 17678 10044 17684 10056
rect 17451 10016 17684 10044
rect 17451 10013 17463 10016
rect 17405 10007 17463 10013
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 18046 10044 18052 10056
rect 18007 10016 18052 10044
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 19426 10044 19432 10056
rect 19387 10016 19432 10044
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 21910 10044 21916 10056
rect 21871 10016 21916 10044
rect 21910 10004 21916 10016
rect 21968 10004 21974 10056
rect 23198 10004 23204 10056
rect 23256 10044 23262 10056
rect 23753 10047 23811 10053
rect 23753 10044 23765 10047
rect 23256 10016 23765 10044
rect 23256 10004 23262 10016
rect 23676 9988 23704 10016
rect 23753 10013 23765 10016
rect 23799 10013 23811 10047
rect 24026 10044 24032 10056
rect 23753 10007 23811 10013
rect 23952 10016 24032 10044
rect 23952 9988 23980 10016
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 13722 9976 13728 9988
rect 13096 9948 13728 9976
rect 6457 9939 6515 9945
rect 3694 9908 3700 9920
rect 2516 9880 3700 9908
rect 3694 9868 3700 9880
rect 3752 9908 3758 9920
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 3752 9880 3893 9908
rect 3752 9868 3758 9880
rect 3881 9877 3893 9880
rect 3927 9908 3939 9911
rect 4246 9908 4252 9920
rect 3927 9880 4252 9908
rect 3927 9877 3939 9880
rect 3881 9871 3939 9877
rect 4246 9868 4252 9880
rect 4304 9908 4310 9920
rect 6288 9908 6316 9939
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 21450 9936 21456 9988
rect 21508 9976 21514 9988
rect 22554 9976 22560 9988
rect 21508 9948 22560 9976
rect 21508 9936 21514 9948
rect 22554 9936 22560 9948
rect 22612 9936 22618 9988
rect 23658 9936 23664 9988
rect 23716 9936 23722 9988
rect 23934 9936 23940 9988
rect 23992 9936 23998 9988
rect 24302 9936 24308 9988
rect 24360 9936 24366 9988
rect 4304 9880 6316 9908
rect 4304 9868 4310 9880
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 16669 9911 16727 9917
rect 16669 9908 16681 9911
rect 16632 9880 16681 9908
rect 16632 9868 16638 9880
rect 16669 9877 16681 9880
rect 16715 9877 16727 9911
rect 16669 9871 16727 9877
rect 19242 9868 19248 9920
rect 19300 9908 19306 9920
rect 19889 9911 19947 9917
rect 19889 9908 19901 9911
rect 19300 9880 19901 9908
rect 19300 9868 19306 9880
rect 19889 9877 19901 9880
rect 19935 9877 19947 9911
rect 19889 9871 19947 9877
rect 20533 9911 20591 9917
rect 20533 9877 20545 9911
rect 20579 9908 20591 9911
rect 20622 9908 20628 9920
rect 20579 9880 20628 9908
rect 20579 9877 20591 9880
rect 20533 9871 20591 9877
rect 20622 9868 20628 9880
rect 20680 9868 20686 9920
rect 20714 9868 20720 9920
rect 20772 9908 20778 9920
rect 21082 9908 21088 9920
rect 20772 9880 21088 9908
rect 20772 9868 20778 9880
rect 21082 9868 21088 9880
rect 21140 9868 21146 9920
rect 23382 9868 23388 9920
rect 23440 9908 23446 9920
rect 23842 9908 23848 9920
rect 23440 9880 23848 9908
rect 23440 9868 23446 9880
rect 23842 9868 23848 9880
rect 23900 9868 23906 9920
rect 24026 9868 24032 9920
rect 24084 9908 24090 9920
rect 24320 9908 24348 9936
rect 25406 9908 25412 9920
rect 24084 9880 24348 9908
rect 25367 9880 25412 9908
rect 24084 9868 24090 9880
rect 25406 9868 25412 9880
rect 25464 9868 25470 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 4338 9704 4344 9716
rect 2556 9676 4344 9704
rect 2556 9664 2562 9676
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 4614 9664 4620 9716
rect 4672 9704 4678 9716
rect 6362 9704 6368 9716
rect 4672 9676 6368 9704
rect 4672 9664 4678 9676
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 8018 9704 8024 9716
rect 7979 9676 8024 9704
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 8386 9704 8392 9716
rect 8347 9676 8392 9704
rect 8386 9664 8392 9676
rect 8444 9664 8450 9716
rect 9677 9707 9735 9713
rect 9677 9673 9689 9707
rect 9723 9704 9735 9707
rect 10045 9707 10103 9713
rect 10045 9704 10057 9707
rect 9723 9676 10057 9704
rect 9723 9673 9735 9676
rect 9677 9667 9735 9673
rect 10045 9673 10057 9676
rect 10091 9704 10103 9707
rect 10134 9704 10140 9716
rect 10091 9676 10140 9704
rect 10091 9673 10103 9676
rect 10045 9667 10103 9673
rect 10134 9664 10140 9676
rect 10192 9664 10198 9716
rect 11790 9664 11796 9716
rect 11848 9704 11854 9716
rect 11977 9707 12035 9713
rect 11977 9704 11989 9707
rect 11848 9676 11989 9704
rect 11848 9664 11854 9676
rect 11977 9673 11989 9676
rect 12023 9673 12035 9707
rect 11977 9667 12035 9673
rect 12897 9707 12955 9713
rect 12897 9673 12909 9707
rect 12943 9704 12955 9707
rect 13170 9704 13176 9716
rect 12943 9676 13176 9704
rect 12943 9673 12955 9676
rect 12897 9667 12955 9673
rect 13170 9664 13176 9676
rect 13228 9664 13234 9716
rect 13998 9664 14004 9716
rect 14056 9704 14062 9716
rect 15746 9704 15752 9716
rect 14056 9676 14504 9704
rect 14056 9664 14062 9676
rect 1762 9645 1768 9648
rect 1746 9639 1768 9645
rect 1746 9605 1758 9639
rect 1746 9599 1768 9605
rect 1762 9596 1768 9599
rect 1820 9596 1826 9648
rect 1857 9639 1915 9645
rect 1857 9605 1869 9639
rect 1903 9636 1915 9639
rect 2222 9636 2228 9648
rect 1903 9608 2084 9636
rect 2183 9608 2228 9636
rect 1903 9605 1915 9608
rect 1857 9599 1915 9605
rect 1946 9568 1952 9580
rect 1907 9540 1952 9568
rect 1946 9528 1952 9540
rect 2004 9528 2010 9580
rect 2056 9568 2084 9608
rect 2222 9596 2228 9608
rect 2280 9596 2286 9648
rect 2958 9636 2964 9648
rect 2919 9608 2964 9636
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 3142 9596 3148 9648
rect 3200 9636 3206 9648
rect 10778 9636 10784 9648
rect 3200 9608 3648 9636
rect 10739 9608 10784 9636
rect 3200 9596 3206 9608
rect 2130 9568 2136 9580
rect 2043 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9568 2194 9580
rect 2593 9571 2651 9577
rect 2593 9568 2605 9571
rect 2188 9540 2605 9568
rect 2188 9528 2194 9540
rect 2593 9537 2605 9540
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 1302 9460 1308 9512
rect 1360 9500 1366 9512
rect 1581 9503 1639 9509
rect 1581 9500 1593 9503
rect 1360 9472 1593 9500
rect 1360 9460 1366 9472
rect 1581 9469 1593 9472
rect 1627 9469 1639 9503
rect 1964 9500 1992 9528
rect 2222 9500 2228 9512
rect 1964 9472 2228 9500
rect 1581 9463 1639 9469
rect 1596 9432 1624 9463
rect 2222 9460 2228 9472
rect 2280 9460 2286 9512
rect 2976 9500 3004 9596
rect 3620 9512 3648 9608
rect 10778 9596 10784 9608
rect 10836 9596 10842 9648
rect 5258 9568 5264 9580
rect 5219 9540 5264 9568
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 10226 9528 10232 9580
rect 10284 9568 10290 9580
rect 11149 9571 11207 9577
rect 11149 9568 11161 9571
rect 10284 9540 11161 9568
rect 10284 9528 10290 9540
rect 11149 9537 11161 9540
rect 11195 9537 11207 9571
rect 13354 9568 13360 9580
rect 13315 9540 13360 9568
rect 11149 9531 11207 9537
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 14274 9528 14280 9580
rect 14332 9568 14338 9580
rect 14476 9568 14504 9676
rect 15120 9676 15752 9704
rect 14921 9639 14979 9645
rect 14921 9605 14933 9639
rect 14967 9636 14979 9639
rect 15120 9636 15148 9676
rect 15746 9664 15752 9676
rect 15804 9704 15810 9716
rect 17405 9707 17463 9713
rect 15804 9676 16620 9704
rect 15804 9664 15810 9676
rect 14967 9608 15148 9636
rect 16592 9636 16620 9676
rect 17405 9673 17417 9707
rect 17451 9704 17463 9707
rect 17494 9704 17500 9716
rect 17451 9676 17500 9704
rect 17451 9673 17463 9676
rect 17405 9667 17463 9673
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 19334 9704 19340 9716
rect 19260 9676 19340 9704
rect 17310 9636 17316 9648
rect 16592 9608 17316 9636
rect 14967 9605 14979 9608
rect 14921 9599 14979 9605
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 18233 9639 18291 9645
rect 18233 9605 18245 9639
rect 18279 9636 18291 9639
rect 19260 9636 19288 9676
rect 19334 9664 19340 9676
rect 19392 9664 19398 9716
rect 20254 9704 20260 9716
rect 20167 9676 20260 9704
rect 20254 9664 20260 9676
rect 20312 9704 20318 9716
rect 20990 9704 20996 9716
rect 20312 9676 20996 9704
rect 20312 9664 20318 9676
rect 20990 9664 20996 9676
rect 21048 9704 21054 9716
rect 22002 9704 22008 9716
rect 21048 9676 22008 9704
rect 21048 9664 21054 9676
rect 22002 9664 22008 9676
rect 22060 9664 22066 9716
rect 22738 9704 22744 9716
rect 22699 9676 22744 9704
rect 22738 9664 22744 9676
rect 22796 9664 22802 9716
rect 24765 9707 24823 9713
rect 24765 9673 24777 9707
rect 24811 9704 24823 9707
rect 24854 9704 24860 9716
rect 24811 9676 24860 9704
rect 24811 9673 24823 9676
rect 24765 9667 24823 9673
rect 24854 9664 24860 9676
rect 24912 9664 24918 9716
rect 25314 9664 25320 9716
rect 25372 9704 25378 9716
rect 26053 9707 26111 9713
rect 26053 9704 26065 9707
rect 25372 9676 26065 9704
rect 25372 9664 25378 9676
rect 26053 9673 26065 9676
rect 26099 9673 26111 9707
rect 26053 9667 26111 9673
rect 18279 9608 19288 9636
rect 18279 9605 18291 9608
rect 18233 9599 18291 9605
rect 19242 9568 19248 9580
rect 14332 9540 14504 9568
rect 19203 9540 19248 9568
rect 14332 9528 14338 9540
rect 19242 9528 19248 9540
rect 19300 9528 19306 9580
rect 21818 9568 21824 9580
rect 21779 9540 21824 9568
rect 21818 9528 21824 9540
rect 21876 9528 21882 9580
rect 23014 9528 23020 9580
rect 23072 9568 23078 9580
rect 23753 9571 23811 9577
rect 23753 9568 23765 9571
rect 23072 9540 23765 9568
rect 23072 9528 23078 9540
rect 23753 9537 23765 9540
rect 23799 9568 23811 9571
rect 24026 9568 24032 9580
rect 23799 9540 24032 9568
rect 23799 9537 23811 9540
rect 23753 9531 23811 9537
rect 24026 9528 24032 9540
rect 24084 9528 24090 9580
rect 24210 9568 24216 9580
rect 24171 9540 24216 9568
rect 24210 9528 24216 9540
rect 24268 9528 24274 9580
rect 3145 9503 3203 9509
rect 3145 9500 3157 9503
rect 2976 9472 3157 9500
rect 3145 9469 3157 9472
rect 3191 9469 3203 9503
rect 3602 9500 3608 9512
rect 3563 9472 3608 9500
rect 3145 9463 3203 9469
rect 3602 9460 3608 9472
rect 3660 9460 3666 9512
rect 4798 9500 4804 9512
rect 4759 9472 4804 9500
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 4890 9460 4896 9512
rect 4948 9500 4954 9512
rect 4948 9472 5041 9500
rect 4948 9460 4954 9472
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5997 9503 6055 9509
rect 5997 9500 6009 9503
rect 5132 9472 6009 9500
rect 5132 9460 5138 9472
rect 5997 9469 6009 9472
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 7098 9500 7104 9512
rect 6696 9472 7104 9500
rect 6696 9460 6702 9472
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9500 7527 9503
rect 7650 9500 7656 9512
rect 7515 9472 7656 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 14826 9460 14832 9512
rect 14884 9500 14890 9512
rect 15013 9503 15071 9509
rect 15013 9500 15025 9503
rect 14884 9472 15025 9500
rect 14884 9460 14890 9472
rect 15013 9469 15025 9472
rect 15059 9500 15071 9503
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 15059 9472 15485 9500
rect 15059 9469 15071 9472
rect 15013 9463 15071 9469
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 15473 9463 15531 9469
rect 17402 9460 17408 9512
rect 17460 9500 17466 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17460 9472 18061 9500
rect 17460 9460 17466 9472
rect 18049 9469 18061 9472
rect 18095 9500 18107 9503
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 18095 9472 18521 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 18509 9469 18521 9472
rect 18555 9500 18567 9503
rect 19058 9500 19064 9512
rect 18555 9472 19064 9500
rect 18555 9469 18567 9472
rect 18509 9463 18567 9469
rect 19058 9460 19064 9472
rect 19116 9460 19122 9512
rect 20784 9503 20842 9509
rect 20784 9469 20796 9503
rect 20830 9500 20842 9503
rect 20830 9472 21036 9500
rect 20830 9469 20842 9472
rect 20784 9463 20842 9469
rect 1946 9432 1952 9444
rect 1596 9404 1952 9432
rect 1946 9392 1952 9404
rect 2004 9392 2010 9444
rect 2866 9392 2872 9444
rect 2924 9432 2930 9444
rect 4614 9432 4620 9444
rect 2924 9404 4620 9432
rect 2924 9392 2930 9404
rect 4614 9392 4620 9404
rect 4672 9392 4678 9444
rect 4908 9432 4936 9460
rect 5258 9432 5264 9444
rect 4908 9404 5264 9432
rect 5258 9392 5264 9404
rect 5316 9392 5322 9444
rect 8665 9435 8723 9441
rect 8665 9401 8677 9435
rect 8711 9401 8723 9435
rect 8665 9395 8723 9401
rect 3142 9324 3148 9376
rect 3200 9364 3206 9376
rect 3237 9367 3295 9373
rect 3237 9364 3249 9367
rect 3200 9336 3249 9364
rect 3200 9324 3206 9336
rect 3237 9333 3249 9336
rect 3283 9333 3295 9367
rect 4338 9364 4344 9376
rect 4299 9336 4344 9364
rect 3237 9327 3295 9333
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 7006 9364 7012 9376
rect 6967 9336 7012 9364
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 8680 9364 8708 9395
rect 8754 9392 8760 9444
rect 8812 9432 8818 9444
rect 9309 9435 9367 9441
rect 8812 9404 8857 9432
rect 8812 9392 8818 9404
rect 9309 9401 9321 9435
rect 9355 9432 9367 9435
rect 9582 9432 9588 9444
rect 9355 9404 9588 9432
rect 9355 9401 9367 9404
rect 9309 9395 9367 9401
rect 9582 9392 9588 9404
rect 9640 9392 9646 9444
rect 10226 9432 10232 9444
rect 10187 9404 10232 9432
rect 10226 9392 10232 9404
rect 10284 9392 10290 9444
rect 10321 9435 10379 9441
rect 10321 9401 10333 9435
rect 10367 9401 10379 9435
rect 10321 9395 10379 9401
rect 13081 9435 13139 9441
rect 13081 9401 13093 9435
rect 13127 9401 13139 9435
rect 13081 9395 13139 9401
rect 9214 9364 9220 9376
rect 8680 9336 9220 9364
rect 9214 9324 9220 9336
rect 9272 9324 9278 9376
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10336 9364 10364 9395
rect 10192 9336 10364 9364
rect 13096 9364 13124 9395
rect 13170 9392 13176 9444
rect 13228 9432 13234 9444
rect 13228 9404 13273 9432
rect 13228 9392 13234 9404
rect 15562 9392 15568 9444
rect 15620 9432 15626 9444
rect 16117 9435 16175 9441
rect 16117 9432 16129 9435
rect 15620 9404 16129 9432
rect 15620 9392 15626 9404
rect 16117 9401 16129 9404
rect 16163 9401 16175 9435
rect 16117 9395 16175 9401
rect 16209 9435 16267 9441
rect 16209 9401 16221 9435
rect 16255 9432 16267 9435
rect 16390 9432 16396 9444
rect 16255 9404 16396 9432
rect 16255 9401 16267 9404
rect 16209 9395 16267 9401
rect 13722 9364 13728 9376
rect 13096 9336 13728 9364
rect 10192 9324 10198 9336
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 14090 9364 14096 9376
rect 13872 9336 14096 9364
rect 13872 9324 13878 9336
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 15197 9367 15255 9373
rect 15197 9333 15209 9367
rect 15243 9364 15255 9367
rect 15378 9364 15384 9376
rect 15243 9336 15384 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 15746 9324 15752 9376
rect 15804 9364 15810 9376
rect 15841 9367 15899 9373
rect 15841 9364 15853 9367
rect 15804 9336 15853 9364
rect 15804 9324 15810 9336
rect 15841 9333 15853 9336
rect 15887 9333 15899 9367
rect 16132 9364 16160 9395
rect 16390 9392 16396 9404
rect 16448 9392 16454 9444
rect 16761 9435 16819 9441
rect 16761 9401 16773 9435
rect 16807 9432 16819 9435
rect 17862 9432 17868 9444
rect 16807 9404 17868 9432
rect 16807 9401 16819 9404
rect 16761 9395 16819 9401
rect 17862 9392 17868 9404
rect 17920 9392 17926 9444
rect 19334 9392 19340 9444
rect 19392 9432 19398 9444
rect 19889 9435 19947 9441
rect 19392 9404 19437 9432
rect 19392 9392 19398 9404
rect 19889 9401 19901 9435
rect 19935 9432 19947 9435
rect 20070 9432 20076 9444
rect 19935 9404 20076 9432
rect 19935 9401 19947 9404
rect 19889 9395 19947 9401
rect 20070 9392 20076 9404
rect 20128 9392 20134 9444
rect 16482 9364 16488 9376
rect 16132 9336 16488 9364
rect 15841 9327 15899 9333
rect 16482 9324 16488 9336
rect 16540 9324 16546 9376
rect 17678 9364 17684 9376
rect 17639 9336 17684 9364
rect 17678 9324 17684 9336
rect 17736 9324 17742 9376
rect 18874 9364 18880 9376
rect 18835 9336 18880 9364
rect 18874 9324 18880 9336
rect 18932 9324 18938 9376
rect 20254 9324 20260 9376
rect 20312 9364 20318 9376
rect 20855 9367 20913 9373
rect 20855 9364 20867 9367
rect 20312 9336 20867 9364
rect 20312 9324 20318 9336
rect 20855 9333 20867 9336
rect 20901 9333 20913 9367
rect 21008 9364 21036 9472
rect 25222 9460 25228 9512
rect 25280 9509 25286 9512
rect 25280 9503 25318 9509
rect 25306 9500 25318 9503
rect 25685 9503 25743 9509
rect 25685 9500 25697 9503
rect 25306 9472 25697 9500
rect 25306 9469 25318 9472
rect 25280 9463 25318 9469
rect 25685 9469 25697 9472
rect 25731 9469 25743 9503
rect 25685 9463 25743 9469
rect 25280 9460 25286 9463
rect 21269 9435 21327 9441
rect 21269 9401 21281 9435
rect 21315 9432 21327 9435
rect 21634 9432 21640 9444
rect 21315 9404 21640 9432
rect 21315 9401 21327 9404
rect 21269 9395 21327 9401
rect 21634 9392 21640 9404
rect 21692 9392 21698 9444
rect 22186 9441 22192 9444
rect 22183 9395 22192 9441
rect 22244 9432 22250 9444
rect 23017 9435 23075 9441
rect 23017 9432 23029 9435
rect 22244 9404 23029 9432
rect 22186 9392 22192 9395
rect 22244 9392 22250 9404
rect 23017 9401 23029 9404
rect 23063 9432 23075 9435
rect 23385 9435 23443 9441
rect 23385 9432 23397 9435
rect 23063 9404 23397 9432
rect 23063 9401 23075 9404
rect 23017 9395 23075 9401
rect 23385 9401 23397 9404
rect 23431 9401 23443 9435
rect 23842 9432 23848 9444
rect 23755 9404 23848 9432
rect 23385 9395 23443 9401
rect 23842 9392 23848 9404
rect 23900 9432 23906 9444
rect 25041 9435 25099 9441
rect 25041 9432 25053 9435
rect 23900 9404 25053 9432
rect 23900 9392 23906 9404
rect 25041 9401 25053 9404
rect 25087 9401 25099 9435
rect 25041 9395 25099 9401
rect 21542 9364 21548 9376
rect 21008 9336 21548 9364
rect 20855 9327 20913 9333
rect 21542 9324 21548 9336
rect 21600 9324 21606 9376
rect 25130 9324 25136 9376
rect 25188 9364 25194 9376
rect 25363 9367 25421 9373
rect 25363 9364 25375 9367
rect 25188 9336 25375 9364
rect 25188 9324 25194 9336
rect 25363 9333 25375 9336
rect 25409 9333 25421 9367
rect 25363 9327 25421 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 2682 9160 2688 9172
rect 1995 9132 2688 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1964 9024 1992 9123
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 4798 9160 4804 9172
rect 3160 9132 4804 9160
rect 2314 9092 2320 9104
rect 2275 9064 2320 9092
rect 2314 9052 2320 9064
rect 2372 9052 2378 9104
rect 3160 9101 3188 9132
rect 4798 9120 4804 9132
rect 4856 9160 4862 9172
rect 5813 9163 5871 9169
rect 5813 9160 5825 9163
rect 4856 9132 5825 9160
rect 4856 9120 4862 9132
rect 5813 9129 5825 9132
rect 5859 9129 5871 9163
rect 5813 9123 5871 9129
rect 10042 9120 10048 9172
rect 10100 9160 10106 9172
rect 10689 9163 10747 9169
rect 10689 9160 10701 9163
rect 10100 9132 10701 9160
rect 10100 9120 10106 9132
rect 10689 9129 10701 9132
rect 10735 9129 10747 9163
rect 10689 9123 10747 9129
rect 11974 9120 11980 9172
rect 12032 9160 12038 9172
rect 16206 9160 16212 9172
rect 12032 9132 16212 9160
rect 12032 9120 12038 9132
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 17862 9160 17868 9172
rect 17696 9132 17868 9160
rect 3145 9095 3203 9101
rect 3145 9061 3157 9095
rect 3191 9061 3203 9095
rect 3878 9092 3884 9104
rect 3839 9064 3884 9092
rect 3145 9055 3203 9061
rect 2866 9024 2872 9036
rect 1443 8996 1992 9024
rect 2827 8996 2872 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 1762 8916 1768 8968
rect 1820 8956 1826 8968
rect 2590 8956 2596 8968
rect 1820 8928 2596 8956
rect 1820 8916 1826 8928
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 3160 8956 3188 9055
rect 3878 9052 3884 9064
rect 3936 9092 3942 9104
rect 7926 9101 7932 9104
rect 4065 9095 4123 9101
rect 4065 9092 4077 9095
rect 3936 9064 4077 9092
rect 3936 9052 3942 9064
rect 4065 9061 4077 9064
rect 4111 9061 4123 9095
rect 7923 9092 7932 9101
rect 7887 9064 7932 9092
rect 4065 9055 4123 9061
rect 7923 9055 7932 9064
rect 7926 9052 7932 9055
rect 7984 9052 7990 9104
rect 9861 9095 9919 9101
rect 9861 9061 9873 9095
rect 9907 9092 9919 9095
rect 10134 9092 10140 9104
rect 9907 9064 10140 9092
rect 9907 9061 9919 9064
rect 9861 9055 9919 9061
rect 10134 9052 10140 9064
rect 10192 9052 10198 9104
rect 12431 9095 12489 9101
rect 12431 9061 12443 9095
rect 12477 9092 12489 9095
rect 12526 9092 12532 9104
rect 12477 9064 12532 9092
rect 12477 9061 12489 9064
rect 12431 9055 12489 9061
rect 12526 9052 12532 9064
rect 12584 9092 12590 9104
rect 12802 9092 12808 9104
rect 12584 9064 12808 9092
rect 12584 9052 12590 9064
rect 12802 9052 12808 9064
rect 12860 9052 12866 9104
rect 13722 9092 13728 9104
rect 13683 9064 13728 9092
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 15565 9095 15623 9101
rect 15565 9061 15577 9095
rect 15611 9092 15623 9095
rect 16114 9092 16120 9104
rect 15611 9064 16120 9092
rect 15611 9061 15623 9064
rect 15565 9055 15623 9061
rect 16114 9052 16120 9064
rect 16172 9052 16178 9104
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 17129 9095 17187 9101
rect 17129 9092 17141 9095
rect 17092 9064 17141 9092
rect 17092 9052 17098 9064
rect 17129 9061 17141 9064
rect 17175 9092 17187 9095
rect 17494 9092 17500 9104
rect 17175 9064 17500 9092
rect 17175 9061 17187 9064
rect 17129 9055 17187 9061
rect 17494 9052 17500 9064
rect 17552 9052 17558 9104
rect 17696 9101 17724 9132
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 22557 9163 22615 9169
rect 22557 9129 22569 9163
rect 22603 9160 22615 9163
rect 23842 9160 23848 9172
rect 22603 9132 23848 9160
rect 22603 9129 22615 9132
rect 22557 9123 22615 9129
rect 23842 9120 23848 9132
rect 23900 9120 23906 9172
rect 18966 9101 18972 9104
rect 17681 9095 17739 9101
rect 17681 9061 17693 9095
rect 17727 9061 17739 9095
rect 18963 9092 18972 9101
rect 18927 9064 18972 9092
rect 17681 9055 17739 9061
rect 18963 9055 18972 9064
rect 18966 9052 18972 9055
rect 19024 9052 19030 9104
rect 20990 9052 20996 9104
rect 21048 9092 21054 9104
rect 21726 9092 21732 9104
rect 21048 9064 21732 9092
rect 21048 9052 21054 9064
rect 21726 9052 21732 9064
rect 21784 9052 21790 9104
rect 21818 9052 21824 9104
rect 21876 9092 21882 9104
rect 21999 9095 22057 9101
rect 21999 9092 22011 9095
rect 21876 9064 22011 9092
rect 21876 9052 21882 9064
rect 21999 9061 22011 9064
rect 22045 9092 22057 9095
rect 22094 9092 22100 9104
rect 22045 9064 22100 9092
rect 22045 9061 22057 9064
rect 21999 9055 22057 9061
rect 22094 9052 22100 9064
rect 22152 9052 22158 9104
rect 22925 9095 22983 9101
rect 22925 9061 22937 9095
rect 22971 9092 22983 9095
rect 23014 9092 23020 9104
rect 22971 9064 23020 9092
rect 22971 9061 22983 9064
rect 22925 9055 22983 9061
rect 23014 9052 23020 9064
rect 23072 9052 23078 9104
rect 23566 9052 23572 9104
rect 23624 9092 23630 9104
rect 24397 9095 24455 9101
rect 24397 9092 24409 9095
rect 23624 9064 24409 9092
rect 23624 9052 23630 9064
rect 24397 9061 24409 9064
rect 24443 9061 24455 9095
rect 24397 9055 24455 9061
rect 24854 9052 24860 9104
rect 24912 9092 24918 9104
rect 25087 9095 25145 9101
rect 25087 9092 25099 9095
rect 24912 9064 25099 9092
rect 24912 9052 24918 9064
rect 25087 9061 25099 9064
rect 25133 9061 25145 9095
rect 25087 9055 25145 9061
rect 4338 9024 4344 9036
rect 4299 8996 4344 9024
rect 4338 8984 4344 8996
rect 4396 9024 4402 9036
rect 5074 9024 5080 9036
rect 4396 8996 5080 9024
rect 4396 8984 4402 8996
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 6086 9024 6092 9036
rect 6047 8996 6092 9024
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 6454 8984 6460 9036
rect 6512 9024 6518 9036
rect 6549 9027 6607 9033
rect 6549 9024 6561 9027
rect 6512 8996 6561 9024
rect 6512 8984 6518 8996
rect 6549 8993 6561 8996
rect 6595 9024 6607 9027
rect 7650 9024 7656 9036
rect 6595 8996 7656 9024
rect 6595 8993 6607 8996
rect 6549 8987 6607 8993
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 14252 9027 14310 9033
rect 14252 8993 14264 9027
rect 14298 9024 14310 9027
rect 14458 9024 14464 9036
rect 14298 8996 14464 9024
rect 14298 8993 14310 8996
rect 14252 8987 14310 8993
rect 14458 8984 14464 8996
rect 14516 8984 14522 9036
rect 17862 8984 17868 9036
rect 17920 9024 17926 9036
rect 18601 9027 18659 9033
rect 18601 9024 18613 9027
rect 17920 8996 18613 9024
rect 17920 8984 17926 8996
rect 18601 8993 18613 8996
rect 18647 9024 18659 9027
rect 19426 9024 19432 9036
rect 18647 8996 19432 9024
rect 18647 8993 18659 8996
rect 18601 8987 18659 8993
rect 19426 8984 19432 8996
rect 19484 8984 19490 9036
rect 23658 9024 23664 9036
rect 23619 8996 23664 9024
rect 23658 8984 23664 8996
rect 23716 8984 23722 9036
rect 23842 9024 23848 9036
rect 23803 8996 23848 9024
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 24995 9027 25053 9033
rect 24995 8993 25007 9027
rect 25041 8993 25053 9027
rect 24995 8987 25053 8993
rect 2740 8928 3188 8956
rect 6733 8959 6791 8965
rect 2740 8916 2746 8928
rect 6733 8925 6745 8959
rect 6779 8956 6791 8959
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 6779 8928 7573 8956
rect 6779 8925 6791 8928
rect 6733 8919 6791 8925
rect 7561 8925 7573 8928
rect 7607 8956 7619 8959
rect 8662 8956 8668 8968
rect 7607 8928 8668 8956
rect 7607 8925 7619 8928
rect 7561 8919 7619 8925
rect 8662 8916 8668 8928
rect 8720 8916 8726 8968
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 9858 8956 9864 8968
rect 9815 8928 9864 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 9858 8916 9864 8928
rect 9916 8916 9922 8968
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 2958 8888 2964 8900
rect 1627 8860 2964 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 2958 8848 2964 8860
rect 3016 8848 3022 8900
rect 8481 8891 8539 8897
rect 8481 8857 8493 8891
rect 8527 8888 8539 8891
rect 8938 8888 8944 8900
rect 8527 8860 8944 8888
rect 8527 8857 8539 8860
rect 8481 8851 8539 8857
rect 8938 8848 8944 8860
rect 8996 8848 9002 8900
rect 9214 8888 9220 8900
rect 9175 8860 9220 8888
rect 9214 8848 9220 8860
rect 9272 8848 9278 8900
rect 9398 8848 9404 8900
rect 9456 8888 9462 8900
rect 10060 8888 10088 8919
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 12069 8959 12127 8965
rect 12069 8956 12081 8959
rect 11296 8928 12081 8956
rect 11296 8916 11302 8928
rect 12069 8925 12081 8928
rect 12115 8925 12127 8959
rect 12069 8919 12127 8925
rect 15473 8959 15531 8965
rect 15473 8925 15485 8959
rect 15519 8925 15531 8959
rect 15473 8919 15531 8925
rect 16117 8959 16175 8965
rect 16117 8925 16129 8959
rect 16163 8956 16175 8959
rect 16206 8956 16212 8968
rect 16163 8928 16212 8956
rect 16163 8925 16175 8928
rect 16117 8919 16175 8925
rect 9456 8860 10088 8888
rect 12989 8891 13047 8897
rect 9456 8848 9462 8860
rect 12989 8857 13001 8891
rect 13035 8888 13047 8891
rect 13170 8888 13176 8900
rect 13035 8860 13176 8888
rect 13035 8857 13047 8860
rect 12989 8851 13047 8857
rect 13170 8848 13176 8860
rect 13228 8888 13234 8900
rect 13357 8891 13415 8897
rect 13357 8888 13369 8891
rect 13228 8860 13369 8888
rect 13228 8848 13234 8860
rect 13357 8857 13369 8860
rect 13403 8888 13415 8891
rect 13722 8888 13728 8900
rect 13403 8860 13728 8888
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 13722 8848 13728 8860
rect 13780 8848 13786 8900
rect 14323 8891 14381 8897
rect 14323 8857 14335 8891
rect 14369 8888 14381 8891
rect 15013 8891 15071 8897
rect 15013 8888 15025 8891
rect 14369 8860 15025 8888
rect 14369 8857 14381 8860
rect 14323 8851 14381 8857
rect 15013 8857 15025 8860
rect 15059 8888 15071 8891
rect 15488 8888 15516 8919
rect 16206 8916 16212 8928
rect 16264 8916 16270 8968
rect 16574 8916 16580 8968
rect 16632 8956 16638 8968
rect 17037 8959 17095 8965
rect 17037 8956 17049 8959
rect 16632 8928 17049 8956
rect 16632 8916 16638 8928
rect 17037 8925 17049 8928
rect 17083 8925 17095 8959
rect 17037 8919 17095 8925
rect 21637 8959 21695 8965
rect 21637 8925 21649 8959
rect 21683 8956 21695 8959
rect 21726 8956 21732 8968
rect 21683 8928 21732 8956
rect 21683 8925 21695 8928
rect 21637 8919 21695 8925
rect 21726 8916 21732 8928
rect 21784 8916 21790 8968
rect 23937 8959 23995 8965
rect 23937 8925 23949 8959
rect 23983 8925 23995 8959
rect 23937 8919 23995 8925
rect 15059 8860 15516 8888
rect 15059 8857 15071 8860
rect 15013 8851 15071 8857
rect 19150 8848 19156 8900
rect 19208 8888 19214 8900
rect 19426 8888 19432 8900
rect 19208 8860 19432 8888
rect 19208 8848 19214 8860
rect 19426 8848 19432 8860
rect 19484 8848 19490 8900
rect 21545 8891 21603 8897
rect 21545 8857 21557 8891
rect 21591 8888 21603 8891
rect 21910 8888 21916 8900
rect 21591 8860 21916 8888
rect 21591 8857 21603 8860
rect 21545 8851 21603 8857
rect 21910 8848 21916 8860
rect 21968 8888 21974 8900
rect 23952 8888 23980 8919
rect 25015 8900 25043 8987
rect 25015 8888 25044 8900
rect 21968 8860 23980 8888
rect 24951 8860 25044 8888
rect 21968 8848 21974 8860
rect 25038 8848 25044 8860
rect 25096 8888 25102 8900
rect 25222 8888 25228 8900
rect 25096 8860 25228 8888
rect 25096 8848 25102 8860
rect 25222 8848 25228 8860
rect 25280 8848 25286 8900
rect 3513 8823 3571 8829
rect 3513 8789 3525 8823
rect 3559 8820 3571 8823
rect 3602 8820 3608 8832
rect 3559 8792 3608 8820
rect 3559 8789 3571 8792
rect 3513 8783 3571 8789
rect 3602 8780 3608 8792
rect 3660 8820 3666 8832
rect 3878 8820 3884 8832
rect 3660 8792 3884 8820
rect 3660 8780 3666 8792
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 5258 8780 5264 8832
rect 5316 8820 5322 8832
rect 5445 8823 5503 8829
rect 5445 8820 5457 8823
rect 5316 8792 5457 8820
rect 5316 8780 5322 8792
rect 5445 8789 5457 8792
rect 5491 8789 5503 8823
rect 7098 8820 7104 8832
rect 7059 8792 7104 8820
rect 5445 8783 5503 8789
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 7469 8823 7527 8829
rect 7469 8789 7481 8823
rect 7515 8820 7527 8823
rect 7650 8820 7656 8832
rect 7515 8792 7656 8820
rect 7515 8789 7527 8792
rect 7469 8783 7527 8789
rect 7650 8780 7656 8792
rect 7708 8820 7714 8832
rect 8202 8820 8208 8832
rect 7708 8792 8208 8820
rect 7708 8780 7714 8792
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 8754 8820 8760 8832
rect 8628 8792 8760 8820
rect 8628 8780 8634 8792
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 14826 8820 14832 8832
rect 9824 8792 14832 8820
rect 9824 8780 9830 8792
rect 14826 8780 14832 8792
rect 14884 8780 14890 8832
rect 16114 8780 16120 8832
rect 16172 8820 16178 8832
rect 16390 8820 16396 8832
rect 16172 8792 16396 8820
rect 16172 8780 16178 8792
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 19334 8780 19340 8832
rect 19392 8820 19398 8832
rect 19521 8823 19579 8829
rect 19521 8820 19533 8823
rect 19392 8792 19533 8820
rect 19392 8780 19398 8792
rect 19521 8789 19533 8792
rect 19567 8820 19579 8823
rect 19797 8823 19855 8829
rect 19797 8820 19809 8823
rect 19567 8792 19809 8820
rect 19567 8789 19579 8792
rect 19521 8783 19579 8789
rect 19797 8789 19809 8792
rect 19843 8789 19855 8823
rect 21174 8820 21180 8832
rect 21135 8792 21180 8820
rect 19797 8783 19855 8789
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 23198 8820 23204 8832
rect 23159 8792 23204 8820
rect 23198 8780 23204 8792
rect 23256 8780 23262 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 4706 8576 4712 8628
rect 4764 8616 4770 8628
rect 4801 8619 4859 8625
rect 4801 8616 4813 8619
rect 4764 8588 4813 8616
rect 4764 8576 4770 8588
rect 4801 8585 4813 8588
rect 4847 8585 4859 8619
rect 6086 8616 6092 8628
rect 6047 8588 6092 8616
rect 4801 8579 4859 8585
rect 1302 8508 1308 8560
rect 1360 8548 1366 8560
rect 3050 8548 3056 8560
rect 1360 8520 3056 8548
rect 1360 8508 1366 8520
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8480 2743 8483
rect 2958 8480 2964 8492
rect 2731 8452 2964 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 1762 8412 1768 8424
rect 1723 8384 1768 8412
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 3142 8412 3148 8424
rect 3103 8384 3148 8412
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 4816 8412 4844 8579
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 6454 8616 6460 8628
rect 6415 8588 6460 8616
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 7006 8616 7012 8628
rect 6967 8588 7012 8616
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 8481 8619 8539 8625
rect 8481 8585 8493 8619
rect 8527 8616 8539 8619
rect 8570 8616 8576 8628
rect 8527 8588 8576 8616
rect 8527 8585 8539 8588
rect 8481 8579 8539 8585
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 8662 8576 8668 8628
rect 8720 8616 8726 8628
rect 8757 8619 8815 8625
rect 8757 8616 8769 8619
rect 8720 8588 8769 8616
rect 8720 8576 8726 8588
rect 8757 8585 8769 8588
rect 8803 8585 8815 8619
rect 8757 8579 8815 8585
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 9125 8619 9183 8625
rect 9125 8616 9137 8619
rect 8996 8588 9137 8616
rect 8996 8576 9002 8588
rect 9125 8585 9137 8588
rect 9171 8616 9183 8619
rect 9490 8616 9496 8628
rect 9171 8588 9496 8616
rect 9171 8585 9183 8588
rect 9125 8579 9183 8585
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 11698 8576 11704 8628
rect 11756 8616 11762 8628
rect 11793 8619 11851 8625
rect 11793 8616 11805 8619
rect 11756 8588 11805 8616
rect 11756 8576 11762 8588
rect 11793 8585 11805 8588
rect 11839 8585 11851 8619
rect 11793 8579 11851 8585
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 13357 8619 13415 8625
rect 13357 8616 13369 8619
rect 13320 8588 13369 8616
rect 13320 8576 13326 8588
rect 13357 8585 13369 8588
rect 13403 8585 13415 8619
rect 13357 8579 13415 8585
rect 14277 8619 14335 8625
rect 14277 8585 14289 8619
rect 14323 8616 14335 8619
rect 14458 8616 14464 8628
rect 14323 8588 14464 8616
rect 14323 8585 14335 8588
rect 14277 8579 14335 8585
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 14599 8619 14657 8625
rect 14599 8585 14611 8619
rect 14645 8616 14657 8619
rect 15562 8616 15568 8628
rect 14645 8588 15568 8616
rect 14645 8585 14657 8588
rect 14599 8579 14657 8585
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 17034 8616 17040 8628
rect 16995 8588 17040 8616
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 17862 8616 17868 8628
rect 17823 8588 17868 8616
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18279 8619 18337 8625
rect 18279 8585 18291 8619
rect 18325 8616 18337 8619
rect 19242 8616 19248 8628
rect 18325 8588 19248 8616
rect 18325 8585 18337 8588
rect 18279 8579 18337 8585
rect 19242 8576 19248 8588
rect 19300 8576 19306 8628
rect 20254 8616 20260 8628
rect 20215 8588 20260 8616
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 20714 8576 20720 8628
rect 20772 8616 20778 8628
rect 20855 8619 20913 8625
rect 20855 8616 20867 8619
rect 20772 8588 20867 8616
rect 20772 8576 20778 8588
rect 20855 8585 20867 8588
rect 20901 8585 20913 8619
rect 20855 8579 20913 8585
rect 22094 8576 22100 8628
rect 22152 8616 22158 8628
rect 22830 8616 22836 8628
rect 22152 8588 22836 8616
rect 22152 8576 22158 8588
rect 22830 8576 22836 8588
rect 22888 8616 22894 8628
rect 23017 8619 23075 8625
rect 23017 8616 23029 8619
rect 22888 8588 23029 8616
rect 22888 8576 22894 8588
rect 23017 8585 23029 8588
rect 23063 8616 23075 8619
rect 23842 8616 23848 8628
rect 23063 8588 23848 8616
rect 23063 8585 23075 8588
rect 23017 8579 23075 8585
rect 23842 8576 23848 8588
rect 23900 8576 23906 8628
rect 24854 8576 24860 8628
rect 24912 8616 24918 8628
rect 25363 8619 25421 8625
rect 25363 8616 25375 8619
rect 24912 8588 25375 8616
rect 24912 8576 24918 8588
rect 25363 8585 25375 8588
rect 25409 8585 25421 8619
rect 25363 8579 25421 8585
rect 5534 8480 5540 8492
rect 5495 8452 5540 8480
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 7024 8480 7052 8576
rect 11471 8551 11529 8557
rect 11471 8517 11483 8551
rect 11517 8548 11529 8551
rect 12158 8548 12164 8560
rect 11517 8520 12164 8548
rect 11517 8517 11529 8520
rect 11471 8511 11529 8517
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 14366 8508 14372 8560
rect 14424 8548 14430 8560
rect 18049 8551 18107 8557
rect 18049 8548 18061 8551
rect 14424 8520 18061 8548
rect 14424 8508 14430 8520
rect 18049 8517 18061 8520
rect 18095 8548 18107 8551
rect 18601 8551 18659 8557
rect 18601 8548 18613 8551
rect 18095 8520 18613 8548
rect 18095 8517 18107 8520
rect 18049 8511 18107 8517
rect 18601 8517 18613 8520
rect 18647 8517 18659 8551
rect 19794 8548 19800 8560
rect 19755 8520 19800 8548
rect 18601 8511 18659 8517
rect 19794 8508 19800 8520
rect 19852 8508 19858 8560
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 7024 8452 7573 8480
rect 7561 8449 7573 8452
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 9582 8440 9588 8492
rect 9640 8480 9646 8492
rect 9677 8483 9735 8489
rect 9677 8480 9689 8483
rect 9640 8452 9689 8480
rect 9640 8440 9646 8452
rect 9677 8449 9689 8452
rect 9723 8449 9735 8483
rect 9677 8443 9735 8449
rect 15194 8440 15200 8492
rect 15252 8480 15258 8492
rect 15473 8483 15531 8489
rect 15473 8480 15485 8483
rect 15252 8452 15485 8480
rect 15252 8440 15258 8452
rect 15473 8449 15485 8452
rect 15519 8480 15531 8483
rect 15838 8480 15844 8492
rect 15519 8452 15844 8480
rect 15519 8449 15531 8452
rect 15473 8443 15531 8449
rect 15838 8440 15844 8452
rect 15896 8440 15902 8492
rect 17954 8480 17960 8492
rect 16776 8452 17960 8480
rect 16776 8424 16804 8452
rect 17954 8440 17960 8452
rect 18012 8480 18018 8492
rect 18966 8480 18972 8492
rect 18012 8452 18972 8480
rect 18012 8440 18018 8452
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8480 19303 8483
rect 20272 8480 20300 8576
rect 23477 8551 23535 8557
rect 23477 8517 23489 8551
rect 23523 8548 23535 8551
rect 23658 8548 23664 8560
rect 23523 8520 23664 8548
rect 23523 8517 23535 8520
rect 23477 8511 23535 8517
rect 23658 8508 23664 8520
rect 23716 8548 23722 8560
rect 24762 8548 24768 8560
rect 23716 8520 24768 8548
rect 23716 8508 23722 8520
rect 24762 8508 24768 8520
rect 24820 8508 24826 8560
rect 19291 8452 20300 8480
rect 19291 8449 19303 8452
rect 19245 8443 19303 8449
rect 21174 8440 21180 8492
rect 21232 8480 21238 8492
rect 21818 8480 21824 8492
rect 21232 8452 21824 8480
rect 21232 8440 21238 8452
rect 21818 8440 21824 8452
rect 21876 8440 21882 8492
rect 23566 8440 23572 8492
rect 23624 8480 23630 8492
rect 23753 8483 23811 8489
rect 23753 8480 23765 8483
rect 23624 8452 23765 8480
rect 23624 8440 23630 8452
rect 23753 8449 23765 8452
rect 23799 8449 23811 8483
rect 24210 8480 24216 8492
rect 24171 8452 24216 8480
rect 23753 8443 23811 8449
rect 24210 8440 24216 8452
rect 24268 8440 24274 8492
rect 4985 8415 5043 8421
rect 4985 8412 4997 8415
rect 4816 8384 4997 8412
rect 4985 8381 4997 8384
rect 5031 8381 5043 8415
rect 4985 8375 5043 8381
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8381 5503 8415
rect 5445 8375 5503 8381
rect 11400 8415 11458 8421
rect 11400 8381 11412 8415
rect 11446 8412 11458 8415
rect 11698 8412 11704 8424
rect 11446 8384 11704 8412
rect 11446 8381 11458 8384
rect 11400 8375 11458 8381
rect 1486 8304 1492 8356
rect 1544 8344 1550 8356
rect 1581 8347 1639 8353
rect 1581 8344 1593 8347
rect 1544 8316 1593 8344
rect 1544 8304 1550 8316
rect 1581 8313 1593 8316
rect 1627 8313 1639 8347
rect 1581 8307 1639 8313
rect 3466 8347 3524 8353
rect 3466 8313 3478 8347
rect 3512 8313 3524 8347
rect 3466 8307 3524 8313
rect 3053 8279 3111 8285
rect 3053 8245 3065 8279
rect 3099 8276 3111 8279
rect 3142 8276 3148 8288
rect 3099 8248 3148 8276
rect 3099 8245 3111 8248
rect 3053 8239 3111 8245
rect 3142 8236 3148 8248
rect 3200 8276 3206 8288
rect 3481 8276 3509 8307
rect 3200 8248 3509 8276
rect 4065 8279 4123 8285
rect 3200 8236 3206 8248
rect 4065 8245 4077 8279
rect 4111 8276 4123 8279
rect 4246 8276 4252 8288
rect 4111 8248 4252 8276
rect 4111 8245 4123 8248
rect 4065 8239 4123 8245
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 4338 8236 4344 8288
rect 4396 8276 4402 8288
rect 4396 8248 4441 8276
rect 4396 8236 4402 8248
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 5460 8276 5488 8375
rect 11698 8372 11704 8384
rect 11756 8372 11762 8424
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 12986 8412 12992 8424
rect 12483 8384 12992 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 12986 8372 12992 8384
rect 13044 8372 13050 8424
rect 13906 8372 13912 8424
rect 13964 8412 13970 8424
rect 14496 8415 14554 8421
rect 14496 8412 14508 8415
rect 13964 8384 14508 8412
rect 13964 8372 13970 8384
rect 14496 8381 14508 8384
rect 14542 8412 14554 8415
rect 14921 8415 14979 8421
rect 14921 8412 14933 8415
rect 14542 8384 14933 8412
rect 14542 8381 14554 8384
rect 14496 8375 14554 8381
rect 14921 8381 14933 8384
rect 14967 8381 14979 8415
rect 14921 8375 14979 8381
rect 15381 8415 15439 8421
rect 15381 8381 15393 8415
rect 15427 8412 15439 8415
rect 16758 8412 16764 8424
rect 15427 8384 16764 8412
rect 15427 8381 15439 8384
rect 15381 8375 15439 8381
rect 7926 8353 7932 8356
rect 7469 8347 7527 8353
rect 7469 8313 7481 8347
rect 7515 8344 7527 8347
rect 7923 8344 7932 8353
rect 7515 8316 7932 8344
rect 7515 8313 7527 8316
rect 7469 8307 7527 8313
rect 7923 8307 7932 8316
rect 7926 8304 7932 8307
rect 7984 8304 7990 8356
rect 9398 8344 9404 8356
rect 9359 8316 9404 8344
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 9548 8316 9593 8344
rect 9548 8304 9554 8316
rect 9858 8304 9864 8356
rect 9916 8344 9922 8356
rect 10689 8347 10747 8353
rect 10689 8344 10701 8347
rect 9916 8316 10701 8344
rect 9916 8304 9922 8316
rect 10689 8313 10701 8316
rect 10735 8313 10747 8347
rect 11238 8344 11244 8356
rect 11199 8316 11244 8344
rect 10689 8307 10747 8313
rect 11238 8304 11244 8316
rect 11296 8304 11302 8356
rect 12526 8344 12532 8356
rect 12176 8316 12532 8344
rect 5224 8248 5488 8276
rect 5224 8236 5230 8248
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 10321 8279 10379 8285
rect 10321 8276 10333 8279
rect 10192 8248 10333 8276
rect 10192 8236 10198 8248
rect 10321 8245 10333 8248
rect 10367 8245 10379 8279
rect 10321 8239 10379 8245
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 12176 8285 12204 8316
rect 12526 8304 12532 8316
rect 12584 8344 12590 8356
rect 12758 8347 12816 8353
rect 12758 8344 12770 8347
rect 12584 8316 12770 8344
rect 12584 8304 12590 8316
rect 12758 8313 12770 8316
rect 12804 8313 12816 8347
rect 13630 8344 13636 8356
rect 13591 8316 13636 8344
rect 12758 8307 12816 8313
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 15850 8353 15878 8384
rect 16758 8372 16764 8384
rect 16816 8372 16822 8424
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8412 18107 8415
rect 18176 8415 18234 8421
rect 18176 8412 18188 8415
rect 18095 8384 18188 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18176 8381 18188 8384
rect 18222 8381 18234 8415
rect 18176 8375 18234 8381
rect 20714 8372 20720 8424
rect 20772 8421 20778 8424
rect 20772 8415 20810 8421
rect 20798 8412 20810 8415
rect 21269 8415 21327 8421
rect 21269 8412 21281 8415
rect 20798 8384 21281 8412
rect 20798 8381 20810 8384
rect 20772 8375 20810 8381
rect 21269 8381 21281 8384
rect 21315 8381 21327 8415
rect 21269 8375 21327 8381
rect 22741 8415 22799 8421
rect 22741 8381 22753 8415
rect 22787 8381 22799 8415
rect 22741 8375 22799 8381
rect 20772 8372 20778 8375
rect 15835 8347 15893 8353
rect 15835 8313 15847 8347
rect 15881 8344 15893 8347
rect 15881 8316 15915 8344
rect 15881 8313 15893 8316
rect 15835 8307 15893 8313
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 17313 8347 17371 8353
rect 17313 8344 17325 8347
rect 16632 8316 17325 8344
rect 16632 8304 16638 8316
rect 17313 8313 17325 8316
rect 17359 8313 17371 8347
rect 17313 8307 17371 8313
rect 19334 8304 19340 8356
rect 19392 8344 19398 8356
rect 22142 8347 22200 8353
rect 22142 8344 22154 8347
rect 19392 8316 19437 8344
rect 21928 8316 22154 8344
rect 19392 8304 19398 8316
rect 21928 8288 21956 8316
rect 22142 8313 22154 8316
rect 22188 8313 22200 8347
rect 22756 8344 22784 8375
rect 25038 8372 25044 8424
rect 25096 8412 25102 8424
rect 25260 8415 25318 8421
rect 25260 8412 25272 8415
rect 25096 8384 25272 8412
rect 25096 8372 25102 8384
rect 25260 8381 25272 8384
rect 25306 8412 25318 8415
rect 25682 8412 25688 8424
rect 25306 8384 25688 8412
rect 25306 8381 25318 8384
rect 25260 8375 25318 8381
rect 25682 8372 25688 8384
rect 25740 8372 25746 8424
rect 22756 8316 23520 8344
rect 22142 8307 22200 8313
rect 12161 8279 12219 8285
rect 12161 8276 12173 8279
rect 11756 8248 12173 8276
rect 11756 8236 11762 8248
rect 12161 8245 12173 8248
rect 12207 8245 12219 8279
rect 12161 8239 12219 8245
rect 16114 8236 16120 8288
rect 16172 8276 16178 8288
rect 16393 8279 16451 8285
rect 16393 8276 16405 8279
rect 16172 8248 16405 8276
rect 16172 8236 16178 8248
rect 16393 8245 16405 8248
rect 16439 8245 16451 8279
rect 16393 8239 16451 8245
rect 21729 8279 21787 8285
rect 21729 8245 21741 8279
rect 21775 8276 21787 8279
rect 21910 8276 21916 8288
rect 21775 8248 21916 8276
rect 21775 8245 21787 8248
rect 21729 8239 21787 8245
rect 21910 8236 21916 8248
rect 21968 8236 21974 8288
rect 23492 8276 23520 8316
rect 23842 8304 23848 8356
rect 23900 8344 23906 8356
rect 23900 8316 23945 8344
rect 23900 8304 23906 8316
rect 23658 8276 23664 8288
rect 23492 8248 23664 8276
rect 23658 8236 23664 8248
rect 23716 8236 23722 8288
rect 25041 8279 25099 8285
rect 25041 8245 25053 8279
rect 25087 8276 25099 8279
rect 25222 8276 25228 8288
rect 25087 8248 25228 8276
rect 25087 8245 25099 8248
rect 25041 8239 25099 8245
rect 25222 8236 25228 8248
rect 25280 8276 25286 8288
rect 26142 8276 26148 8288
rect 25280 8248 26148 8276
rect 25280 8236 25286 8248
rect 26142 8236 26148 8248
rect 26200 8236 26206 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2041 8075 2099 8081
rect 2041 8041 2053 8075
rect 2087 8072 2099 8075
rect 2682 8072 2688 8084
rect 2087 8044 2688 8072
rect 2087 8041 2099 8044
rect 2041 8035 2099 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 3237 8075 3295 8081
rect 3237 8041 3249 8075
rect 3283 8072 3295 8075
rect 3694 8072 3700 8084
rect 3283 8044 3700 8072
rect 3283 8041 3295 8044
rect 3237 8035 3295 8041
rect 3694 8032 3700 8044
rect 3752 8032 3758 8084
rect 4706 8072 4712 8084
rect 4147 8044 4712 8072
rect 2314 8004 2320 8016
rect 2275 7976 2320 8004
rect 2314 7964 2320 7976
rect 2372 7964 2378 8016
rect 3510 7964 3516 8016
rect 3568 8004 3574 8016
rect 4147 8004 4175 8044
rect 4706 8032 4712 8044
rect 4764 8072 4770 8084
rect 5166 8072 5172 8084
rect 4764 8044 5172 8072
rect 4764 8032 4770 8044
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 5810 8072 5816 8084
rect 5771 8044 5816 8072
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 7653 8075 7711 8081
rect 7653 8041 7665 8075
rect 7699 8072 7711 8075
rect 7742 8072 7748 8084
rect 7699 8044 7748 8072
rect 7699 8041 7711 8044
rect 7653 8035 7711 8041
rect 7742 8032 7748 8044
rect 7800 8072 7806 8084
rect 7926 8072 7932 8084
rect 7800 8044 7932 8072
rect 7800 8032 7806 8044
rect 7926 8032 7932 8044
rect 7984 8072 7990 8084
rect 12342 8072 12348 8084
rect 7984 8044 10082 8072
rect 12303 8044 12348 8072
rect 7984 8032 7990 8044
rect 4246 8004 4252 8016
rect 3568 7976 4175 8004
rect 4207 7976 4252 8004
rect 3568 7964 3574 7976
rect 4246 7964 4252 7976
rect 4304 7964 4310 8016
rect 6270 7964 6276 8016
rect 6328 8004 6334 8016
rect 6641 8007 6699 8013
rect 6641 8004 6653 8007
rect 6328 7976 6653 8004
rect 6328 7964 6334 7976
rect 6641 7973 6653 7976
rect 6687 7973 6699 8007
rect 8754 8004 8760 8016
rect 8715 7976 8760 8004
rect 6641 7967 6699 7973
rect 8754 7964 8760 7976
rect 8812 7964 8818 8016
rect 10054 8013 10082 8044
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 12986 8072 12992 8084
rect 12947 8044 12992 8072
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 15102 8072 15108 8084
rect 13320 8044 13860 8072
rect 15063 8044 15108 8072
rect 13320 8032 13326 8044
rect 10039 8007 10097 8013
rect 10039 7973 10051 8007
rect 10085 8004 10097 8007
rect 11698 8004 11704 8016
rect 10085 7976 11704 8004
rect 10085 7973 10097 7976
rect 10039 7967 10097 7973
rect 11698 7964 11704 7976
rect 11756 8013 11762 8016
rect 11756 8007 11804 8013
rect 11756 7973 11758 8007
rect 11792 7973 11804 8007
rect 11756 7967 11804 7973
rect 13541 8007 13599 8013
rect 13541 7973 13553 8007
rect 13587 8004 13599 8007
rect 13722 8004 13728 8016
rect 13587 7976 13728 8004
rect 13587 7973 13599 7976
rect 13541 7967 13599 7973
rect 11756 7964 11762 7967
rect 13722 7964 13728 7976
rect 13780 7964 13786 8016
rect 13832 8013 13860 8044
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 16114 8072 16120 8084
rect 16075 8044 16120 8072
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 17034 8032 17040 8084
rect 17092 8072 17098 8084
rect 17497 8075 17555 8081
rect 17497 8072 17509 8075
rect 17092 8044 17509 8072
rect 17092 8032 17098 8044
rect 17497 8041 17509 8044
rect 17543 8041 17555 8075
rect 17497 8035 17555 8041
rect 18417 8075 18475 8081
rect 18417 8041 18429 8075
rect 18463 8041 18475 8075
rect 19334 8072 19340 8084
rect 19295 8044 19340 8072
rect 18417 8035 18475 8041
rect 13817 8007 13875 8013
rect 13817 7973 13829 8007
rect 13863 7973 13875 8007
rect 13817 7967 13875 7973
rect 15703 8007 15761 8013
rect 15703 7973 15715 8007
rect 15749 8004 15761 8007
rect 16482 8004 16488 8016
rect 15749 7976 16488 8004
rect 15749 7973 15761 7976
rect 15703 7967 15761 7973
rect 16482 7964 16488 7976
rect 16540 7964 16546 8016
rect 16758 7964 16764 8016
rect 16816 8004 16822 8016
rect 16898 8007 16956 8013
rect 16898 8004 16910 8007
rect 16816 7976 16910 8004
rect 16816 7964 16822 7976
rect 16898 7973 16910 7976
rect 16944 7973 16956 8007
rect 18432 8004 18460 8035
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 22741 8075 22799 8081
rect 22741 8041 22753 8075
rect 22787 8072 22799 8075
rect 23477 8075 23535 8081
rect 23477 8072 23489 8075
rect 22787 8044 23489 8072
rect 22787 8041 22799 8044
rect 22741 8035 22799 8041
rect 23477 8041 23489 8044
rect 23523 8072 23535 8075
rect 23842 8072 23848 8084
rect 23523 8044 23848 8072
rect 23523 8041 23535 8044
rect 23477 8035 23535 8041
rect 23842 8032 23848 8044
rect 23900 8032 23906 8084
rect 16898 7967 16956 7973
rect 17696 7976 18460 8004
rect 7926 7896 7932 7948
rect 7984 7936 7990 7948
rect 8021 7939 8079 7945
rect 8021 7936 8033 7939
rect 7984 7908 8033 7936
rect 7984 7896 7990 7908
rect 8021 7905 8033 7908
rect 8067 7936 8079 7939
rect 8067 7908 8248 7936
rect 8067 7905 8079 7908
rect 8021 7899 8079 7905
rect 1854 7828 1860 7880
rect 1912 7868 1918 7880
rect 2225 7871 2283 7877
rect 2225 7868 2237 7871
rect 1912 7840 2237 7868
rect 1912 7828 1918 7840
rect 2225 7837 2237 7840
rect 2271 7837 2283 7871
rect 2593 7871 2651 7877
rect 2593 7868 2605 7871
rect 2225 7831 2283 7837
rect 2516 7840 2605 7868
rect 2516 7812 2544 7840
rect 2593 7837 2605 7840
rect 2639 7837 2651 7871
rect 4154 7868 4160 7880
rect 4115 7840 4160 7868
rect 2593 7831 2651 7837
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7868 4491 7871
rect 5442 7868 5448 7880
rect 4479 7840 5448 7868
rect 4479 7837 4491 7840
rect 4433 7831 4491 7837
rect 2498 7760 2504 7812
rect 2556 7800 2562 7812
rect 4448 7800 4476 7831
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 6365 7871 6423 7877
rect 6365 7837 6377 7871
rect 6411 7868 6423 7871
rect 6546 7868 6552 7880
rect 6411 7840 6552 7868
rect 6411 7837 6423 7840
rect 6365 7831 6423 7837
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 8220 7868 8248 7908
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 8573 7939 8631 7945
rect 8573 7936 8585 7939
rect 8352 7908 8585 7936
rect 8352 7896 8358 7908
rect 8573 7905 8585 7908
rect 8619 7936 8631 7939
rect 8662 7936 8668 7948
rect 8619 7908 8668 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 8662 7896 8668 7908
rect 8720 7896 8726 7948
rect 15562 7896 15568 7948
rect 15620 7945 15626 7948
rect 15620 7939 15658 7945
rect 15646 7905 15658 7939
rect 15620 7899 15658 7905
rect 16577 7939 16635 7945
rect 16577 7905 16589 7939
rect 16623 7936 16635 7939
rect 17402 7936 17408 7948
rect 16623 7908 17408 7936
rect 16623 7905 16635 7908
rect 16577 7899 16635 7905
rect 15620 7896 15626 7899
rect 17402 7896 17408 7908
rect 17460 7936 17466 7948
rect 17696 7936 17724 7976
rect 21910 7964 21916 8016
rect 21968 8004 21974 8016
rect 22142 8007 22200 8013
rect 22142 8004 22154 8007
rect 21968 7976 22154 8004
rect 21968 7964 21974 7976
rect 22142 7973 22154 7976
rect 22188 7973 22200 8007
rect 22142 7967 22200 7973
rect 23658 7964 23664 8016
rect 23716 8004 23722 8016
rect 23753 8007 23811 8013
rect 23753 8004 23765 8007
rect 23716 7976 23765 8004
rect 23716 7964 23722 7976
rect 23753 7973 23765 7976
rect 23799 7973 23811 8007
rect 23753 7967 23811 7973
rect 18322 7936 18328 7948
rect 17460 7908 17724 7936
rect 18283 7908 18328 7936
rect 17460 7896 17466 7908
rect 18322 7896 18328 7908
rect 18380 7896 18386 7948
rect 18785 7939 18843 7945
rect 18785 7905 18797 7939
rect 18831 7905 18843 7939
rect 18785 7899 18843 7905
rect 25184 7939 25242 7945
rect 25184 7905 25196 7939
rect 25230 7936 25242 7939
rect 25774 7936 25780 7948
rect 25230 7908 25780 7936
rect 25230 7905 25242 7908
rect 25184 7899 25242 7905
rect 8754 7868 8760 7880
rect 8220 7840 8760 7868
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 9677 7871 9735 7877
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 9766 7868 9772 7880
rect 9723 7840 9772 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 9766 7828 9772 7840
rect 9824 7828 9830 7880
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 11296 7840 11437 7868
rect 11296 7828 11302 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 13998 7868 14004 7880
rect 13959 7840 14004 7868
rect 11425 7831 11483 7837
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 17310 7828 17316 7880
rect 17368 7868 17374 7880
rect 18800 7868 18828 7899
rect 25774 7896 25780 7908
rect 25832 7896 25838 7948
rect 17368 7840 18828 7868
rect 21821 7871 21879 7877
rect 17368 7828 17374 7840
rect 21821 7837 21833 7871
rect 21867 7868 21879 7871
rect 22002 7868 22008 7880
rect 21867 7840 22008 7868
rect 21867 7837 21879 7840
rect 21821 7831 21879 7837
rect 22002 7828 22008 7840
rect 22060 7828 22066 7880
rect 23661 7871 23719 7877
rect 23661 7837 23673 7871
rect 23707 7868 23719 7871
rect 25038 7868 25044 7880
rect 23707 7840 25044 7868
rect 23707 7837 23719 7840
rect 23661 7831 23719 7837
rect 25038 7828 25044 7840
rect 25096 7868 25102 7880
rect 25271 7871 25329 7877
rect 25271 7868 25283 7871
rect 25096 7840 25283 7868
rect 25096 7828 25102 7840
rect 25271 7837 25283 7840
rect 25317 7837 25329 7871
rect 25271 7831 25329 7837
rect 2556 7772 4476 7800
rect 7101 7803 7159 7809
rect 2556 7760 2562 7772
rect 7101 7769 7113 7803
rect 7147 7800 7159 7803
rect 8018 7800 8024 7812
rect 7147 7772 8024 7800
rect 7147 7769 7159 7772
rect 7101 7763 7159 7769
rect 8018 7760 8024 7772
rect 8076 7760 8082 7812
rect 14734 7760 14740 7812
rect 14792 7800 14798 7812
rect 16666 7800 16672 7812
rect 14792 7772 16672 7800
rect 14792 7760 14798 7772
rect 16666 7760 16672 7772
rect 16724 7760 16730 7812
rect 21361 7803 21419 7809
rect 21361 7769 21373 7803
rect 21407 7800 21419 7803
rect 21726 7800 21732 7812
rect 21407 7772 21732 7800
rect 21407 7769 21419 7772
rect 21361 7763 21419 7769
rect 21726 7760 21732 7772
rect 21784 7760 21790 7812
rect 24210 7800 24216 7812
rect 24171 7772 24216 7800
rect 24210 7760 24216 7772
rect 24268 7760 24274 7812
rect 1673 7735 1731 7741
rect 1673 7701 1685 7735
rect 1719 7732 1731 7735
rect 1762 7732 1768 7744
rect 1719 7704 1768 7732
rect 1719 7701 1731 7704
rect 1673 7695 1731 7701
rect 1762 7692 1768 7704
rect 1820 7692 1826 7744
rect 3602 7732 3608 7744
rect 3563 7704 3608 7732
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 5442 7732 5448 7744
rect 5403 7704 5448 7732
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 9398 7732 9404 7744
rect 9359 7704 9404 7732
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 9674 7692 9680 7744
rect 9732 7732 9738 7744
rect 10134 7732 10140 7744
rect 9732 7704 10140 7732
rect 9732 7692 9738 7704
rect 10134 7692 10140 7704
rect 10192 7732 10198 7744
rect 10597 7735 10655 7741
rect 10597 7732 10609 7735
rect 10192 7704 10609 7732
rect 10192 7692 10198 7704
rect 10597 7701 10609 7704
rect 10643 7701 10655 7735
rect 10597 7695 10655 7701
rect 11698 7692 11704 7744
rect 11756 7732 11762 7744
rect 12621 7735 12679 7741
rect 12621 7732 12633 7735
rect 11756 7704 12633 7732
rect 11756 7692 11762 7704
rect 12621 7701 12633 7704
rect 12667 7701 12679 7735
rect 12621 7695 12679 7701
rect 21637 7735 21695 7741
rect 21637 7701 21649 7735
rect 21683 7732 21695 7735
rect 21818 7732 21824 7744
rect 21683 7704 21824 7732
rect 21683 7701 21695 7704
rect 21637 7695 21695 7701
rect 21818 7692 21824 7704
rect 21876 7692 21882 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1670 7488 1676 7540
rect 1728 7537 1734 7540
rect 1728 7531 1777 7537
rect 1728 7497 1731 7531
rect 1765 7497 1777 7531
rect 1728 7491 1777 7497
rect 2225 7531 2283 7537
rect 2225 7497 2237 7531
rect 2271 7528 2283 7531
rect 2314 7528 2320 7540
rect 2271 7500 2320 7528
rect 2271 7497 2283 7500
rect 2225 7491 2283 7497
rect 1728 7488 1734 7491
rect 2314 7488 2320 7500
rect 2372 7488 2378 7540
rect 3878 7488 3884 7540
rect 3936 7528 3942 7540
rect 3973 7531 4031 7537
rect 3973 7528 3985 7531
rect 3936 7500 3985 7528
rect 3936 7488 3942 7500
rect 3973 7497 3985 7500
rect 4019 7497 4031 7531
rect 3973 7491 4031 7497
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4341 7531 4399 7537
rect 4341 7528 4353 7531
rect 4212 7500 4353 7528
rect 4212 7488 4218 7500
rect 4341 7497 4353 7500
rect 4387 7497 4399 7531
rect 4341 7491 4399 7497
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 6270 7528 6276 7540
rect 5951 7500 6276 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 8527 7531 8585 7537
rect 8527 7528 8539 7531
rect 8352 7500 8539 7528
rect 8352 7488 8358 7500
rect 8527 7497 8539 7500
rect 8573 7497 8585 7531
rect 8846 7528 8852 7540
rect 8807 7500 8852 7528
rect 8527 7491 8585 7497
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 11333 7531 11391 7537
rect 11333 7497 11345 7531
rect 11379 7528 11391 7531
rect 11422 7528 11428 7540
rect 11379 7500 11428 7528
rect 11379 7497 11391 7500
rect 11333 7491 11391 7497
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 13262 7488 13268 7540
rect 13320 7528 13326 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 13320 7500 13461 7528
rect 13320 7488 13326 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 15562 7488 15568 7540
rect 15620 7528 15626 7540
rect 16209 7531 16267 7537
rect 16209 7528 16221 7531
rect 15620 7500 16221 7528
rect 15620 7488 15626 7500
rect 16209 7497 16221 7500
rect 16255 7497 16267 7531
rect 16209 7491 16267 7497
rect 17083 7531 17141 7537
rect 17083 7497 17095 7531
rect 17129 7528 17141 7531
rect 17678 7528 17684 7540
rect 17129 7500 17684 7528
rect 17129 7497 17141 7500
rect 17083 7491 17141 7497
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 18322 7528 18328 7540
rect 18283 7500 18328 7528
rect 18322 7488 18328 7500
rect 18380 7528 18386 7540
rect 22830 7528 22836 7540
rect 18380 7500 19748 7528
rect 22791 7500 22836 7528
rect 18380 7488 18386 7500
rect 2332 7460 2360 7488
rect 3697 7463 3755 7469
rect 3697 7460 3709 7463
rect 2332 7432 3709 7460
rect 3697 7429 3709 7432
rect 3743 7429 3755 7463
rect 3697 7423 3755 7429
rect 10042 7420 10048 7472
rect 10100 7460 10106 7472
rect 10137 7463 10195 7469
rect 10137 7460 10149 7463
rect 10100 7432 10149 7460
rect 10100 7420 10106 7432
rect 10137 7429 10149 7432
rect 10183 7429 10195 7463
rect 10137 7423 10195 7429
rect 13630 7420 13636 7472
rect 13688 7460 13694 7472
rect 13688 7432 13768 7460
rect 13688 7420 13694 7432
rect 4890 7352 4896 7404
rect 4948 7392 4954 7404
rect 4985 7395 5043 7401
rect 4985 7392 4997 7395
rect 4948 7364 4997 7392
rect 4948 7352 4954 7364
rect 4985 7361 4997 7364
rect 5031 7392 5043 7395
rect 5442 7392 5448 7404
rect 5031 7364 5448 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7926 7392 7932 7404
rect 6972 7364 7932 7392
rect 6972 7352 6978 7364
rect 7926 7352 7932 7364
rect 7984 7392 7990 7404
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 7984 7364 8033 7392
rect 7984 7352 7990 7364
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 9766 7352 9772 7404
rect 9824 7392 9830 7404
rect 13740 7401 13768 7432
rect 17310 7420 17316 7472
rect 17368 7460 17374 7472
rect 17773 7463 17831 7469
rect 17773 7460 17785 7463
rect 17368 7432 17785 7460
rect 17368 7420 17374 7432
rect 17773 7429 17785 7432
rect 17819 7429 17831 7463
rect 17773 7423 17831 7429
rect 19150 7420 19156 7472
rect 19208 7460 19214 7472
rect 19245 7463 19303 7469
rect 19245 7460 19257 7463
rect 19208 7432 19257 7460
rect 19208 7420 19214 7432
rect 19245 7429 19257 7432
rect 19291 7429 19303 7463
rect 19245 7423 19303 7429
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 9824 7364 10885 7392
rect 9824 7352 9830 7364
rect 10873 7361 10885 7364
rect 10919 7361 10931 7395
rect 10873 7355 10931 7361
rect 13725 7395 13783 7401
rect 13725 7361 13737 7395
rect 13771 7361 13783 7395
rect 13998 7392 14004 7404
rect 13959 7364 14004 7392
rect 13725 7355 13783 7361
rect 13998 7352 14004 7364
rect 14056 7352 14062 7404
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7392 18751 7395
rect 19518 7392 19524 7404
rect 18739 7364 19524 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 19518 7352 19524 7364
rect 19576 7392 19582 7404
rect 19613 7395 19671 7401
rect 19613 7392 19625 7395
rect 19576 7364 19625 7392
rect 19576 7352 19582 7364
rect 19613 7361 19625 7364
rect 19659 7361 19671 7395
rect 19613 7355 19671 7361
rect 1648 7327 1706 7333
rect 1648 7293 1660 7327
rect 1694 7324 1706 7327
rect 2498 7324 2504 7336
rect 1694 7296 2504 7324
rect 1694 7293 1706 7296
rect 1648 7287 1706 7293
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 2777 7327 2835 7333
rect 2777 7293 2789 7327
rect 2823 7324 2835 7327
rect 3602 7324 3608 7336
rect 2823 7296 3608 7324
rect 2823 7293 2835 7296
rect 2777 7287 2835 7293
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 7098 7324 7104 7336
rect 6687 7296 7104 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 7282 7324 7288 7336
rect 7243 7296 7288 7324
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 8456 7327 8514 7333
rect 8456 7293 8468 7327
rect 8502 7324 8514 7327
rect 8846 7324 8852 7336
rect 8502 7296 8852 7324
rect 8502 7293 8514 7296
rect 8456 7287 8514 7293
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 11112 7296 11161 7324
rect 11112 7284 11118 7296
rect 11149 7293 11161 7296
rect 11195 7324 11207 7327
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11195 7296 11989 7324
rect 11195 7293 11207 7296
rect 11149 7287 11207 7293
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 12504 7327 12562 7333
rect 12504 7293 12516 7327
rect 12550 7293 12562 7327
rect 12504 7287 12562 7293
rect 2685 7259 2743 7265
rect 2685 7225 2697 7259
rect 2731 7256 2743 7259
rect 3139 7259 3197 7265
rect 3139 7256 3151 7259
rect 2731 7228 3151 7256
rect 2731 7225 2743 7228
rect 2685 7219 2743 7225
rect 3139 7225 3151 7228
rect 3185 7256 3197 7259
rect 3234 7256 3240 7268
rect 3185 7228 3240 7256
rect 3185 7225 3197 7228
rect 3139 7219 3197 7225
rect 3234 7216 3240 7228
rect 3292 7256 3298 7268
rect 4893 7259 4951 7265
rect 4893 7256 4905 7259
rect 3292 7228 4905 7256
rect 3292 7216 3298 7228
rect 4893 7225 4905 7228
rect 4939 7256 4951 7259
rect 5347 7259 5405 7265
rect 5347 7256 5359 7259
rect 4939 7228 5359 7256
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 5347 7225 5359 7228
rect 5393 7256 5405 7259
rect 5994 7256 6000 7268
rect 5393 7228 6000 7256
rect 5393 7225 5405 7228
rect 5347 7219 5405 7225
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 9582 7256 9588 7268
rect 9543 7228 9588 7256
rect 9582 7216 9588 7228
rect 9640 7216 9646 7268
rect 9674 7216 9680 7268
rect 9732 7256 9738 7268
rect 12519 7256 12547 7287
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 15197 7327 15255 7333
rect 15197 7324 15209 7327
rect 15068 7296 15209 7324
rect 15068 7284 15074 7296
rect 15197 7293 15209 7296
rect 15243 7324 15255 7327
rect 15378 7324 15384 7336
rect 15243 7296 15384 7324
rect 15243 7293 15255 7296
rect 15197 7287 15255 7293
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 15746 7324 15752 7336
rect 15707 7296 15752 7324
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 16850 7284 16856 7336
rect 16908 7324 16914 7336
rect 16980 7327 17038 7333
rect 16980 7324 16992 7327
rect 16908 7296 16992 7324
rect 16908 7284 16914 7296
rect 16980 7293 16992 7296
rect 17026 7324 17038 7327
rect 17405 7327 17463 7333
rect 17405 7324 17417 7327
rect 17026 7296 17417 7324
rect 17026 7293 17038 7296
rect 16980 7287 17038 7293
rect 17405 7293 17417 7296
rect 17451 7293 17463 7327
rect 19720 7324 19748 7500
rect 22830 7488 22836 7500
rect 22888 7488 22894 7540
rect 25038 7528 25044 7540
rect 24999 7500 25044 7528
rect 25038 7488 25044 7500
rect 25096 7488 25102 7540
rect 25130 7488 25136 7540
rect 25188 7528 25194 7540
rect 25363 7531 25421 7537
rect 25363 7528 25375 7531
rect 25188 7500 25375 7528
rect 25188 7488 25194 7500
rect 25363 7497 25375 7500
rect 25409 7497 25421 7531
rect 25774 7528 25780 7540
rect 25735 7500 25780 7528
rect 25363 7491 25421 7497
rect 25774 7488 25780 7500
rect 25832 7488 25838 7540
rect 21637 7395 21695 7401
rect 21637 7361 21649 7395
rect 21683 7392 21695 7395
rect 21818 7392 21824 7404
rect 21683 7364 21824 7392
rect 21683 7361 21695 7364
rect 21637 7355 21695 7361
rect 21818 7352 21824 7364
rect 21876 7352 21882 7404
rect 24578 7352 24584 7404
rect 24636 7392 24642 7404
rect 24636 7364 24900 7392
rect 24636 7352 24642 7364
rect 20165 7327 20223 7333
rect 20165 7324 20177 7327
rect 19720 7296 20177 7324
rect 17405 7287 17463 7293
rect 20165 7293 20177 7296
rect 20211 7324 20223 7327
rect 20254 7324 20260 7336
rect 20211 7296 20260 7324
rect 20211 7293 20223 7296
rect 20165 7287 20223 7293
rect 20254 7284 20260 7296
rect 20312 7284 20318 7336
rect 20622 7324 20628 7336
rect 20535 7296 20628 7324
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 21729 7327 21787 7333
rect 21729 7324 21741 7327
rect 21192 7296 21741 7324
rect 13446 7256 13452 7268
rect 9732 7228 9825 7256
rect 12519 7228 13452 7256
rect 9732 7216 9738 7228
rect 6914 7188 6920 7200
rect 6875 7160 6920 7188
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 9401 7191 9459 7197
rect 9401 7157 9413 7191
rect 9447 7188 9459 7191
rect 9692 7188 9720 7216
rect 13004 7200 13032 7228
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 13872 7228 13917 7256
rect 13872 7216 13878 7228
rect 13998 7216 14004 7268
rect 14056 7256 14062 7268
rect 14737 7259 14795 7265
rect 14737 7256 14749 7259
rect 14056 7228 14749 7256
rect 14056 7216 14062 7228
rect 14737 7225 14749 7228
rect 14783 7256 14795 7259
rect 15764 7256 15792 7284
rect 14783 7228 15792 7256
rect 14783 7225 14795 7228
rect 14737 7219 14795 7225
rect 18782 7216 18788 7268
rect 18840 7256 18846 7268
rect 18840 7228 18885 7256
rect 18840 7216 18846 7228
rect 19058 7216 19064 7268
rect 19116 7256 19122 7268
rect 19981 7259 20039 7265
rect 19981 7256 19993 7259
rect 19116 7228 19993 7256
rect 19116 7216 19122 7228
rect 19981 7225 19993 7228
rect 20027 7256 20039 7259
rect 20640 7256 20668 7284
rect 20027 7228 20668 7256
rect 20027 7225 20039 7228
rect 19981 7219 20039 7225
rect 21192 7200 21220 7296
rect 21729 7293 21741 7296
rect 21775 7293 21787 7327
rect 21729 7287 21787 7293
rect 22281 7327 22339 7333
rect 22281 7293 22293 7327
rect 22327 7324 22339 7327
rect 22830 7324 22836 7336
rect 22327 7296 22836 7324
rect 22327 7293 22339 7296
rect 22281 7287 22339 7293
rect 22830 7284 22836 7296
rect 22888 7284 22894 7336
rect 23382 7284 23388 7336
rect 23440 7324 23446 7336
rect 23661 7327 23719 7333
rect 23661 7324 23673 7327
rect 23440 7296 23673 7324
rect 23440 7284 23446 7296
rect 23661 7293 23673 7296
rect 23707 7293 23719 7327
rect 23661 7287 23719 7293
rect 24121 7327 24179 7333
rect 24121 7293 24133 7327
rect 24167 7324 24179 7327
rect 24673 7327 24731 7333
rect 24673 7324 24685 7327
rect 24167 7296 24685 7324
rect 24167 7293 24179 7296
rect 24121 7287 24179 7293
rect 24673 7293 24685 7296
rect 24719 7293 24731 7327
rect 24872 7324 24900 7364
rect 25260 7327 25318 7333
rect 25260 7324 25272 7327
rect 24872 7296 25272 7324
rect 24673 7287 24731 7293
rect 25260 7293 25272 7296
rect 25306 7324 25318 7327
rect 26053 7327 26111 7333
rect 26053 7324 26065 7327
rect 25306 7296 26065 7324
rect 25306 7293 25318 7296
rect 25260 7287 25318 7293
rect 26053 7293 26065 7296
rect 26099 7293 26111 7327
rect 26053 7287 26111 7293
rect 22848 7256 22876 7284
rect 24136 7256 24164 7287
rect 22848 7228 24164 7256
rect 9447 7160 9720 7188
rect 10597 7191 10655 7197
rect 9447 7157 9459 7160
rect 9401 7151 9459 7157
rect 10597 7157 10609 7191
rect 10643 7188 10655 7191
rect 11698 7188 11704 7200
rect 10643 7160 11704 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 12618 7197 12624 7200
rect 12575 7191 12624 7197
rect 12575 7157 12587 7191
rect 12621 7157 12624 7191
rect 12575 7151 12624 7157
rect 12618 7148 12624 7151
rect 12676 7148 12682 7200
rect 12986 7188 12992 7200
rect 12947 7160 12992 7188
rect 12986 7148 12992 7160
rect 13044 7148 13050 7200
rect 15010 7188 15016 7200
rect 14971 7160 15016 7188
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 15473 7191 15531 7197
rect 15473 7157 15485 7191
rect 15519 7188 15531 7191
rect 15654 7188 15660 7200
rect 15519 7160 15660 7188
rect 15519 7157 15531 7160
rect 15473 7151 15531 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 16669 7191 16727 7197
rect 16669 7157 16681 7191
rect 16715 7188 16727 7191
rect 16758 7188 16764 7200
rect 16715 7160 16764 7188
rect 16715 7157 16727 7160
rect 16669 7151 16727 7157
rect 16758 7148 16764 7160
rect 16816 7188 16822 7200
rect 17862 7188 17868 7200
rect 16816 7160 17868 7188
rect 16816 7148 16822 7160
rect 17862 7148 17868 7160
rect 17920 7148 17926 7200
rect 20162 7148 20168 7200
rect 20220 7188 20226 7200
rect 20257 7191 20315 7197
rect 20257 7188 20269 7191
rect 20220 7160 20269 7188
rect 20220 7148 20226 7160
rect 20257 7157 20269 7160
rect 20303 7157 20315 7191
rect 21174 7188 21180 7200
rect 21135 7160 21180 7188
rect 20257 7151 20315 7157
rect 21174 7148 21180 7160
rect 21232 7148 21238 7200
rect 21726 7148 21732 7200
rect 21784 7188 21790 7200
rect 21821 7191 21879 7197
rect 21821 7188 21833 7191
rect 21784 7160 21833 7188
rect 21784 7148 21790 7160
rect 21821 7157 21833 7160
rect 21867 7157 21879 7191
rect 23382 7188 23388 7200
rect 23343 7160 23388 7188
rect 21821 7151 21879 7157
rect 23382 7148 23388 7160
rect 23440 7148 23446 7200
rect 23750 7188 23756 7200
rect 23711 7160 23756 7188
rect 23750 7148 23756 7160
rect 23808 7148 23814 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1210 6944 1216 6996
rect 1268 6984 1274 6996
rect 1857 6987 1915 6993
rect 1857 6984 1869 6987
rect 1268 6956 1869 6984
rect 1268 6944 1274 6956
rect 1479 6857 1507 6956
rect 1857 6953 1869 6956
rect 1903 6953 1915 6987
rect 1857 6947 1915 6953
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 5537 6987 5595 6993
rect 5537 6984 5549 6987
rect 4304 6956 5549 6984
rect 4304 6944 4310 6956
rect 5537 6953 5549 6956
rect 5583 6953 5595 6987
rect 9766 6984 9772 6996
rect 9727 6956 9772 6984
rect 5537 6947 5595 6953
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 13725 6987 13783 6993
rect 13725 6953 13737 6987
rect 13771 6984 13783 6987
rect 13814 6984 13820 6996
rect 13771 6956 13820 6984
rect 13771 6953 13783 6956
rect 13725 6947 13783 6953
rect 13814 6944 13820 6956
rect 13872 6944 13878 6996
rect 17402 6984 17408 6996
rect 17363 6956 17408 6984
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 18782 6984 18788 6996
rect 18743 6956 18788 6984
rect 18782 6944 18788 6956
rect 18840 6984 18846 6996
rect 19061 6987 19119 6993
rect 19061 6984 19073 6987
rect 18840 6956 19073 6984
rect 18840 6944 18846 6956
rect 19061 6953 19073 6956
rect 19107 6953 19119 6987
rect 19061 6947 19119 6953
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 19751 6987 19809 6993
rect 19751 6984 19763 6987
rect 19576 6956 19763 6984
rect 19576 6944 19582 6956
rect 19751 6953 19763 6956
rect 19797 6953 19809 6987
rect 20254 6984 20260 6996
rect 20215 6956 20260 6984
rect 19751 6947 19809 6953
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 22738 6944 22744 6996
rect 22796 6984 22802 6996
rect 23290 6984 23296 6996
rect 22796 6956 23296 6984
rect 22796 6944 22802 6956
rect 23290 6944 23296 6956
rect 23348 6944 23354 6996
rect 23658 6944 23664 6996
rect 23716 6984 23722 6996
rect 24305 6987 24363 6993
rect 24305 6984 24317 6987
rect 23716 6956 24317 6984
rect 23716 6944 23722 6956
rect 24305 6953 24317 6956
rect 24351 6953 24363 6987
rect 25130 6984 25136 6996
rect 25091 6956 25136 6984
rect 24305 6947 24363 6953
rect 25130 6944 25136 6956
rect 25188 6944 25194 6996
rect 4890 6916 4896 6928
rect 4851 6888 4896 6916
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 6086 6925 6092 6928
rect 6083 6879 6092 6925
rect 6144 6916 6150 6928
rect 7650 6916 7656 6928
rect 6144 6888 6183 6916
rect 7611 6888 7656 6916
rect 6086 6876 6092 6879
rect 6144 6876 6150 6888
rect 7650 6876 7656 6888
rect 7708 6876 7714 6928
rect 9030 6876 9036 6928
rect 9088 6916 9094 6928
rect 12713 6919 12771 6925
rect 12713 6916 12725 6919
rect 9088 6888 9904 6916
rect 9088 6876 9094 6888
rect 1464 6851 1522 6857
rect 1464 6817 1476 6851
rect 1510 6817 1522 6851
rect 1464 6811 1522 6817
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6817 2467 6851
rect 2409 6811 2467 6817
rect 2556 6851 2614 6857
rect 2556 6817 2568 6851
rect 2602 6848 2614 6851
rect 2866 6848 2872 6860
rect 2602 6820 2872 6848
rect 2602 6817 2614 6820
rect 2556 6811 2614 6817
rect 2424 6712 2452 6811
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 3513 6851 3571 6857
rect 3513 6817 3525 6851
rect 3559 6848 3571 6851
rect 3970 6848 3976 6860
rect 3559 6820 3976 6848
rect 3559 6817 3571 6820
rect 3513 6811 3571 6817
rect 3970 6808 3976 6820
rect 4028 6848 4034 6860
rect 4433 6851 4491 6857
rect 4433 6848 4445 6851
rect 4028 6820 4445 6848
rect 4028 6808 4034 6820
rect 4433 6817 4445 6820
rect 4479 6848 4491 6851
rect 4522 6848 4528 6860
rect 4479 6820 4528 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 4706 6848 4712 6860
rect 4667 6820 4712 6848
rect 4706 6808 4712 6820
rect 4764 6808 4770 6860
rect 5534 6808 5540 6860
rect 5592 6848 5598 6860
rect 5721 6851 5779 6857
rect 5721 6848 5733 6851
rect 5592 6820 5733 6848
rect 5592 6808 5598 6820
rect 5721 6817 5733 6820
rect 5767 6817 5779 6851
rect 5721 6811 5779 6817
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 9876 6848 9904 6888
rect 12452 6888 12725 6916
rect 12452 6860 12480 6888
rect 12713 6885 12725 6888
rect 12759 6885 12771 6919
rect 12713 6879 12771 6885
rect 15746 6876 15752 6928
rect 15804 6916 15810 6928
rect 15804 6888 16620 6916
rect 15804 6876 15810 6888
rect 10137 6851 10195 6857
rect 10137 6848 10149 6851
rect 9732 6820 9777 6848
rect 9876 6820 10149 6848
rect 9732 6808 9738 6820
rect 10137 6817 10149 6820
rect 10183 6848 10195 6851
rect 10689 6851 10747 6857
rect 10689 6848 10701 6851
rect 10183 6820 10701 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10689 6817 10701 6820
rect 10735 6848 10747 6851
rect 10778 6848 10784 6860
rect 10735 6820 10784 6848
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 10778 6808 10784 6820
rect 10836 6808 10842 6860
rect 11292 6851 11350 6857
rect 11292 6817 11304 6851
rect 11338 6848 11350 6851
rect 11606 6848 11612 6860
rect 11338 6820 11612 6848
rect 11338 6817 11350 6820
rect 11292 6811 11350 6817
rect 11606 6808 11612 6820
rect 11664 6848 11670 6860
rect 12066 6848 12072 6860
rect 11664 6820 12072 6848
rect 11664 6808 11670 6820
rect 12066 6808 12072 6820
rect 12124 6808 12130 6860
rect 12434 6808 12440 6860
rect 12492 6808 12498 6860
rect 14252 6851 14310 6857
rect 14252 6817 14264 6851
rect 14298 6848 14310 6851
rect 14642 6848 14648 6860
rect 14298 6820 14648 6848
rect 14298 6817 14310 6820
rect 14252 6811 14310 6817
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 15286 6808 15292 6860
rect 15344 6857 15350 6860
rect 15470 6857 15476 6860
rect 15344 6851 15382 6857
rect 15370 6817 15382 6851
rect 15344 6811 15382 6817
rect 15427 6851 15476 6857
rect 15427 6817 15439 6851
rect 15473 6817 15476 6851
rect 15427 6811 15476 6817
rect 15344 6808 15350 6811
rect 15470 6808 15476 6811
rect 15528 6808 15534 6860
rect 16482 6848 16488 6860
rect 16443 6820 16488 6848
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 16592 6848 16620 6888
rect 17862 6876 17868 6928
rect 17920 6916 17926 6928
rect 18186 6919 18244 6925
rect 18186 6916 18198 6919
rect 17920 6888 18198 6916
rect 17920 6876 17926 6888
rect 18186 6885 18198 6888
rect 18232 6885 18244 6919
rect 18186 6879 18244 6885
rect 21818 6876 21824 6928
rect 21876 6925 21882 6928
rect 21876 6919 21924 6925
rect 21876 6885 21878 6919
rect 21912 6885 21924 6919
rect 23477 6919 23535 6925
rect 23477 6916 23489 6919
rect 21876 6879 21924 6885
rect 23216 6888 23489 6916
rect 21876 6876 21882 6879
rect 16758 6848 16764 6860
rect 16592 6820 16764 6848
rect 16758 6808 16764 6820
rect 16816 6808 16822 6860
rect 19426 6808 19432 6860
rect 19484 6848 19490 6860
rect 19648 6851 19706 6857
rect 19648 6848 19660 6851
rect 19484 6820 19660 6848
rect 19484 6808 19490 6820
rect 19648 6817 19660 6820
rect 19694 6817 19706 6851
rect 23216 6848 23244 6888
rect 23477 6885 23489 6888
rect 23523 6885 23535 6919
rect 23477 6879 23535 6885
rect 19648 6811 19706 6817
rect 23124 6820 23244 6848
rect 24029 6851 24087 6857
rect 2682 6740 2688 6792
rect 2740 6780 2746 6792
rect 2777 6783 2835 6789
rect 2777 6780 2789 6783
rect 2740 6752 2789 6780
rect 2740 6740 2746 6752
rect 2777 6749 2789 6752
rect 2823 6749 2835 6783
rect 2958 6780 2964 6792
rect 2919 6752 2964 6780
rect 2777 6743 2835 6749
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 4724 6780 4752 6808
rect 6917 6783 6975 6789
rect 6917 6780 6929 6783
rect 4724 6752 6929 6780
rect 6917 6749 6929 6752
rect 6963 6780 6975 6783
rect 7282 6780 7288 6792
rect 6963 6752 7288 6780
rect 6963 6749 6975 6752
rect 6917 6743 6975 6749
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7374 6740 7380 6792
rect 7432 6780 7438 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7432 6752 7573 6780
rect 7432 6740 7438 6752
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 8018 6780 8024 6792
rect 7979 6752 8024 6780
rect 7561 6743 7619 6749
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8846 6780 8852 6792
rect 8807 6752 8852 6780
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6780 9551 6783
rect 9582 6780 9588 6792
rect 9539 6752 9588 6780
rect 9539 6749 9551 6752
rect 9493 6743 9551 6749
rect 9582 6740 9588 6752
rect 9640 6780 9646 6792
rect 11379 6783 11437 6789
rect 11379 6780 11391 6783
rect 9640 6752 11391 6780
rect 9640 6740 9646 6752
rect 11379 6749 11391 6752
rect 11425 6749 11437 6783
rect 12618 6780 12624 6792
rect 12531 6752 12624 6780
rect 11379 6743 11437 6749
rect 12618 6740 12624 6752
rect 12676 6780 12682 6792
rect 13078 6780 13084 6792
rect 12676 6752 13084 6780
rect 12676 6740 12682 6752
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 17037 6783 17095 6789
rect 17037 6749 17049 6783
rect 17083 6780 17095 6783
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 17083 6752 17877 6780
rect 17083 6749 17095 6752
rect 17037 6743 17095 6749
rect 17865 6749 17877 6752
rect 17911 6780 17923 6783
rect 18414 6780 18420 6792
rect 17911 6752 18420 6780
rect 17911 6749 17923 6752
rect 17865 6743 17923 6749
rect 18414 6740 18420 6752
rect 18472 6740 18478 6792
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6780 21603 6783
rect 22370 6780 22376 6792
rect 21591 6752 22376 6780
rect 21591 6749 21603 6752
rect 21545 6743 21603 6749
rect 22370 6740 22376 6752
rect 22428 6740 22434 6792
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 2424 6684 3801 6712
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 3789 6675 3847 6681
rect 6641 6715 6699 6721
rect 6641 6681 6653 6715
rect 6687 6712 6699 6715
rect 7650 6712 7656 6724
rect 6687 6684 7656 6712
rect 6687 6681 6699 6684
rect 6641 6675 6699 6681
rect 1535 6647 1593 6653
rect 1535 6613 1547 6647
rect 1581 6644 1593 6647
rect 1762 6644 1768 6656
rect 1581 6616 1768 6644
rect 1581 6613 1593 6616
rect 1535 6607 1593 6613
rect 1762 6604 1768 6616
rect 1820 6604 1826 6656
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2685 6647 2743 6653
rect 2685 6613 2697 6647
rect 2731 6644 2743 6647
rect 2958 6644 2964 6656
rect 2731 6616 2964 6644
rect 2731 6613 2743 6616
rect 2685 6607 2743 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 3804 6644 3832 6675
rect 7650 6672 7656 6684
rect 7708 6672 7714 6724
rect 9674 6672 9680 6724
rect 9732 6712 9738 6724
rect 9950 6712 9956 6724
rect 9732 6684 9956 6712
rect 9732 6672 9738 6684
rect 9950 6672 9956 6684
rect 10008 6712 10014 6724
rect 10870 6712 10876 6724
rect 10008 6684 10876 6712
rect 10008 6672 10014 6684
rect 10870 6672 10876 6684
rect 10928 6672 10934 6724
rect 13170 6712 13176 6724
rect 13131 6684 13176 6712
rect 13170 6672 13176 6684
rect 13228 6672 13234 6724
rect 23124 6721 23152 6820
rect 24029 6817 24041 6851
rect 24075 6848 24087 6851
rect 24210 6848 24216 6860
rect 24075 6820 24216 6848
rect 24075 6817 24087 6820
rect 24029 6811 24087 6817
rect 24210 6808 24216 6820
rect 24268 6808 24274 6860
rect 24670 6848 24676 6860
rect 24631 6820 24676 6848
rect 24670 6808 24676 6820
rect 24728 6808 24734 6860
rect 24854 6848 24860 6860
rect 24815 6820 24860 6848
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 25314 6808 25320 6860
rect 25372 6848 25378 6860
rect 25409 6851 25467 6857
rect 25409 6848 25421 6851
rect 25372 6820 25421 6848
rect 25372 6808 25378 6820
rect 25409 6817 25421 6820
rect 25455 6848 25467 6851
rect 25866 6848 25872 6860
rect 25455 6820 25872 6848
rect 25455 6817 25467 6820
rect 25409 6811 25467 6817
rect 25866 6808 25872 6820
rect 25924 6808 25930 6860
rect 23385 6783 23443 6789
rect 23385 6749 23397 6783
rect 23431 6780 23443 6783
rect 24688 6780 24716 6808
rect 23431 6752 24716 6780
rect 24872 6780 24900 6808
rect 25590 6780 25596 6792
rect 24872 6752 25596 6780
rect 23431 6749 23443 6752
rect 23385 6743 23443 6749
rect 25590 6740 25596 6752
rect 25648 6740 25654 6792
rect 22465 6715 22523 6721
rect 22465 6681 22477 6715
rect 22511 6712 22523 6715
rect 23109 6715 23167 6721
rect 23109 6712 23121 6715
rect 22511 6684 23121 6712
rect 22511 6681 22523 6684
rect 22465 6675 22523 6681
rect 23109 6681 23121 6684
rect 23155 6681 23167 6715
rect 23109 6675 23167 6681
rect 3878 6644 3884 6656
rect 3804 6616 3884 6644
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 5166 6644 5172 6656
rect 5127 6616 5172 6644
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 7282 6644 7288 6656
rect 7243 6616 7288 6644
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 8662 6644 8668 6656
rect 8619 6616 8668 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 8662 6604 8668 6616
rect 8720 6604 8726 6656
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11701 6647 11759 6653
rect 11701 6644 11713 6647
rect 11296 6616 11713 6644
rect 11296 6604 11302 6616
rect 11701 6613 11713 6616
rect 11747 6613 11759 6647
rect 11701 6607 11759 6613
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 14093 6647 14151 6653
rect 14093 6644 14105 6647
rect 13872 6616 14105 6644
rect 13872 6604 13878 6616
rect 14093 6613 14105 6616
rect 14139 6644 14151 6647
rect 14323 6647 14381 6653
rect 14323 6644 14335 6647
rect 14139 6616 14335 6644
rect 14139 6613 14151 6616
rect 14093 6607 14151 6613
rect 14323 6613 14335 6616
rect 14369 6613 14381 6647
rect 15746 6644 15752 6656
rect 15707 6616 15752 6644
rect 14323 6607 14381 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 16209 6647 16267 6653
rect 16209 6613 16221 6647
rect 16255 6644 16267 6647
rect 16390 6644 16396 6656
rect 16255 6616 16396 6644
rect 16255 6613 16267 6616
rect 16209 6607 16267 6613
rect 16390 6604 16396 6616
rect 16448 6604 16454 6656
rect 17773 6647 17831 6653
rect 17773 6613 17785 6647
rect 17819 6644 17831 6647
rect 18138 6644 18144 6656
rect 17819 6616 18144 6644
rect 17819 6613 17831 6616
rect 17773 6607 17831 6613
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 21453 6647 21511 6653
rect 21453 6613 21465 6647
rect 21499 6644 21511 6647
rect 21542 6644 21548 6656
rect 21499 6616 21548 6644
rect 21499 6613 21511 6616
rect 21453 6607 21511 6613
rect 21542 6604 21548 6616
rect 21600 6604 21606 6656
rect 22002 6604 22008 6656
rect 22060 6644 22066 6656
rect 22833 6647 22891 6653
rect 22833 6644 22845 6647
rect 22060 6616 22845 6644
rect 22060 6604 22066 6616
rect 22833 6613 22845 6616
rect 22879 6644 22891 6647
rect 23750 6644 23756 6656
rect 22879 6616 23756 6644
rect 22879 6613 22891 6616
rect 22833 6607 22891 6613
rect 23750 6604 23756 6616
rect 23808 6604 23814 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 2866 6440 2872 6452
rect 2823 6412 2872 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 2866 6400 2872 6412
rect 2924 6400 2930 6452
rect 2958 6400 2964 6452
rect 3016 6440 3022 6452
rect 3053 6443 3111 6449
rect 3053 6440 3065 6443
rect 3016 6412 3065 6440
rect 3016 6400 3022 6412
rect 3053 6409 3065 6412
rect 3099 6409 3111 6443
rect 4706 6440 4712 6452
rect 4667 6412 4712 6440
rect 3053 6403 3111 6409
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 6181 6443 6239 6449
rect 6181 6440 6193 6443
rect 5592 6412 6193 6440
rect 5592 6400 5598 6412
rect 6181 6409 6193 6412
rect 6227 6409 6239 6443
rect 7374 6440 7380 6452
rect 7335 6412 7380 6440
rect 6181 6403 6239 6409
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 8481 6443 8539 6449
rect 8481 6440 8493 6443
rect 7708 6412 8493 6440
rect 7708 6400 7714 6412
rect 8481 6409 8493 6412
rect 8527 6409 8539 6443
rect 9030 6440 9036 6452
rect 8991 6412 9036 6440
rect 8481 6403 8539 6409
rect 9030 6400 9036 6412
rect 9088 6400 9094 6452
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 9401 6443 9459 6449
rect 9401 6440 9413 6443
rect 9364 6412 9413 6440
rect 9364 6400 9370 6412
rect 9401 6409 9413 6412
rect 9447 6440 9459 6443
rect 9674 6440 9680 6452
rect 9447 6412 9680 6440
rect 9447 6409 9459 6412
rect 9401 6403 9459 6409
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 11606 6440 11612 6452
rect 11567 6412 11612 6440
rect 11606 6400 11612 6412
rect 11664 6400 11670 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 12434 6440 12440 6452
rect 12299 6412 12440 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 14642 6400 14648 6452
rect 14700 6440 14706 6452
rect 14737 6443 14795 6449
rect 14737 6440 14749 6443
rect 14700 6412 14749 6440
rect 14700 6400 14706 6412
rect 14737 6409 14749 6412
rect 14783 6409 14795 6443
rect 14737 6403 14795 6409
rect 15197 6443 15255 6449
rect 15197 6409 15209 6443
rect 15243 6440 15255 6443
rect 15286 6440 15292 6452
rect 15243 6412 15292 6440
rect 15243 6409 15255 6412
rect 15197 6403 15255 6409
rect 15286 6400 15292 6412
rect 15344 6400 15350 6452
rect 16393 6443 16451 6449
rect 16393 6409 16405 6443
rect 16439 6440 16451 6443
rect 16482 6440 16488 6452
rect 16439 6412 16488 6440
rect 16439 6409 16451 6412
rect 16393 6403 16451 6409
rect 16482 6400 16488 6412
rect 16540 6400 16546 6452
rect 16942 6400 16948 6452
rect 17000 6449 17006 6452
rect 17000 6443 17049 6449
rect 17000 6409 17003 6443
rect 17037 6409 17049 6443
rect 17000 6403 17049 6409
rect 17000 6400 17006 6403
rect 19426 6400 19432 6452
rect 19484 6440 19490 6452
rect 19613 6443 19671 6449
rect 19613 6440 19625 6443
rect 19484 6412 19625 6440
rect 19484 6400 19490 6412
rect 19613 6409 19625 6412
rect 19659 6409 19671 6443
rect 19613 6403 19671 6409
rect 22830 6400 22836 6452
rect 22888 6440 22894 6452
rect 23017 6443 23075 6449
rect 23017 6440 23029 6443
rect 22888 6412 23029 6440
rect 22888 6400 22894 6412
rect 23017 6409 23029 6412
rect 23063 6409 23075 6443
rect 23017 6403 23075 6409
rect 13265 6375 13323 6381
rect 13265 6341 13277 6375
rect 13311 6372 13323 6375
rect 16022 6372 16028 6384
rect 13311 6344 16028 6372
rect 13311 6341 13323 6344
rect 13265 6335 13323 6341
rect 2409 6307 2467 6313
rect 2409 6273 2421 6307
rect 2455 6304 2467 6307
rect 2682 6304 2688 6316
rect 2455 6276 2688 6304
rect 2455 6273 2467 6276
rect 2409 6267 2467 6273
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 3602 6264 3608 6316
rect 3660 6304 3666 6316
rect 3789 6307 3847 6313
rect 3789 6304 3801 6307
rect 3660 6276 3801 6304
rect 3660 6264 3666 6276
rect 3789 6273 3801 6276
rect 3835 6273 3847 6307
rect 4890 6304 4896 6316
rect 4851 6276 4896 6304
rect 3789 6267 3847 6273
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6304 5595 6307
rect 7006 6304 7012 6316
rect 5583 6276 7012 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 7006 6264 7012 6276
rect 7064 6304 7070 6316
rect 7558 6304 7564 6316
rect 7064 6276 7564 6304
rect 7064 6264 7070 6276
rect 7558 6264 7564 6276
rect 7616 6264 7622 6316
rect 8018 6304 8024 6316
rect 7979 6276 8024 6304
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 11238 6304 11244 6316
rect 11199 6276 11244 6304
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 2317 6239 2375 6245
rect 2317 6205 2329 6239
rect 2363 6236 2375 6239
rect 2498 6236 2504 6248
rect 2363 6208 2504 6236
rect 2363 6205 2375 6208
rect 2317 6199 2375 6205
rect 2498 6196 2504 6208
rect 2556 6196 2562 6248
rect 3513 6239 3571 6245
rect 3513 6205 3525 6239
rect 3559 6205 3571 6239
rect 3513 6199 3571 6205
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6236 3755 6239
rect 3970 6236 3976 6248
rect 3743 6208 3976 6236
rect 3743 6205 3755 6208
rect 3697 6199 3755 6205
rect 3528 6168 3556 6199
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 4341 6239 4399 6245
rect 4341 6205 4353 6239
rect 4387 6236 4399 6239
rect 4522 6236 4528 6248
rect 4387 6208 4528 6236
rect 4387 6205 4399 6208
rect 4341 6199 4399 6205
rect 4356 6168 4384 6199
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 8202 6196 8208 6248
rect 8260 6236 8266 6248
rect 9493 6239 9551 6245
rect 9493 6236 9505 6239
rect 8260 6208 9505 6236
rect 8260 6196 8266 6208
rect 9493 6205 9505 6208
rect 9539 6236 9551 6239
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9539 6208 9965 6236
rect 9539 6205 9551 6208
rect 9493 6199 9551 6205
rect 9953 6205 9965 6208
rect 9999 6205 10011 6239
rect 10502 6236 10508 6248
rect 9953 6199 10011 6205
rect 10336 6208 10508 6236
rect 3528 6140 4384 6168
rect 4985 6171 5043 6177
rect 4985 6137 4997 6171
rect 5031 6168 5043 6171
rect 5166 6168 5172 6180
rect 5031 6140 5172 6168
rect 5031 6137 5043 6140
rect 4985 6131 5043 6137
rect 5166 6128 5172 6140
rect 5224 6128 5230 6180
rect 6641 6171 6699 6177
rect 6641 6137 6653 6171
rect 6687 6168 6699 6171
rect 7653 6171 7711 6177
rect 6687 6140 7512 6168
rect 6687 6137 6699 6140
rect 6641 6131 6699 6137
rect 5905 6103 5963 6109
rect 5905 6069 5917 6103
rect 5951 6100 5963 6103
rect 5994 6100 6000 6112
rect 5951 6072 6000 6100
rect 5951 6069 5963 6072
rect 5905 6063 5963 6069
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 7484 6100 7512 6140
rect 7653 6137 7665 6171
rect 7699 6137 7711 6171
rect 7653 6131 7711 6137
rect 7668 6100 7696 6131
rect 7926 6100 7932 6112
rect 7484 6072 7932 6100
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 9766 6100 9772 6112
rect 9723 6072 9772 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10134 6060 10140 6112
rect 10192 6100 10198 6112
rect 10336 6109 10364 6208
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 10778 6196 10784 6248
rect 10836 6236 10842 6248
rect 12802 6245 12808 6248
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 10836 6208 10977 6236
rect 10836 6196 10842 6208
rect 10965 6205 10977 6208
rect 11011 6205 11023 6239
rect 10965 6199 11023 6205
rect 12764 6239 12808 6245
rect 12764 6205 12776 6239
rect 12860 6236 12866 6248
rect 13280 6236 13308 6335
rect 16022 6332 16028 6344
rect 16080 6332 16086 6384
rect 13814 6304 13820 6316
rect 13775 6276 13820 6304
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 14182 6304 14188 6316
rect 14143 6276 14188 6304
rect 14182 6264 14188 6276
rect 14240 6264 14246 6316
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6304 15439 6307
rect 16390 6304 16396 6316
rect 15427 6276 16396 6304
rect 15427 6273 15439 6276
rect 15381 6267 15439 6273
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 16758 6304 16764 6316
rect 16671 6276 16764 6304
rect 16758 6264 16764 6276
rect 16816 6304 16822 6316
rect 23032 6304 23060 6403
rect 23382 6332 23388 6384
rect 23440 6372 23446 6384
rect 23477 6375 23535 6381
rect 23477 6372 23489 6375
rect 23440 6344 23489 6372
rect 23440 6332 23446 6344
rect 23477 6341 23489 6344
rect 23523 6341 23535 6375
rect 23477 6335 23535 6341
rect 16816 6276 20484 6304
rect 23032 6276 24164 6304
rect 16816 6264 16822 6276
rect 20456 6248 20484 6276
rect 12860 6208 13308 6236
rect 16920 6239 16978 6245
rect 12764 6199 12808 6205
rect 12802 6196 12808 6199
rect 12860 6196 12866 6208
rect 16920 6205 16932 6239
rect 16966 6236 16978 6239
rect 18138 6236 18144 6248
rect 16966 6208 17448 6236
rect 18051 6208 18144 6236
rect 16966 6205 16978 6208
rect 16920 6199 16978 6205
rect 13909 6171 13967 6177
rect 13909 6137 13921 6171
rect 13955 6137 13967 6171
rect 13909 6131 13967 6137
rect 10321 6103 10379 6109
rect 10321 6100 10333 6103
rect 10192 6072 10333 6100
rect 10192 6060 10198 6072
rect 10321 6069 10333 6072
rect 10367 6069 10379 6103
rect 10321 6063 10379 6069
rect 12851 6103 12909 6109
rect 12851 6069 12863 6103
rect 12897 6100 12909 6103
rect 13446 6100 13452 6112
rect 12897 6072 13452 6100
rect 12897 6069 12909 6072
rect 12851 6063 12909 6069
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 13633 6103 13691 6109
rect 13633 6069 13645 6103
rect 13679 6100 13691 6103
rect 13924 6100 13952 6131
rect 14642 6128 14648 6180
rect 14700 6168 14706 6180
rect 15473 6171 15531 6177
rect 14700 6140 15240 6168
rect 14700 6128 14706 6140
rect 14660 6100 14688 6128
rect 13679 6072 14688 6100
rect 15212 6100 15240 6140
rect 15473 6137 15485 6171
rect 15519 6168 15531 6171
rect 15746 6168 15752 6180
rect 15519 6140 15752 6168
rect 15519 6137 15531 6140
rect 15473 6131 15531 6137
rect 15488 6100 15516 6131
rect 15746 6128 15752 6140
rect 15804 6128 15810 6180
rect 16025 6171 16083 6177
rect 16025 6137 16037 6171
rect 16071 6168 16083 6171
rect 16206 6168 16212 6180
rect 16071 6140 16212 6168
rect 16071 6137 16083 6140
rect 16025 6131 16083 6137
rect 16206 6128 16212 6140
rect 16264 6128 16270 6180
rect 17420 6112 17448 6208
rect 18138 6196 18144 6208
rect 18196 6236 18202 6248
rect 20162 6236 20168 6248
rect 18196 6208 18644 6236
rect 20123 6208 20168 6236
rect 18196 6196 18202 6208
rect 18462 6171 18520 6177
rect 18462 6137 18474 6171
rect 18508 6137 18520 6171
rect 18616 6168 18644 6208
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 20438 6236 20444 6248
rect 20399 6208 20444 6236
rect 20438 6196 20444 6208
rect 20496 6196 20502 6248
rect 21542 6236 21548 6248
rect 21503 6208 21548 6236
rect 21542 6196 21548 6208
rect 21600 6196 21606 6248
rect 23382 6196 23388 6248
rect 23440 6236 23446 6248
rect 23661 6239 23719 6245
rect 23661 6236 23673 6239
rect 23440 6208 23673 6236
rect 23440 6196 23446 6208
rect 23661 6205 23673 6208
rect 23707 6236 23719 6239
rect 23842 6236 23848 6248
rect 23707 6208 23848 6236
rect 23707 6205 23719 6208
rect 23661 6199 23719 6205
rect 23842 6196 23848 6208
rect 23900 6196 23906 6248
rect 24136 6245 24164 6276
rect 24121 6239 24179 6245
rect 24121 6205 24133 6239
rect 24167 6205 24179 6239
rect 25222 6236 25228 6248
rect 25183 6208 25228 6236
rect 24121 6199 24179 6205
rect 25222 6196 25228 6208
rect 25280 6236 25286 6248
rect 25777 6239 25835 6245
rect 25777 6236 25789 6239
rect 25280 6208 25789 6236
rect 25280 6196 25286 6208
rect 25777 6205 25789 6208
rect 25823 6205 25835 6239
rect 25777 6199 25835 6205
rect 18616 6140 20024 6168
rect 18462 6131 18520 6137
rect 17402 6100 17408 6112
rect 15212 6072 15516 6100
rect 17363 6072 17408 6100
rect 13679 6069 13691 6072
rect 13633 6063 13691 6069
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 17862 6100 17868 6112
rect 17823 6072 17868 6100
rect 17862 6060 17868 6072
rect 17920 6100 17926 6112
rect 18477 6100 18505 6131
rect 17920 6072 18505 6100
rect 19061 6103 19119 6109
rect 17920 6060 17926 6072
rect 19061 6069 19073 6103
rect 19107 6100 19119 6103
rect 19242 6100 19248 6112
rect 19107 6072 19248 6100
rect 19107 6069 19119 6072
rect 19061 6063 19119 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 19996 6109 20024 6140
rect 20714 6128 20720 6180
rect 20772 6168 20778 6180
rect 20990 6168 20996 6180
rect 20772 6140 20996 6168
rect 20772 6128 20778 6140
rect 20990 6128 20996 6140
rect 21048 6128 21054 6180
rect 21818 6168 21824 6180
rect 21376 6140 21824 6168
rect 19981 6103 20039 6109
rect 19981 6069 19993 6103
rect 20027 6069 20039 6103
rect 21082 6100 21088 6112
rect 21043 6072 21088 6100
rect 19981 6063 20039 6069
rect 21082 6060 21088 6072
rect 21140 6100 21146 6112
rect 21376 6109 21404 6140
rect 21818 6128 21824 6140
rect 21876 6177 21882 6180
rect 21876 6171 21924 6177
rect 21876 6137 21878 6171
rect 21912 6137 21924 6171
rect 21876 6131 21924 6137
rect 21876 6128 21882 6131
rect 21361 6103 21419 6109
rect 21361 6100 21373 6103
rect 21140 6072 21373 6100
rect 21140 6060 21146 6072
rect 21361 6069 21373 6072
rect 21407 6069 21419 6103
rect 22462 6100 22468 6112
rect 22423 6072 22468 6100
rect 21361 6063 21419 6069
rect 22462 6060 22468 6072
rect 22520 6060 22526 6112
rect 23750 6100 23756 6112
rect 23711 6072 23756 6100
rect 23750 6060 23756 6072
rect 23808 6060 23814 6112
rect 24854 6100 24860 6112
rect 24815 6072 24860 6100
rect 24854 6060 24860 6072
rect 24912 6060 24918 6112
rect 25409 6103 25467 6109
rect 25409 6069 25421 6103
rect 25455 6100 25467 6103
rect 26510 6100 26516 6112
rect 25455 6072 26516 6100
rect 25455 6069 25467 6072
rect 25409 6063 25467 6069
rect 26510 6060 26516 6072
rect 26568 6060 26574 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1578 5905 1584 5908
rect 1535 5899 1584 5905
rect 1535 5865 1547 5899
rect 1581 5865 1584 5899
rect 1535 5859 1584 5865
rect 1578 5856 1584 5859
rect 1636 5856 1642 5908
rect 1949 5899 2007 5905
rect 1949 5865 1961 5899
rect 1995 5896 2007 5899
rect 2498 5896 2504 5908
rect 1995 5868 2504 5896
rect 1995 5865 2007 5868
rect 1949 5859 2007 5865
rect 2498 5856 2504 5868
rect 2556 5856 2562 5908
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 5261 5899 5319 5905
rect 5261 5896 5273 5899
rect 5224 5868 5273 5896
rect 5224 5856 5230 5868
rect 5261 5865 5273 5868
rect 5307 5865 5319 5899
rect 6270 5896 6276 5908
rect 6231 5868 6276 5896
rect 5261 5859 5319 5865
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 6914 5896 6920 5908
rect 6875 5868 6920 5896
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7926 5896 7932 5908
rect 7887 5868 7932 5896
rect 7926 5856 7932 5868
rect 7984 5856 7990 5908
rect 10962 5896 10968 5908
rect 10923 5868 10968 5896
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 13446 5896 13452 5908
rect 13407 5868 13452 5896
rect 13446 5856 13452 5868
rect 13504 5896 13510 5908
rect 16209 5899 16267 5905
rect 13504 5868 13768 5896
rect 13504 5856 13510 5868
rect 3145 5831 3203 5837
rect 3145 5797 3157 5831
rect 3191 5828 3203 5831
rect 3786 5828 3792 5840
rect 3191 5800 3792 5828
rect 3191 5797 3203 5800
rect 3145 5791 3203 5797
rect 3786 5788 3792 5800
rect 3844 5788 3850 5840
rect 4522 5788 4528 5840
rect 4580 5828 4586 5840
rect 4703 5831 4761 5837
rect 4703 5828 4715 5831
rect 4580 5800 4715 5828
rect 4580 5788 4586 5800
rect 4703 5797 4715 5800
rect 4749 5828 4761 5831
rect 5994 5828 6000 5840
rect 4749 5800 6000 5828
rect 4749 5797 4761 5800
rect 4703 5791 4761 5797
rect 5994 5788 6000 5800
rect 6052 5788 6058 5840
rect 7371 5831 7429 5837
rect 7371 5797 7383 5831
rect 7417 5828 7429 5831
rect 7417 5800 7512 5828
rect 7417 5797 7429 5800
rect 7371 5791 7429 5797
rect 1118 5720 1124 5772
rect 1176 5760 1182 5772
rect 1432 5763 1490 5769
rect 1432 5760 1444 5763
rect 1176 5732 1444 5760
rect 1176 5720 1182 5732
rect 1432 5729 1444 5732
rect 1478 5729 1490 5763
rect 1432 5723 1490 5729
rect 2314 5720 2320 5772
rect 2372 5760 2378 5772
rect 2409 5763 2467 5769
rect 2409 5760 2421 5763
rect 2372 5732 2421 5760
rect 2372 5720 2378 5732
rect 2409 5729 2421 5732
rect 2455 5760 2467 5763
rect 2498 5760 2504 5772
rect 2455 5732 2504 5760
rect 2455 5729 2467 5732
rect 2409 5723 2467 5729
rect 2498 5720 2504 5732
rect 2556 5720 2562 5772
rect 7484 5760 7512 5800
rect 7558 5788 7564 5840
rect 7616 5828 7622 5840
rect 8205 5831 8263 5837
rect 8205 5828 8217 5831
rect 7616 5800 8217 5828
rect 7616 5788 7622 5800
rect 8205 5797 8217 5800
rect 8251 5797 8263 5831
rect 13078 5828 13084 5840
rect 13039 5800 13084 5828
rect 8205 5791 8263 5797
rect 13078 5788 13084 5800
rect 13136 5788 13142 5840
rect 13740 5837 13768 5868
rect 16209 5865 16221 5899
rect 16255 5896 16267 5899
rect 18414 5896 18420 5908
rect 16255 5868 17264 5896
rect 18375 5868 18420 5896
rect 16255 5865 16267 5868
rect 16209 5859 16267 5865
rect 17236 5840 17264 5868
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 19981 5899 20039 5905
rect 19981 5865 19993 5899
rect 20027 5896 20039 5899
rect 20162 5896 20168 5908
rect 20027 5868 20168 5896
rect 20027 5865 20039 5868
rect 19981 5859 20039 5865
rect 20162 5856 20168 5868
rect 20220 5856 20226 5908
rect 20990 5896 20996 5908
rect 20951 5868 20996 5896
rect 20990 5856 20996 5868
rect 21048 5856 21054 5908
rect 23474 5856 23480 5908
rect 23532 5896 23538 5908
rect 23750 5896 23756 5908
rect 23532 5868 23756 5896
rect 23532 5856 23538 5868
rect 23750 5856 23756 5868
rect 23808 5856 23814 5908
rect 24210 5896 24216 5908
rect 24171 5868 24216 5896
rect 24210 5856 24216 5868
rect 24268 5856 24274 5908
rect 25225 5899 25283 5905
rect 25225 5865 25237 5899
rect 25271 5896 25283 5899
rect 25314 5896 25320 5908
rect 25271 5868 25320 5896
rect 25271 5865 25283 5868
rect 25225 5859 25283 5865
rect 25314 5856 25320 5868
rect 25372 5856 25378 5908
rect 13725 5831 13783 5837
rect 13725 5797 13737 5831
rect 13771 5797 13783 5831
rect 13725 5791 13783 5797
rect 13814 5788 13820 5840
rect 13872 5828 13878 5840
rect 13872 5800 13917 5828
rect 13872 5788 13878 5800
rect 15562 5788 15568 5840
rect 15620 5837 15626 5840
rect 15620 5831 15668 5837
rect 15620 5797 15622 5831
rect 15656 5797 15668 5831
rect 17218 5828 17224 5840
rect 17131 5800 17224 5828
rect 15620 5791 15668 5797
rect 15620 5788 15626 5791
rect 17218 5788 17224 5800
rect 17276 5788 17282 5840
rect 18966 5828 18972 5840
rect 18927 5800 18972 5828
rect 18966 5788 18972 5800
rect 19024 5788 19030 5840
rect 19061 5831 19119 5837
rect 19061 5797 19073 5831
rect 19107 5828 19119 5831
rect 19242 5828 19248 5840
rect 19107 5800 19248 5828
rect 19107 5797 19119 5800
rect 19061 5791 19119 5797
rect 19242 5788 19248 5800
rect 19300 5788 19306 5840
rect 20349 5831 20407 5837
rect 20349 5797 20361 5831
rect 20395 5828 20407 5831
rect 20438 5828 20444 5840
rect 20395 5800 20444 5828
rect 20395 5797 20407 5800
rect 20349 5791 20407 5797
rect 20438 5788 20444 5800
rect 20496 5828 20502 5840
rect 20496 5800 21404 5828
rect 20496 5788 20502 5800
rect 21376 5772 21404 5800
rect 22462 5788 22468 5840
rect 22520 5828 22526 5840
rect 22741 5831 22799 5837
rect 22741 5828 22753 5831
rect 22520 5800 22753 5828
rect 22520 5788 22526 5800
rect 22741 5797 22753 5800
rect 22787 5797 22799 5831
rect 22741 5791 22799 5797
rect 23293 5831 23351 5837
rect 23293 5797 23305 5831
rect 23339 5828 23351 5831
rect 23934 5828 23940 5840
rect 23339 5800 23940 5828
rect 23339 5797 23351 5800
rect 23293 5791 23351 5797
rect 23934 5788 23940 5800
rect 23992 5828 23998 5840
rect 24302 5828 24308 5840
rect 23992 5800 24308 5828
rect 23992 5788 23998 5800
rect 24302 5788 24308 5800
rect 24360 5788 24366 5840
rect 7742 5760 7748 5772
rect 7484 5732 7748 5760
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 10045 5763 10103 5769
rect 10045 5729 10057 5763
rect 10091 5760 10103 5763
rect 10321 5763 10379 5769
rect 10321 5760 10333 5763
rect 10091 5732 10333 5760
rect 10091 5729 10103 5732
rect 10045 5723 10103 5729
rect 10321 5729 10333 5732
rect 10367 5729 10379 5763
rect 12066 5760 12072 5772
rect 12027 5732 12072 5760
rect 10321 5723 10379 5729
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 12618 5760 12624 5772
rect 12579 5732 12624 5760
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 14734 5760 14740 5772
rect 14695 5732 14740 5760
rect 14734 5720 14740 5732
rect 14792 5720 14798 5772
rect 20530 5720 20536 5772
rect 20588 5760 20594 5772
rect 20898 5760 20904 5772
rect 20588 5732 20904 5760
rect 20588 5720 20594 5732
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 21358 5760 21364 5772
rect 21319 5732 21364 5760
rect 21358 5720 21364 5732
rect 21416 5720 21422 5772
rect 23842 5720 23848 5772
rect 23900 5760 23906 5772
rect 24121 5763 24179 5769
rect 24121 5760 24133 5763
rect 23900 5732 24133 5760
rect 23900 5720 23906 5732
rect 24121 5729 24133 5732
rect 24167 5729 24179 5763
rect 24121 5723 24179 5729
rect 2682 5652 2688 5704
rect 2740 5692 2746 5704
rect 2777 5695 2835 5701
rect 2777 5692 2789 5695
rect 2740 5664 2789 5692
rect 2740 5652 2746 5664
rect 2777 5661 2789 5664
rect 2823 5692 2835 5695
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 2823 5664 3801 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 3789 5661 3801 5664
rect 3835 5692 3847 5695
rect 3970 5692 3976 5704
rect 3835 5664 3976 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4341 5695 4399 5701
rect 4341 5692 4353 5695
rect 4120 5664 4353 5692
rect 4120 5652 4126 5664
rect 4341 5661 4353 5664
rect 4387 5692 4399 5695
rect 5537 5695 5595 5701
rect 5537 5692 5549 5695
rect 4387 5664 5549 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 5537 5661 5549 5664
rect 5583 5661 5595 5695
rect 5902 5692 5908 5704
rect 5863 5664 5908 5692
rect 5537 5655 5595 5661
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7009 5695 7067 5701
rect 7009 5692 7021 5695
rect 6972 5664 7021 5692
rect 6972 5652 6978 5664
rect 7009 5661 7021 5664
rect 7055 5692 7067 5695
rect 8202 5692 8208 5704
rect 7055 5664 8208 5692
rect 7055 5661 7067 5664
rect 7009 5655 7067 5661
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 9766 5652 9772 5704
rect 9824 5692 9830 5704
rect 10502 5692 10508 5704
rect 9824 5664 10508 5692
rect 9824 5652 9830 5664
rect 10502 5652 10508 5664
rect 10560 5692 10566 5704
rect 10689 5695 10747 5701
rect 10689 5692 10701 5695
rect 10560 5664 10701 5692
rect 10560 5652 10566 5664
rect 10689 5661 10701 5664
rect 10735 5661 10747 5695
rect 10689 5655 10747 5661
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5692 12863 5695
rect 14826 5692 14832 5704
rect 12851 5664 14832 5692
rect 12851 5661 12863 5664
rect 12805 5655 12863 5661
rect 14826 5652 14832 5664
rect 14884 5692 14890 5704
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 14884 5664 15301 5692
rect 14884 5652 14890 5664
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5661 17187 5695
rect 22646 5692 22652 5704
rect 22607 5664 22652 5692
rect 17129 5655 17187 5661
rect 2547 5627 2605 5633
rect 2547 5624 2559 5627
rect 2240 5596 2559 5624
rect 2240 5568 2268 5596
rect 2547 5593 2559 5596
rect 2593 5624 2605 5627
rect 2866 5624 2872 5636
rect 2593 5596 2872 5624
rect 2593 5593 2605 5596
rect 2547 5587 2605 5593
rect 2866 5584 2872 5596
rect 2924 5584 2930 5636
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 10597 5627 10655 5633
rect 10597 5624 10609 5627
rect 9732 5596 10609 5624
rect 9732 5584 9738 5596
rect 10597 5593 10609 5596
rect 10643 5593 10655 5627
rect 10597 5587 10655 5593
rect 14182 5584 14188 5636
rect 14240 5624 14246 5636
rect 14277 5627 14335 5633
rect 14277 5624 14289 5627
rect 14240 5596 14289 5624
rect 14240 5584 14246 5596
rect 14277 5593 14289 5596
rect 14323 5624 14335 5627
rect 17034 5624 17040 5636
rect 14323 5596 17040 5624
rect 14323 5593 14335 5596
rect 14277 5587 14335 5593
rect 17034 5584 17040 5596
rect 17092 5624 17098 5636
rect 17144 5624 17172 5655
rect 22646 5652 22652 5664
rect 22704 5652 22710 5704
rect 24136 5692 24164 5723
rect 24210 5720 24216 5772
rect 24268 5760 24274 5772
rect 24581 5763 24639 5769
rect 24581 5760 24593 5763
rect 24268 5732 24593 5760
rect 24268 5720 24274 5732
rect 24581 5729 24593 5732
rect 24627 5729 24639 5763
rect 24581 5723 24639 5729
rect 24670 5692 24676 5704
rect 24136 5664 24676 5692
rect 24670 5652 24676 5664
rect 24728 5652 24734 5704
rect 17092 5596 17172 5624
rect 17092 5584 17098 5596
rect 17310 5584 17316 5636
rect 17368 5624 17374 5636
rect 17681 5627 17739 5633
rect 17681 5624 17693 5627
rect 17368 5596 17693 5624
rect 17368 5584 17374 5596
rect 17681 5593 17693 5596
rect 17727 5624 17739 5627
rect 19150 5624 19156 5636
rect 17727 5596 19156 5624
rect 17727 5593 17739 5596
rect 17681 5587 17739 5593
rect 19150 5584 19156 5596
rect 19208 5624 19214 5636
rect 19518 5624 19524 5636
rect 19208 5596 19524 5624
rect 19208 5584 19214 5596
rect 19518 5584 19524 5596
rect 19576 5584 19582 5636
rect 2222 5556 2228 5568
rect 2183 5528 2228 5556
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 2682 5556 2688 5568
rect 2643 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 3326 5516 3332 5568
rect 3384 5556 3390 5568
rect 3421 5559 3479 5565
rect 3421 5556 3433 5559
rect 3384 5528 3433 5556
rect 3384 5516 3390 5528
rect 3421 5525 3433 5528
rect 3467 5525 3479 5559
rect 3421 5519 3479 5525
rect 3786 5516 3792 5568
rect 3844 5556 3850 5568
rect 4154 5556 4160 5568
rect 3844 5528 4160 5556
rect 3844 5516 3850 5528
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 9858 5516 9864 5568
rect 9916 5556 9922 5568
rect 10045 5559 10103 5565
rect 10045 5556 10057 5559
rect 9916 5528 10057 5556
rect 9916 5516 9922 5528
rect 10045 5525 10057 5528
rect 10091 5556 10103 5559
rect 10137 5559 10195 5565
rect 10137 5556 10149 5559
rect 10091 5528 10149 5556
rect 10091 5525 10103 5528
rect 10045 5519 10103 5525
rect 10137 5525 10149 5528
rect 10183 5525 10195 5559
rect 10137 5519 10195 5525
rect 10410 5516 10416 5568
rect 10468 5565 10474 5568
rect 10468 5559 10517 5565
rect 10468 5525 10471 5559
rect 10505 5556 10517 5559
rect 10778 5556 10784 5568
rect 10505 5528 10784 5556
rect 10505 5525 10517 5528
rect 10468 5519 10517 5525
rect 10468 5516 10474 5519
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 10870 5516 10876 5568
rect 10928 5556 10934 5568
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 10928 5528 11345 5556
rect 10928 5516 10934 5528
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 11333 5519 11391 5525
rect 17862 5516 17868 5568
rect 17920 5556 17926 5568
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 17920 5528 18061 5556
rect 17920 5516 17926 5528
rect 18049 5525 18061 5528
rect 18095 5525 18107 5559
rect 21910 5556 21916 5568
rect 21871 5528 21916 5556
rect 18049 5519 18107 5525
rect 21910 5516 21916 5528
rect 21968 5516 21974 5568
rect 22370 5556 22376 5568
rect 22283 5528 22376 5556
rect 22370 5516 22376 5528
rect 22428 5556 22434 5568
rect 23382 5556 23388 5568
rect 22428 5528 23388 5556
rect 22428 5516 22434 5528
rect 23382 5516 23388 5528
rect 23440 5516 23446 5568
rect 23753 5559 23811 5565
rect 23753 5525 23765 5559
rect 23799 5556 23811 5559
rect 24210 5556 24216 5568
rect 23799 5528 24216 5556
rect 23799 5525 23811 5528
rect 23753 5519 23811 5525
rect 24210 5516 24216 5528
rect 24268 5516 24274 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1838 5355 1896 5361
rect 1838 5321 1850 5355
rect 1884 5352 1896 5355
rect 2222 5352 2228 5364
rect 1884 5324 2228 5352
rect 1884 5321 1896 5324
rect 1838 5315 1896 5321
rect 2222 5312 2228 5324
rect 2280 5312 2286 5364
rect 2317 5355 2375 5361
rect 2317 5321 2329 5355
rect 2363 5352 2375 5355
rect 2406 5352 2412 5364
rect 2363 5324 2412 5352
rect 2363 5321 2375 5324
rect 2317 5315 2375 5321
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 4433 5355 4491 5361
rect 4433 5321 4445 5355
rect 4479 5352 4491 5355
rect 4522 5352 4528 5364
rect 4479 5324 4528 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 6273 5355 6331 5361
rect 6273 5321 6285 5355
rect 6319 5352 6331 5355
rect 6914 5352 6920 5364
rect 6319 5324 6920 5352
rect 6319 5321 6331 5324
rect 6273 5315 6331 5321
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 8386 5352 8392 5364
rect 8347 5324 8392 5352
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 10781 5355 10839 5361
rect 10781 5352 10793 5355
rect 9824 5324 10793 5352
rect 9824 5312 9830 5324
rect 10781 5321 10793 5324
rect 10827 5352 10839 5355
rect 10962 5352 10968 5364
rect 10827 5324 10968 5352
rect 10827 5321 10839 5324
rect 10781 5315 10839 5321
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11146 5352 11152 5364
rect 11107 5324 11152 5352
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 12066 5352 12072 5364
rect 12027 5324 12072 5352
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 12618 5312 12624 5364
rect 12676 5352 12682 5364
rect 12713 5355 12771 5361
rect 12713 5352 12725 5355
rect 12676 5324 12725 5352
rect 12676 5312 12682 5324
rect 12713 5321 12725 5324
rect 12759 5352 12771 5355
rect 13081 5355 13139 5361
rect 13081 5352 13093 5355
rect 12759 5324 13093 5352
rect 12759 5321 12771 5324
rect 12713 5315 12771 5321
rect 13081 5321 13093 5324
rect 13127 5352 13139 5355
rect 13998 5352 14004 5364
rect 13127 5324 14004 5352
rect 13127 5321 13139 5324
rect 13081 5315 13139 5321
rect 13998 5312 14004 5324
rect 14056 5312 14062 5364
rect 14642 5312 14648 5364
rect 14700 5352 14706 5364
rect 14829 5355 14887 5361
rect 14829 5352 14841 5355
rect 14700 5324 14841 5352
rect 14700 5312 14706 5324
rect 14829 5321 14841 5324
rect 14875 5321 14887 5355
rect 17218 5352 17224 5364
rect 17179 5324 17224 5352
rect 14829 5315 14887 5321
rect 17218 5312 17224 5324
rect 17276 5312 17282 5364
rect 19242 5312 19248 5364
rect 19300 5352 19306 5364
rect 19613 5355 19671 5361
rect 19613 5352 19625 5355
rect 19300 5324 19625 5352
rect 19300 5312 19306 5324
rect 19613 5321 19625 5324
rect 19659 5321 19671 5355
rect 19613 5315 19671 5321
rect 20717 5355 20775 5361
rect 20717 5321 20729 5355
rect 20763 5352 20775 5355
rect 21266 5352 21272 5364
rect 20763 5324 21272 5352
rect 20763 5321 20775 5324
rect 20717 5315 20775 5321
rect 1949 5287 2007 5293
rect 1949 5253 1961 5287
rect 1995 5284 2007 5287
rect 2130 5284 2136 5296
rect 1995 5256 2136 5284
rect 1995 5253 2007 5256
rect 1949 5247 2007 5253
rect 2130 5244 2136 5256
rect 2188 5284 2194 5296
rect 2774 5284 2780 5296
rect 2188 5256 2780 5284
rect 2188 5244 2194 5256
rect 2774 5244 2780 5256
rect 2832 5284 2838 5296
rect 3053 5287 3111 5293
rect 3053 5284 3065 5287
rect 2832 5256 3065 5284
rect 2832 5244 2838 5256
rect 3053 5253 3065 5256
rect 3099 5253 3111 5287
rect 10134 5284 10140 5296
rect 3053 5247 3111 5253
rect 3896 5256 10140 5284
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2314 5216 2320 5228
rect 2087 5188 2320 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2314 5176 2320 5188
rect 2372 5216 2378 5228
rect 2869 5219 2927 5225
rect 2869 5216 2881 5219
rect 2372 5188 2881 5216
rect 2372 5176 2378 5188
rect 2869 5185 2881 5188
rect 2915 5185 2927 5219
rect 2869 5179 2927 5185
rect 2958 5176 2964 5228
rect 3016 5216 3022 5228
rect 3896 5216 3924 5256
rect 10134 5244 10140 5256
rect 10192 5284 10198 5296
rect 10410 5284 10416 5296
rect 10192 5256 10416 5284
rect 10192 5244 10198 5256
rect 10410 5244 10416 5256
rect 10468 5284 10474 5296
rect 10643 5287 10701 5293
rect 10643 5284 10655 5287
rect 10468 5256 10655 5284
rect 10468 5244 10474 5256
rect 10643 5253 10655 5256
rect 10689 5253 10701 5287
rect 19334 5284 19340 5296
rect 19295 5256 19340 5284
rect 10643 5247 10701 5253
rect 19334 5244 19340 5256
rect 19392 5244 19398 5296
rect 3016 5188 3924 5216
rect 3973 5219 4031 5225
rect 3016 5176 3022 5188
rect 3973 5185 3985 5219
rect 4019 5216 4031 5219
rect 4062 5216 4068 5228
rect 4019 5188 4068 5216
rect 4019 5185 4031 5188
rect 3973 5179 4031 5185
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4890 5216 4896 5228
rect 4851 5188 4896 5216
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 6822 5216 6828 5228
rect 6783 5188 6828 5216
rect 6822 5176 6828 5188
rect 6880 5176 6886 5228
rect 10229 5219 10287 5225
rect 10229 5185 10241 5219
rect 10275 5216 10287 5219
rect 10502 5216 10508 5228
rect 10275 5188 10508 5216
rect 10275 5185 10287 5188
rect 10229 5179 10287 5185
rect 10502 5176 10508 5188
rect 10560 5216 10566 5228
rect 10873 5219 10931 5225
rect 10873 5216 10885 5219
rect 10560 5188 10885 5216
rect 10560 5176 10566 5188
rect 10873 5185 10885 5188
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 13909 5219 13967 5225
rect 13909 5185 13921 5219
rect 13955 5216 13967 5219
rect 14734 5216 14740 5228
rect 13955 5188 14740 5216
rect 13955 5185 13967 5188
rect 13909 5179 13967 5185
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 15654 5216 15660 5228
rect 15615 5188 15660 5216
rect 15654 5176 15660 5188
rect 15712 5216 15718 5228
rect 16853 5219 16911 5225
rect 16853 5216 16865 5219
rect 15712 5188 16865 5216
rect 15712 5176 15718 5188
rect 16853 5185 16865 5188
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 2130 5108 2136 5160
rect 2188 5148 2194 5160
rect 3513 5151 3571 5157
rect 3513 5148 3525 5151
rect 2188 5120 3525 5148
rect 2188 5108 2194 5120
rect 3513 5117 3525 5120
rect 3559 5117 3571 5151
rect 3513 5111 3571 5117
rect 3789 5151 3847 5157
rect 3789 5117 3801 5151
rect 3835 5148 3847 5151
rect 4706 5148 4712 5160
rect 3835 5120 4712 5148
rect 3835 5117 3847 5120
rect 3789 5111 3847 5117
rect 1673 5083 1731 5089
rect 1673 5049 1685 5083
rect 1719 5080 1731 5083
rect 2498 5080 2504 5092
rect 1719 5052 2504 5080
rect 1719 5049 1731 5052
rect 1673 5043 1731 5049
rect 2498 5040 2504 5052
rect 2556 5040 2562 5092
rect 2777 5083 2835 5089
rect 2777 5049 2789 5083
rect 2823 5080 2835 5083
rect 2866 5080 2872 5092
rect 2823 5052 2872 5080
rect 2823 5049 2835 5052
rect 2777 5043 2835 5049
rect 2866 5040 2872 5052
rect 2924 5040 2930 5092
rect 3528 5080 3556 5111
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 6641 5151 6699 5157
rect 6641 5148 6653 5151
rect 6052 5120 6653 5148
rect 6052 5108 6058 5120
rect 6641 5117 6653 5120
rect 6687 5148 6699 5151
rect 6914 5148 6920 5160
rect 6687 5120 6920 5148
rect 6687 5117 6699 5120
rect 6641 5111 6699 5117
rect 6914 5108 6920 5120
rect 6972 5148 6978 5160
rect 7742 5148 7748 5160
rect 6972 5120 7748 5148
rect 6972 5108 6978 5120
rect 3878 5080 3884 5092
rect 3528 5052 3884 5080
rect 3878 5040 3884 5052
rect 3936 5040 3942 5092
rect 4985 5083 5043 5089
rect 4985 5049 4997 5083
rect 5031 5080 5043 5083
rect 5166 5080 5172 5092
rect 5031 5052 5172 5080
rect 5031 5049 5043 5052
rect 4985 5043 5043 5049
rect 5166 5040 5172 5052
rect 5224 5040 5230 5092
rect 5537 5083 5595 5089
rect 5537 5049 5549 5083
rect 5583 5080 5595 5083
rect 5626 5080 5632 5092
rect 5583 5052 5632 5080
rect 5583 5049 5595 5052
rect 5537 5043 5595 5049
rect 5626 5040 5632 5052
rect 5684 5040 5690 5092
rect 7202 5089 7230 5120
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 8386 5108 8392 5160
rect 8444 5148 8450 5160
rect 8573 5151 8631 5157
rect 8573 5148 8585 5151
rect 8444 5120 8585 5148
rect 8444 5108 8450 5120
rect 8573 5117 8585 5120
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 8662 5108 8668 5160
rect 8720 5148 8726 5160
rect 9033 5151 9091 5157
rect 9033 5148 9045 5151
rect 8720 5120 9045 5148
rect 8720 5108 8726 5120
rect 9033 5117 9045 5120
rect 9079 5117 9091 5151
rect 9033 5111 9091 5117
rect 12526 5108 12532 5160
rect 12584 5148 12590 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12584 5120 12909 5148
rect 12584 5108 12590 5120
rect 12897 5117 12909 5120
rect 12943 5148 12955 5151
rect 13357 5151 13415 5157
rect 13357 5148 13369 5151
rect 12943 5120 13369 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 13357 5117 13369 5120
rect 13403 5117 13415 5151
rect 13357 5111 13415 5117
rect 18969 5151 19027 5157
rect 18969 5117 18981 5151
rect 19015 5148 19027 5151
rect 19242 5148 19248 5160
rect 19015 5120 19248 5148
rect 19015 5117 19027 5120
rect 18969 5111 19027 5117
rect 19242 5108 19248 5120
rect 19300 5108 19306 5160
rect 20073 5151 20131 5157
rect 20073 5117 20085 5151
rect 20119 5148 20131 5151
rect 20732 5148 20760 5315
rect 21266 5312 21272 5324
rect 21324 5312 21330 5364
rect 22646 5312 22652 5364
rect 22704 5352 22710 5364
rect 22741 5355 22799 5361
rect 22741 5352 22753 5355
rect 22704 5324 22753 5352
rect 22704 5312 22710 5324
rect 22741 5321 22753 5324
rect 22787 5321 22799 5355
rect 22741 5315 22799 5321
rect 23290 5312 23296 5364
rect 23348 5352 23354 5364
rect 23385 5355 23443 5361
rect 23385 5352 23397 5355
rect 23348 5324 23397 5352
rect 23348 5312 23354 5324
rect 23385 5321 23397 5324
rect 23431 5321 23443 5355
rect 24670 5352 24676 5364
rect 24631 5324 24676 5352
rect 23385 5315 23443 5321
rect 21177 5219 21235 5225
rect 21177 5185 21189 5219
rect 21223 5216 21235 5219
rect 21910 5216 21916 5228
rect 21223 5188 21916 5216
rect 21223 5185 21235 5188
rect 21177 5179 21235 5185
rect 21910 5176 21916 5188
rect 21968 5176 21974 5228
rect 20119 5120 20760 5148
rect 23400 5148 23428 5315
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 23661 5151 23719 5157
rect 23661 5148 23673 5151
rect 23400 5120 23673 5148
rect 20119 5117 20131 5120
rect 20073 5111 20131 5117
rect 23661 5117 23673 5120
rect 23707 5117 23719 5151
rect 24210 5148 24216 5160
rect 24171 5120 24216 5148
rect 23661 5111 23719 5117
rect 24210 5108 24216 5120
rect 24268 5108 24274 5160
rect 25222 5148 25228 5160
rect 25183 5120 25228 5148
rect 25222 5108 25228 5120
rect 25280 5148 25286 5160
rect 25777 5151 25835 5157
rect 25777 5148 25789 5151
rect 25280 5120 25789 5148
rect 25280 5108 25286 5120
rect 25777 5117 25789 5120
rect 25823 5117 25835 5151
rect 25777 5111 25835 5117
rect 7187 5083 7245 5089
rect 7187 5049 7199 5083
rect 7233 5049 7245 5083
rect 7187 5043 7245 5049
rect 7466 5040 7472 5092
rect 7524 5080 7530 5092
rect 8018 5080 8024 5092
rect 7524 5052 8024 5080
rect 7524 5040 7530 5052
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 8202 5040 8208 5092
rect 8260 5080 8266 5092
rect 8260 5052 8708 5080
rect 8260 5040 8266 5052
rect 5184 5012 5212 5040
rect 5813 5015 5871 5021
rect 5813 5012 5825 5015
rect 5184 4984 5825 5012
rect 5813 4981 5825 4984
rect 5859 4981 5871 5015
rect 7742 5012 7748 5024
rect 7703 4984 7748 5012
rect 5813 4975 5871 4981
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 8680 5021 8708 5052
rect 10042 5040 10048 5092
rect 10100 5080 10106 5092
rect 10505 5083 10563 5089
rect 10505 5080 10517 5083
rect 10100 5052 10517 5080
rect 10100 5040 10106 5052
rect 10505 5049 10517 5052
rect 10551 5080 10563 5083
rect 10870 5080 10876 5092
rect 10551 5052 10876 5080
rect 10551 5049 10563 5052
rect 10505 5043 10563 5049
rect 10870 5040 10876 5052
rect 10928 5040 10934 5092
rect 14271 5083 14329 5089
rect 14271 5049 14283 5083
rect 14317 5080 14329 5083
rect 15978 5083 16036 5089
rect 14317 5052 14351 5080
rect 14317 5049 14329 5052
rect 14271 5043 14329 5049
rect 15978 5049 15990 5083
rect 16024 5049 16036 5083
rect 18322 5080 18328 5092
rect 18283 5052 18328 5080
rect 15978 5043 16036 5049
rect 8665 5015 8723 5021
rect 8665 4981 8677 5015
rect 8711 4981 8723 5015
rect 9674 5012 9680 5024
rect 9635 4984 9680 5012
rect 8665 4975 8723 4981
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 9950 5012 9956 5024
rect 9911 4984 9956 5012
rect 9950 4972 9956 4984
rect 10008 5012 10014 5024
rect 10229 5015 10287 5021
rect 10229 5012 10241 5015
rect 10008 4984 10241 5012
rect 10008 4972 10014 4984
rect 10229 4981 10241 4984
rect 10275 5012 10287 5015
rect 10321 5015 10379 5021
rect 10321 5012 10333 5015
rect 10275 4984 10333 5012
rect 10275 4981 10287 4984
rect 10229 4975 10287 4981
rect 10321 4981 10333 4984
rect 10367 4981 10379 5015
rect 10321 4975 10379 4981
rect 10778 4972 10784 5024
rect 10836 5012 10842 5024
rect 11422 5012 11428 5024
rect 10836 4984 11428 5012
rect 10836 4972 10842 4984
rect 11422 4972 11428 4984
rect 11480 5012 11486 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 11480 4984 11529 5012
rect 11480 4972 11486 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 11517 4975 11575 4981
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 13817 5015 13875 5021
rect 13817 5012 13829 5015
rect 11756 4984 13829 5012
rect 11756 4972 11762 4984
rect 13817 4981 13829 4984
rect 13863 5012 13875 5015
rect 14286 5012 14314 5043
rect 15289 5015 15347 5021
rect 15289 5012 15301 5015
rect 13863 4984 15301 5012
rect 13863 4981 13875 4984
rect 13817 4975 13875 4981
rect 15289 4981 15301 4984
rect 15335 5012 15347 5015
rect 15654 5012 15660 5024
rect 15335 4984 15660 5012
rect 15335 4981 15347 4984
rect 15289 4975 15347 4981
rect 15654 4972 15660 4984
rect 15712 5012 15718 5024
rect 15993 5012 16021 5043
rect 18322 5040 18328 5052
rect 18380 5040 18386 5092
rect 18414 5040 18420 5092
rect 18472 5089 18478 5092
rect 18472 5080 18484 5089
rect 21498 5083 21556 5089
rect 21498 5080 21510 5083
rect 18472 5052 18517 5080
rect 21100 5052 21510 5080
rect 18472 5043 18484 5052
rect 18472 5040 18478 5043
rect 21100 5024 21128 5052
rect 21498 5049 21510 5052
rect 21544 5049 21556 5083
rect 22370 5080 22376 5092
rect 22331 5052 22376 5080
rect 21498 5043 21556 5049
rect 22370 5040 22376 5052
rect 22428 5040 22434 5092
rect 16574 5012 16580 5024
rect 15712 4984 16021 5012
rect 16535 4984 16580 5012
rect 15712 4972 15718 4984
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 17494 4972 17500 5024
rect 17552 5012 17558 5024
rect 17773 5015 17831 5021
rect 17773 5012 17785 5015
rect 17552 4984 17785 5012
rect 17552 4972 17558 4984
rect 17773 4981 17785 4984
rect 17819 4981 17831 5015
rect 20254 5012 20260 5024
rect 20215 4984 20260 5012
rect 17773 4975 17831 4981
rect 20254 4972 20260 4984
rect 20312 4972 20318 5024
rect 21082 5012 21088 5024
rect 21043 4984 21088 5012
rect 21082 4972 21088 4984
rect 21140 4972 21146 5024
rect 22094 4972 22100 5024
rect 22152 5012 22158 5024
rect 22152 4984 22197 5012
rect 22152 4972 22158 4984
rect 23474 4972 23480 5024
rect 23532 5012 23538 5024
rect 23753 5015 23811 5021
rect 23753 5012 23765 5015
rect 23532 4984 23765 5012
rect 23532 4972 23538 4984
rect 23753 4981 23765 4984
rect 23799 4981 23811 5015
rect 23753 4975 23811 4981
rect 25409 5015 25467 5021
rect 25409 4981 25421 5015
rect 25455 5012 25467 5015
rect 25498 5012 25504 5024
rect 25455 4984 25504 5012
rect 25455 4981 25467 4984
rect 25409 4975 25467 4981
rect 25498 4972 25504 4984
rect 25556 4972 25562 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1535 4811 1593 4817
rect 1535 4777 1547 4811
rect 1581 4808 1593 4811
rect 1854 4808 1860 4820
rect 1581 4780 1860 4808
rect 1581 4777 1593 4780
rect 1535 4771 1593 4777
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 2317 4811 2375 4817
rect 2317 4777 2329 4811
rect 2363 4808 2375 4811
rect 2774 4808 2780 4820
rect 2363 4780 2780 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 2774 4768 2780 4780
rect 2832 4768 2838 4820
rect 2958 4768 2964 4820
rect 3016 4808 3022 4820
rect 3421 4811 3479 4817
rect 3421 4808 3433 4811
rect 3016 4780 3433 4808
rect 3016 4768 3022 4780
rect 3421 4777 3433 4780
rect 3467 4777 3479 4811
rect 3878 4808 3884 4820
rect 3839 4780 3884 4808
rect 3421 4771 3479 4777
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 4212 4780 4261 4808
rect 4212 4768 4218 4780
rect 4249 4777 4261 4780
rect 4295 4777 4307 4811
rect 4706 4808 4712 4820
rect 4667 4780 4712 4808
rect 4249 4771 4307 4777
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 6914 4808 6920 4820
rect 6875 4780 6920 4808
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 7300 4780 8217 4808
rect 7300 4752 7328 4780
rect 8205 4777 8217 4780
rect 8251 4777 8263 4811
rect 8570 4808 8576 4820
rect 8531 4780 8576 4808
rect 8205 4771 8263 4777
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 9030 4808 9036 4820
rect 8991 4780 9036 4808
rect 9030 4768 9036 4780
rect 9088 4768 9094 4820
rect 10778 4808 10784 4820
rect 10739 4780 10784 4808
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 10962 4768 10968 4820
rect 11020 4808 11026 4820
rect 11057 4811 11115 4817
rect 11057 4808 11069 4811
rect 11020 4780 11069 4808
rect 11020 4768 11026 4780
rect 11057 4777 11069 4780
rect 11103 4777 11115 4811
rect 11330 4808 11336 4820
rect 11291 4780 11336 4808
rect 11057 4771 11115 4777
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14461 4811 14519 4817
rect 14461 4808 14473 4811
rect 13872 4780 14473 4808
rect 13872 4768 13878 4780
rect 14461 4777 14473 4780
rect 14507 4777 14519 4811
rect 14461 4771 14519 4777
rect 14826 4768 14832 4820
rect 14884 4808 14890 4820
rect 15013 4811 15071 4817
rect 15013 4808 15025 4811
rect 14884 4780 15025 4808
rect 14884 4768 14890 4780
rect 15013 4777 15025 4780
rect 15059 4777 15071 4811
rect 15013 4771 15071 4777
rect 17497 4811 17555 4817
rect 17497 4777 17509 4811
rect 17543 4808 17555 4811
rect 17586 4808 17592 4820
rect 17543 4780 17592 4808
rect 17543 4777 17555 4780
rect 17497 4771 17555 4777
rect 17586 4768 17592 4780
rect 17644 4768 17650 4820
rect 18141 4811 18199 4817
rect 18141 4777 18153 4811
rect 18187 4808 18199 4811
rect 18230 4808 18236 4820
rect 18187 4780 18236 4808
rect 18187 4777 18199 4780
rect 18141 4771 18199 4777
rect 18230 4768 18236 4780
rect 18288 4768 18294 4820
rect 18322 4768 18328 4820
rect 18380 4808 18386 4820
rect 19337 4811 19395 4817
rect 19337 4808 19349 4811
rect 18380 4780 19349 4808
rect 18380 4768 18386 4780
rect 19337 4777 19349 4780
rect 19383 4808 19395 4811
rect 20346 4808 20352 4820
rect 19383 4780 20352 4808
rect 19383 4777 19395 4780
rect 19337 4771 19395 4777
rect 20346 4768 20352 4780
rect 20404 4768 20410 4820
rect 22462 4768 22468 4820
rect 22520 4808 22526 4820
rect 22557 4811 22615 4817
rect 22557 4808 22569 4811
rect 22520 4780 22569 4808
rect 22520 4768 22526 4780
rect 22557 4777 22569 4780
rect 22603 4777 22615 4811
rect 22557 4771 22615 4777
rect 1118 4700 1124 4752
rect 1176 4740 1182 4752
rect 1949 4743 2007 4749
rect 1949 4740 1961 4743
rect 1176 4712 1961 4740
rect 1176 4700 1182 4712
rect 1949 4709 1961 4712
rect 1995 4709 2007 4743
rect 1949 4703 2007 4709
rect 3145 4743 3203 4749
rect 3145 4709 3157 4743
rect 3191 4740 3203 4743
rect 3234 4740 3240 4752
rect 3191 4712 3240 4740
rect 3191 4709 3203 4712
rect 3145 4703 3203 4709
rect 3234 4700 3240 4712
rect 3292 4700 3298 4752
rect 5074 4740 5080 4752
rect 5035 4712 5080 4740
rect 5074 4700 5080 4712
rect 5132 4700 5138 4752
rect 5626 4740 5632 4752
rect 5587 4712 5632 4740
rect 5626 4700 5632 4712
rect 5684 4740 5690 4752
rect 7282 4740 7288 4752
rect 5684 4712 7288 4740
rect 5684 4700 5690 4712
rect 7282 4700 7288 4712
rect 7340 4700 7346 4752
rect 7377 4743 7435 4749
rect 7377 4709 7389 4743
rect 7423 4740 7435 4743
rect 7742 4740 7748 4752
rect 7423 4712 7748 4740
rect 7423 4709 7435 4712
rect 7377 4703 7435 4709
rect 7742 4700 7748 4712
rect 7800 4700 7806 4752
rect 9048 4740 9076 4768
rect 9677 4743 9735 4749
rect 9677 4740 9689 4743
rect 9048 4712 9689 4740
rect 9677 4709 9689 4712
rect 9723 4740 9735 4743
rect 9858 4740 9864 4752
rect 9723 4712 9864 4740
rect 9723 4709 9735 4712
rect 9677 4703 9735 4709
rect 9858 4700 9864 4712
rect 9916 4700 9922 4752
rect 10413 4743 10471 4749
rect 10413 4709 10425 4743
rect 10459 4740 10471 4743
rect 10686 4740 10692 4752
rect 10459 4712 10692 4740
rect 10459 4709 10471 4712
rect 10413 4703 10471 4709
rect 10686 4700 10692 4712
rect 10744 4700 10750 4752
rect 13630 4740 13636 4752
rect 13591 4712 13636 4740
rect 13630 4700 13636 4712
rect 13688 4700 13694 4752
rect 14182 4740 14188 4752
rect 14143 4712 14188 4740
rect 14182 4700 14188 4712
rect 14240 4700 14246 4752
rect 16114 4700 16120 4752
rect 16172 4740 16178 4752
rect 16209 4743 16267 4749
rect 16209 4740 16221 4743
rect 16172 4712 16221 4740
rect 16172 4700 16178 4712
rect 16209 4709 16221 4712
rect 16255 4740 16267 4743
rect 16574 4740 16580 4752
rect 16255 4712 16580 4740
rect 16255 4709 16267 4712
rect 16209 4703 16267 4709
rect 16574 4700 16580 4712
rect 16632 4700 16638 4752
rect 16761 4743 16819 4749
rect 16761 4709 16773 4743
rect 16807 4740 16819 4743
rect 17310 4740 17316 4752
rect 16807 4712 17316 4740
rect 16807 4709 16819 4712
rect 16761 4703 16819 4709
rect 17310 4700 17316 4712
rect 17368 4700 17374 4752
rect 18414 4740 18420 4752
rect 17512 4712 18420 4740
rect 17512 4684 17540 4712
rect 18414 4700 18420 4712
rect 18472 4700 18478 4752
rect 21082 4700 21088 4752
rect 21140 4740 21146 4752
rect 21406 4743 21464 4749
rect 21406 4740 21418 4743
rect 21140 4712 21418 4740
rect 21140 4700 21146 4712
rect 21406 4709 21418 4712
rect 21452 4709 21464 4743
rect 21406 4703 21464 4709
rect 22094 4700 22100 4752
rect 22152 4740 22158 4752
rect 22646 4740 22652 4752
rect 22152 4712 22652 4740
rect 22152 4700 22158 4712
rect 22646 4700 22652 4712
rect 22704 4740 22710 4752
rect 23017 4743 23075 4749
rect 23017 4740 23029 4743
rect 22704 4712 23029 4740
rect 22704 4700 22710 4712
rect 23017 4709 23029 4712
rect 23063 4709 23075 4743
rect 23017 4703 23075 4709
rect 23382 4700 23388 4752
rect 23440 4740 23446 4752
rect 23569 4743 23627 4749
rect 23569 4740 23581 4743
rect 23440 4712 23581 4740
rect 23440 4700 23446 4712
rect 23569 4709 23581 4712
rect 23615 4740 23627 4743
rect 23934 4740 23940 4752
rect 23615 4712 23940 4740
rect 23615 4709 23627 4712
rect 23569 4703 23627 4709
rect 23934 4700 23940 4712
rect 23992 4700 23998 4752
rect 24210 4700 24216 4752
rect 24268 4740 24274 4752
rect 24268 4712 24900 4740
rect 24268 4700 24274 4712
rect 1464 4675 1522 4681
rect 1464 4641 1476 4675
rect 1510 4672 1522 4675
rect 2222 4672 2228 4684
rect 1510 4644 2228 4672
rect 1510 4641 1522 4644
rect 1464 4635 1522 4641
rect 2222 4632 2228 4644
rect 2280 4632 2286 4684
rect 2409 4675 2467 4681
rect 2409 4641 2421 4675
rect 2455 4672 2467 4675
rect 2498 4672 2504 4684
rect 2455 4644 2504 4672
rect 2455 4641 2467 4644
rect 2409 4635 2467 4641
rect 2498 4632 2504 4644
rect 2556 4672 2562 4684
rect 3326 4672 3332 4684
rect 2556 4644 3332 4672
rect 2556 4632 2562 4644
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 6549 4675 6607 4681
rect 6549 4641 6561 4675
rect 6595 4672 6607 4675
rect 6730 4672 6736 4684
rect 6595 4644 6736 4672
rect 6595 4641 6607 4644
rect 6549 4635 6607 4641
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 9398 4672 9404 4684
rect 9359 4644 9404 4672
rect 9398 4632 9404 4644
rect 9456 4632 9462 4684
rect 11514 4672 11520 4684
rect 11475 4644 11520 4672
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 11793 4675 11851 4681
rect 11793 4641 11805 4675
rect 11839 4672 11851 4675
rect 12158 4672 12164 4684
rect 11839 4644 12164 4672
rect 11839 4641 11851 4644
rect 11793 4635 11851 4641
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 17494 4632 17500 4684
rect 17552 4632 17558 4684
rect 19702 4632 19708 4684
rect 19760 4672 19766 4684
rect 19864 4675 19922 4681
rect 19864 4672 19876 4675
rect 19760 4644 19876 4672
rect 19760 4632 19766 4644
rect 19864 4641 19876 4644
rect 19910 4672 19922 4675
rect 20622 4672 20628 4684
rect 19910 4644 20628 4672
rect 19910 4641 19922 4644
rect 19864 4635 19922 4641
rect 20622 4632 20628 4644
rect 20680 4632 20686 4684
rect 24673 4675 24731 4681
rect 24673 4641 24685 4675
rect 24719 4672 24731 4675
rect 24762 4672 24768 4684
rect 24719 4644 24768 4672
rect 24719 4641 24731 4644
rect 24673 4635 24731 4641
rect 24762 4632 24768 4644
rect 24820 4632 24826 4684
rect 24872 4681 24900 4712
rect 24857 4675 24915 4681
rect 24857 4641 24869 4675
rect 24903 4641 24915 4675
rect 24857 4635 24915 4641
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4604 2835 4607
rect 2866 4604 2872 4616
rect 2823 4576 2872 4604
rect 2823 4573 2835 4576
rect 2777 4567 2835 4573
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 4430 4564 4436 4616
rect 4488 4604 4494 4616
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 4488 4576 4997 4604
rect 4488 4564 4494 4576
rect 4985 4573 4997 4576
rect 5031 4604 5043 4607
rect 5905 4607 5963 4613
rect 5905 4604 5917 4607
rect 5031 4576 5917 4604
rect 5031 4573 5043 4576
rect 4985 4567 5043 4573
rect 5905 4573 5917 4576
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 7466 4564 7472 4616
rect 7524 4604 7530 4616
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7524 4576 7573 4604
rect 7524 4564 7530 4576
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 9416 4604 9444 4632
rect 10045 4607 10103 4613
rect 10045 4604 10057 4607
rect 9416 4576 10057 4604
rect 7561 4567 7619 4573
rect 10045 4573 10057 4576
rect 10091 4573 10103 4607
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 10045 4567 10103 4573
rect 13280 4576 13553 4604
rect 2682 4536 2688 4548
rect 2643 4508 2688 4536
rect 2682 4496 2688 4508
rect 2740 4496 2746 4548
rect 9842 4539 9900 4545
rect 9842 4505 9854 4539
rect 9888 4536 9900 4539
rect 10778 4536 10784 4548
rect 9888 4508 10784 4536
rect 9888 4505 9900 4508
rect 9842 4499 9900 4505
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 13280 4480 13308 4576
rect 13541 4573 13553 4576
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4604 16175 4607
rect 16206 4604 16212 4616
rect 16163 4576 16212 4604
rect 16163 4573 16175 4576
rect 16117 4567 16175 4573
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 18322 4604 18328 4616
rect 18283 4576 18328 4604
rect 18322 4564 18328 4576
rect 18380 4564 18386 4616
rect 18966 4604 18972 4616
rect 18927 4576 18972 4604
rect 18966 4564 18972 4576
rect 19024 4564 19030 4616
rect 21085 4607 21143 4613
rect 21085 4573 21097 4607
rect 21131 4604 21143 4607
rect 21174 4604 21180 4616
rect 21131 4576 21180 4604
rect 21131 4573 21143 4576
rect 21085 4567 21143 4573
rect 21174 4564 21180 4576
rect 21232 4564 21238 4616
rect 22925 4607 22983 4613
rect 22925 4573 22937 4607
rect 22971 4604 22983 4607
rect 23014 4604 23020 4616
rect 22971 4576 23020 4604
rect 22971 4573 22983 4576
rect 22925 4567 22983 4573
rect 23014 4564 23020 4576
rect 23072 4564 23078 4616
rect 24946 4604 24952 4616
rect 24907 4576 24952 4604
rect 24946 4564 24952 4576
rect 25004 4564 25010 4616
rect 20717 4539 20775 4545
rect 20717 4505 20729 4539
rect 20763 4536 20775 4539
rect 21358 4536 21364 4548
rect 20763 4508 21364 4536
rect 20763 4505 20775 4508
rect 20717 4499 20775 4505
rect 21358 4496 21364 4508
rect 21416 4536 21422 4548
rect 22186 4536 22192 4548
rect 21416 4508 22192 4536
rect 21416 4496 21422 4508
rect 22186 4496 22192 4508
rect 22244 4496 22250 4548
rect 2590 4477 2596 4480
rect 2574 4471 2596 4477
rect 2574 4437 2586 4471
rect 2574 4431 2596 4437
rect 2590 4428 2596 4431
rect 2648 4428 2654 4480
rect 3326 4428 3332 4480
rect 3384 4468 3390 4480
rect 8938 4468 8944 4480
rect 3384 4440 8944 4468
rect 3384 4428 3390 4440
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 9953 4471 10011 4477
rect 9953 4468 9965 4471
rect 9732 4440 9965 4468
rect 9732 4428 9738 4440
rect 9953 4437 9965 4440
rect 9999 4437 10011 4471
rect 9953 4431 10011 4437
rect 11146 4428 11152 4480
rect 11204 4468 11210 4480
rect 12253 4471 12311 4477
rect 12253 4468 12265 4471
rect 11204 4440 12265 4468
rect 11204 4428 11210 4440
rect 12253 4437 12265 4440
rect 12299 4437 12311 4471
rect 13262 4468 13268 4480
rect 13223 4440 13268 4468
rect 12253 4431 12311 4437
rect 13262 4428 13268 4440
rect 13320 4428 13326 4480
rect 15654 4468 15660 4480
rect 15615 4440 15660 4468
rect 15654 4428 15660 4440
rect 15712 4428 15718 4480
rect 17034 4468 17040 4480
rect 16995 4440 17040 4468
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 19334 4428 19340 4480
rect 19392 4468 19398 4480
rect 19935 4471 19993 4477
rect 19935 4468 19947 4471
rect 19392 4440 19947 4468
rect 19392 4428 19398 4440
rect 19935 4437 19947 4440
rect 19981 4437 19993 4471
rect 22002 4468 22008 4480
rect 21963 4440 22008 4468
rect 19935 4431 19993 4437
rect 22002 4428 22008 4440
rect 22060 4428 22066 4480
rect 24210 4468 24216 4480
rect 24171 4440 24216 4468
rect 24210 4428 24216 4440
rect 24268 4428 24274 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1946 4264 1952 4276
rect 1907 4236 1952 4264
rect 1946 4224 1952 4236
rect 2004 4224 2010 4276
rect 2866 4264 2872 4276
rect 2827 4236 2872 4264
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 3326 4264 3332 4276
rect 3287 4236 3332 4264
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 5350 4224 5356 4276
rect 5408 4264 5414 4276
rect 7653 4267 7711 4273
rect 7653 4264 7665 4267
rect 5408 4236 7665 4264
rect 5408 4224 5414 4236
rect 7653 4233 7665 4236
rect 7699 4233 7711 4267
rect 7653 4227 7711 4233
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 7837 4267 7895 4273
rect 7837 4264 7849 4267
rect 7800 4236 7849 4264
rect 7800 4224 7806 4236
rect 7837 4233 7849 4236
rect 7883 4233 7895 4267
rect 9674 4264 9680 4276
rect 9635 4236 9680 4264
rect 7837 4227 7895 4233
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 10042 4264 10048 4276
rect 10003 4236 10048 4264
rect 10042 4224 10048 4236
rect 10100 4224 10106 4276
rect 10778 4264 10784 4276
rect 10739 4236 10784 4264
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 11241 4267 11299 4273
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 11514 4264 11520 4276
rect 11287 4236 11520 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11514 4224 11520 4236
rect 11572 4224 11578 4276
rect 12158 4264 12164 4276
rect 12119 4236 12164 4264
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 16114 4264 16120 4276
rect 16075 4236 16120 4264
rect 16114 4224 16120 4236
rect 16172 4224 16178 4276
rect 17494 4264 17500 4276
rect 17455 4236 17500 4264
rect 17494 4224 17500 4236
rect 17552 4224 17558 4276
rect 18414 4224 18420 4276
rect 18472 4264 18478 4276
rect 18969 4267 19027 4273
rect 18969 4264 18981 4267
rect 18472 4236 18981 4264
rect 18472 4224 18478 4236
rect 18969 4233 18981 4236
rect 19015 4233 19027 4267
rect 19702 4264 19708 4276
rect 19663 4236 19708 4264
rect 18969 4227 19027 4233
rect 19702 4224 19708 4236
rect 19760 4224 19766 4276
rect 21821 4267 21879 4273
rect 21821 4233 21833 4267
rect 21867 4264 21879 4267
rect 22002 4264 22008 4276
rect 21867 4236 22008 4264
rect 21867 4233 21879 4236
rect 21821 4227 21879 4233
rect 22002 4224 22008 4236
rect 22060 4224 22066 4276
rect 24762 4264 24768 4276
rect 24723 4236 24768 4264
rect 24762 4224 24768 4236
rect 24820 4224 24826 4276
rect 6730 4156 6736 4208
rect 6788 4196 6794 4208
rect 6788 4168 6868 4196
rect 6788 4156 6794 4168
rect 5074 4088 5080 4140
rect 5132 4128 5138 4140
rect 5997 4131 6055 4137
rect 5997 4128 6009 4131
rect 5132 4100 6009 4128
rect 5132 4088 5138 4100
rect 5997 4097 6009 4100
rect 6043 4097 6055 4131
rect 6840 4128 6868 4168
rect 9398 4156 9404 4208
rect 9456 4196 9462 4208
rect 9907 4199 9965 4205
rect 9907 4196 9919 4199
rect 9456 4168 9919 4196
rect 9456 4156 9462 4168
rect 9907 4165 9919 4168
rect 9953 4165 9965 4199
rect 9907 4159 9965 4165
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 6840 4100 6929 4128
rect 5997 4091 6055 4097
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 7282 4128 7288 4140
rect 7243 4100 7288 4128
rect 6917 4091 6975 4097
rect 7282 4088 7288 4100
rect 7340 4128 7346 4140
rect 7650 4128 7656 4140
rect 7340 4100 7656 4128
rect 7340 4088 7346 4100
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 8294 4128 8300 4140
rect 8255 4100 8300 4128
rect 8294 4088 8300 4100
rect 8352 4128 8358 4140
rect 8938 4128 8944 4140
rect 8352 4100 8432 4128
rect 8899 4100 8944 4128
rect 8352 4088 8358 4100
rect 1486 4020 1492 4072
rect 1544 4060 1550 4072
rect 1857 4063 1915 4069
rect 1857 4060 1869 4063
rect 1544 4032 1869 4060
rect 1544 4020 1550 4032
rect 1857 4029 1869 4032
rect 1903 4029 1915 4063
rect 1857 4023 1915 4029
rect 2593 4063 2651 4069
rect 2593 4029 2605 4063
rect 2639 4060 2651 4063
rect 2682 4060 2688 4072
rect 2639 4032 2688 4060
rect 2639 4029 2651 4032
rect 2593 4023 2651 4029
rect 1765 3995 1823 4001
rect 1765 3961 1777 3995
rect 1811 3992 1823 3995
rect 2608 3992 2636 4023
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 3142 4020 3148 4072
rect 3200 4060 3206 4072
rect 3421 4063 3479 4069
rect 3421 4060 3433 4063
rect 3200 4032 3433 4060
rect 3200 4020 3206 4032
rect 3421 4029 3433 4032
rect 3467 4060 3479 4063
rect 3694 4060 3700 4072
rect 3467 4032 3700 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 3973 4063 4031 4069
rect 3973 4029 3985 4063
rect 4019 4060 4031 4063
rect 4246 4060 4252 4072
rect 4019 4032 4252 4060
rect 4019 4029 4031 4032
rect 3973 4023 4031 4029
rect 4246 4020 4252 4032
rect 4304 4060 4310 4072
rect 4706 4060 4712 4072
rect 4304 4032 4712 4060
rect 4304 4020 4310 4032
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 8404 4069 8432 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9030 4088 9036 4140
rect 9088 4128 9094 4140
rect 10054 4128 10082 4224
rect 15378 4196 15384 4208
rect 14016 4168 15384 4196
rect 9088 4100 10082 4128
rect 9088 4088 9094 4100
rect 10134 4088 10140 4140
rect 10192 4128 10198 4140
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 10192 4100 10237 4128
rect 12452 4100 13001 4128
rect 10192 4088 10198 4100
rect 8389 4063 8447 4069
rect 8389 4029 8401 4063
rect 8435 4029 8447 4063
rect 8570 4060 8576 4072
rect 8531 4032 8576 4060
rect 8389 4023 8447 4029
rect 4154 3992 4160 4004
rect 1811 3964 2636 3992
rect 4115 3964 4160 3992
rect 1811 3961 1823 3964
rect 1765 3955 1823 3961
rect 4154 3952 4160 3964
rect 4212 3952 4218 4004
rect 4798 3952 4804 4004
rect 4856 3992 4862 4004
rect 5077 3995 5135 4001
rect 5077 3992 5089 3995
rect 4856 3964 5089 3992
rect 4856 3952 4862 3964
rect 5077 3961 5089 3964
rect 5123 3961 5135 3995
rect 5077 3955 5135 3961
rect 5169 3995 5227 4001
rect 5169 3961 5181 3995
rect 5215 3961 5227 3995
rect 5169 3955 5227 3961
rect 4430 3924 4436 3936
rect 4391 3896 4436 3924
rect 4430 3884 4436 3896
rect 4488 3884 4494 3936
rect 4893 3927 4951 3933
rect 4893 3893 4905 3927
rect 4939 3924 4951 3927
rect 5184 3924 5212 3955
rect 5534 3952 5540 4004
rect 5592 3992 5598 4004
rect 5721 3995 5779 4001
rect 5721 3992 5733 3995
rect 5592 3964 5733 3992
rect 5592 3952 5598 3964
rect 5721 3961 5733 3964
rect 5767 3992 5779 3995
rect 6914 3992 6920 4004
rect 5767 3964 6920 3992
rect 5767 3961 5779 3964
rect 5721 3955 5779 3961
rect 6914 3952 6920 3964
rect 6972 3952 6978 4004
rect 7009 3995 7067 4001
rect 7009 3961 7021 3995
rect 7055 3961 7067 3995
rect 8404 3992 8432 4023
rect 8570 4020 8576 4032
rect 8628 4060 8634 4072
rect 9217 4063 9275 4069
rect 9217 4060 9229 4063
rect 8628 4032 9229 4060
rect 8628 4020 8634 4032
rect 9217 4029 9229 4032
rect 9263 4029 9275 4063
rect 9217 4023 9275 4029
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 9769 4063 9827 4069
rect 9769 4060 9781 4063
rect 9732 4032 9781 4060
rect 9732 4020 9738 4032
rect 9769 4029 9781 4032
rect 9815 4029 9827 4063
rect 11330 4060 11336 4072
rect 11291 4032 11336 4060
rect 9769 4023 9827 4029
rect 11330 4020 11336 4032
rect 11388 4060 11394 4072
rect 12452 4069 12480 4100
rect 12989 4097 13001 4100
rect 13035 4128 13047 4131
rect 13078 4128 13084 4140
rect 13035 4100 13084 4128
rect 13035 4097 13047 4100
rect 12989 4091 13047 4097
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 14016 4137 14044 4168
rect 15378 4156 15384 4168
rect 15436 4156 15442 4208
rect 15749 4199 15807 4205
rect 15749 4165 15761 4199
rect 15795 4196 15807 4199
rect 16206 4196 16212 4208
rect 15795 4168 16212 4196
rect 15795 4165 15807 4168
rect 15749 4159 15807 4165
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14424 4100 14657 4128
rect 14424 4088 14430 4100
rect 14645 4097 14657 4100
rect 14691 4128 14703 4131
rect 15764 4128 15792 4159
rect 16206 4156 16212 4168
rect 16264 4156 16270 4208
rect 17586 4196 17592 4208
rect 16500 4168 17592 4196
rect 14691 4100 15792 4128
rect 14691 4097 14703 4100
rect 14645 4091 14703 4097
rect 15838 4088 15844 4140
rect 15896 4128 15902 4140
rect 16298 4128 16304 4140
rect 15896 4100 16304 4128
rect 15896 4088 15902 4100
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 16500 4137 16528 4168
rect 17586 4156 17592 4168
rect 17644 4156 17650 4208
rect 17972 4168 19288 4196
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4097 16543 4131
rect 16485 4091 16543 4097
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17972 4128 18000 4168
rect 19260 4140 19288 4168
rect 19812 4168 20116 4196
rect 17175 4100 18000 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 19242 4088 19248 4140
rect 19300 4128 19306 4140
rect 19812 4128 19840 4168
rect 19300 4100 19840 4128
rect 19889 4131 19947 4137
rect 19300 4088 19306 4100
rect 19889 4097 19901 4131
rect 19935 4128 19947 4131
rect 19978 4128 19984 4140
rect 19935 4100 19984 4128
rect 19935 4097 19947 4100
rect 19889 4091 19947 4097
rect 19978 4088 19984 4100
rect 20036 4088 20042 4140
rect 20088 4128 20116 4168
rect 20162 4156 20168 4208
rect 20220 4196 20226 4208
rect 25314 4196 25320 4208
rect 20220 4168 25320 4196
rect 20220 4156 20226 4168
rect 25314 4156 25320 4168
rect 25372 4156 25378 4208
rect 22649 4131 22707 4137
rect 20088 4100 20576 4128
rect 11793 4063 11851 4069
rect 11793 4060 11805 4063
rect 11388 4032 11805 4060
rect 11388 4020 11394 4032
rect 11793 4029 11805 4032
rect 11839 4029 11851 4063
rect 11793 4023 11851 4029
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4060 18107 4063
rect 18138 4060 18144 4072
rect 18095 4032 18144 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 18138 4020 18144 4032
rect 18196 4020 18202 4072
rect 20548 4004 20576 4100
rect 22649 4097 22661 4131
rect 22695 4128 22707 4131
rect 23382 4128 23388 4140
rect 22695 4100 23388 4128
rect 22695 4097 22707 4100
rect 22649 4091 22707 4097
rect 23382 4088 23388 4100
rect 23440 4088 23446 4140
rect 25682 4128 25688 4140
rect 25240 4100 25688 4128
rect 22830 4020 22836 4072
rect 22888 4060 22894 4072
rect 23017 4063 23075 4069
rect 23017 4060 23029 4063
rect 22888 4032 23029 4060
rect 22888 4020 22894 4032
rect 23017 4029 23029 4032
rect 23063 4029 23075 4063
rect 23017 4023 23075 4029
rect 23477 4063 23535 4069
rect 23477 4029 23489 4063
rect 23523 4060 23535 4063
rect 23661 4063 23719 4069
rect 23661 4060 23673 4063
rect 23523 4032 23673 4060
rect 23523 4029 23535 4032
rect 23477 4023 23535 4029
rect 23661 4029 23673 4032
rect 23707 4060 23719 4063
rect 23750 4060 23756 4072
rect 23707 4032 23756 4060
rect 23707 4029 23719 4032
rect 23661 4023 23719 4029
rect 9122 3992 9128 4004
rect 8404 3964 9128 3992
rect 7009 3955 7067 3961
rect 6086 3924 6092 3936
rect 4939 3896 6092 3924
rect 4939 3893 4951 3896
rect 4893 3887 4951 3893
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6641 3927 6699 3933
rect 6641 3893 6653 3927
rect 6687 3924 6699 3927
rect 7024 3924 7052 3955
rect 9122 3952 9128 3964
rect 9180 3952 9186 4004
rect 14093 3995 14151 4001
rect 14093 3961 14105 3995
rect 14139 3961 14151 3995
rect 15378 3992 15384 4004
rect 15339 3964 15384 3992
rect 14093 3955 14151 3961
rect 7374 3924 7380 3936
rect 6687 3896 7380 3924
rect 6687 3893 6699 3896
rect 6641 3887 6699 3893
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 7653 3927 7711 3933
rect 7653 3893 7665 3927
rect 7699 3924 7711 3927
rect 10413 3927 10471 3933
rect 10413 3924 10425 3927
rect 7699 3896 10425 3924
rect 7699 3893 7711 3896
rect 7653 3887 7711 3893
rect 10413 3893 10425 3896
rect 10459 3893 10471 3927
rect 10413 3887 10471 3893
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11480 3896 11529 3924
rect 11480 3884 11486 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 12618 3924 12624 3936
rect 12579 3896 12624 3924
rect 11517 3887 11575 3893
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 13541 3927 13599 3933
rect 13541 3893 13553 3927
rect 13587 3924 13599 3927
rect 13630 3924 13636 3936
rect 13587 3896 13636 3924
rect 13587 3893 13599 3896
rect 13541 3887 13599 3893
rect 13630 3884 13636 3896
rect 13688 3924 13694 3936
rect 14108 3924 14136 3955
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 16574 3992 16580 4004
rect 16535 3964 16580 3992
rect 16574 3952 16580 3964
rect 16632 3952 16638 4004
rect 18370 3995 18428 4001
rect 18370 3961 18382 3995
rect 18416 3961 18428 3995
rect 19981 3995 20039 4001
rect 19981 3992 19993 3995
rect 18370 3955 18428 3961
rect 19260 3964 19993 3992
rect 14921 3927 14979 3933
rect 14921 3924 14933 3927
rect 13688 3896 14933 3924
rect 13688 3884 13694 3896
rect 14921 3893 14933 3896
rect 14967 3893 14979 3927
rect 17862 3924 17868 3936
rect 17823 3896 17868 3924
rect 14921 3887 14979 3893
rect 17862 3884 17868 3896
rect 17920 3924 17926 3936
rect 18385 3924 18413 3955
rect 19260 3936 19288 3964
rect 19981 3961 19993 3964
rect 20027 3961 20039 3995
rect 20530 3992 20536 4004
rect 20491 3964 20536 3992
rect 19981 3955 20039 3961
rect 20530 3952 20536 3964
rect 20588 3952 20594 4004
rect 21450 3952 21456 4004
rect 21508 3992 21514 4004
rect 22005 3995 22063 4001
rect 22005 3992 22017 3995
rect 21508 3964 22017 3992
rect 21508 3952 21514 3964
rect 22005 3961 22017 3964
rect 22051 3961 22063 3995
rect 22005 3955 22063 3961
rect 22094 3952 22100 4004
rect 22152 3992 22158 4004
rect 23032 3992 23060 4023
rect 23750 4020 23756 4032
rect 23808 4020 23814 4072
rect 24121 4063 24179 4069
rect 24121 4029 24133 4063
rect 24167 4060 24179 4063
rect 24210 4060 24216 4072
rect 24167 4032 24216 4060
rect 24167 4029 24179 4032
rect 24121 4023 24179 4029
rect 24136 3992 24164 4023
rect 24210 4020 24216 4032
rect 24268 4060 24274 4072
rect 24946 4060 24952 4072
rect 24268 4032 24952 4060
rect 24268 4020 24274 4032
rect 24946 4020 24952 4032
rect 25004 4060 25010 4072
rect 25240 4069 25268 4100
rect 25682 4088 25688 4100
rect 25740 4128 25746 4140
rect 25777 4131 25835 4137
rect 25777 4128 25789 4131
rect 25740 4100 25789 4128
rect 25740 4088 25746 4100
rect 25777 4097 25789 4100
rect 25823 4097 25835 4131
rect 25777 4091 25835 4097
rect 25041 4063 25099 4069
rect 25041 4060 25053 4063
rect 25004 4032 25053 4060
rect 25004 4020 25010 4032
rect 25041 4029 25053 4032
rect 25087 4029 25099 4063
rect 25041 4023 25099 4029
rect 25225 4063 25283 4069
rect 25225 4029 25237 4063
rect 25271 4029 25283 4063
rect 25225 4023 25283 4029
rect 22152 3964 22197 3992
rect 23032 3964 24164 3992
rect 22152 3952 22158 3964
rect 19242 3924 19248 3936
rect 17920 3896 18413 3924
rect 19203 3896 19248 3924
rect 17920 3884 17926 3896
rect 19242 3884 19248 3896
rect 19300 3884 19306 3936
rect 21082 3924 21088 3936
rect 21043 3896 21088 3924
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 23750 3924 23756 3936
rect 23711 3896 23756 3924
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 25409 3927 25467 3933
rect 25409 3893 25421 3927
rect 25455 3924 25467 3927
rect 25590 3924 25596 3936
rect 25455 3896 25596 3924
rect 25455 3893 25467 3896
rect 25409 3887 25467 3893
rect 25590 3884 25596 3896
rect 25648 3884 25654 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 2222 3720 2228 3732
rect 2183 3692 2228 3720
rect 2222 3680 2228 3692
rect 2280 3720 2286 3732
rect 2682 3720 2688 3732
rect 2280 3692 2688 3720
rect 2280 3680 2286 3692
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 2869 3723 2927 3729
rect 2869 3720 2881 3723
rect 2832 3692 2881 3720
rect 2832 3680 2838 3692
rect 2869 3689 2881 3692
rect 2915 3720 2927 3723
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 2915 3692 3433 3720
rect 2915 3689 2927 3692
rect 2869 3683 2927 3689
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 3421 3683 3479 3689
rect 3694 3680 3700 3732
rect 3752 3720 3758 3732
rect 3789 3723 3847 3729
rect 3789 3720 3801 3723
rect 3752 3692 3801 3720
rect 3752 3680 3758 3692
rect 3789 3689 3801 3692
rect 3835 3689 3847 3723
rect 4246 3720 4252 3732
rect 4207 3692 4252 3720
rect 3789 3683 3847 3689
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5353 3723 5411 3729
rect 5353 3720 5365 3723
rect 5132 3692 5365 3720
rect 5132 3680 5138 3692
rect 5353 3689 5365 3692
rect 5399 3720 5411 3723
rect 5629 3723 5687 3729
rect 5629 3720 5641 3723
rect 5399 3692 5641 3720
rect 5399 3689 5411 3692
rect 5353 3683 5411 3689
rect 5629 3689 5641 3692
rect 5675 3689 5687 3723
rect 6362 3720 6368 3732
rect 6323 3692 6368 3720
rect 5629 3683 5687 3689
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 8205 3723 8263 3729
rect 8205 3720 8217 3723
rect 7340 3692 8217 3720
rect 7340 3680 7346 3692
rect 8205 3689 8217 3692
rect 8251 3689 8263 3723
rect 9398 3720 9404 3732
rect 9359 3692 9404 3720
rect 8205 3683 8263 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 9861 3723 9919 3729
rect 9861 3720 9873 3723
rect 9732 3692 9873 3720
rect 9732 3680 9738 3692
rect 9861 3689 9873 3692
rect 9907 3689 9919 3723
rect 9861 3683 9919 3689
rect 10134 3680 10140 3732
rect 10192 3720 10198 3732
rect 10229 3723 10287 3729
rect 10229 3720 10241 3723
rect 10192 3692 10241 3720
rect 10192 3680 10198 3692
rect 10229 3689 10241 3692
rect 10275 3689 10287 3723
rect 12437 3723 12495 3729
rect 12437 3720 12449 3723
rect 10229 3683 10287 3689
rect 11992 3692 12449 3720
rect 4798 3661 4804 3664
rect 4795 3652 4804 3661
rect 4759 3624 4804 3652
rect 4795 3615 4804 3624
rect 4798 3612 4804 3615
rect 4856 3612 4862 3664
rect 7374 3652 7380 3664
rect 7335 3624 7380 3652
rect 7374 3612 7380 3624
rect 7432 3612 7438 3664
rect 7742 3612 7748 3664
rect 7800 3652 7806 3664
rect 8665 3655 8723 3661
rect 8665 3652 8677 3655
rect 7800 3624 8677 3652
rect 7800 3612 7806 3624
rect 8665 3621 8677 3624
rect 8711 3652 8723 3655
rect 9214 3652 9220 3664
rect 8711 3624 9220 3652
rect 8711 3621 8723 3624
rect 8665 3615 8723 3621
rect 9214 3612 9220 3624
rect 9272 3612 9278 3664
rect 10042 3612 10048 3664
rect 10100 3652 10106 3664
rect 10597 3655 10655 3661
rect 10597 3652 10609 3655
rect 10100 3624 10609 3652
rect 10100 3612 10106 3624
rect 10597 3621 10609 3624
rect 10643 3652 10655 3655
rect 11609 3655 11667 3661
rect 11609 3652 11621 3655
rect 10643 3624 11621 3652
rect 10643 3621 10655 3624
rect 10597 3615 10655 3621
rect 11609 3621 11621 3624
rect 11655 3621 11667 3655
rect 11609 3615 11667 3621
rect 1486 3593 1492 3596
rect 1464 3587 1492 3593
rect 1464 3553 1476 3587
rect 1464 3547 1492 3553
rect 1486 3544 1492 3547
rect 1544 3544 1550 3596
rect 2866 3584 2872 3596
rect 2827 3556 2872 3584
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4433 3587 4491 3593
rect 4433 3584 4445 3587
rect 4212 3556 4445 3584
rect 4212 3544 4218 3556
rect 4433 3553 4445 3556
rect 4479 3584 4491 3587
rect 5997 3587 6055 3593
rect 5997 3584 6009 3587
rect 4479 3556 6009 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 5997 3553 6009 3556
rect 6043 3553 6055 3587
rect 6178 3584 6184 3596
rect 6139 3556 6184 3584
rect 5997 3547 6055 3553
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 10778 3593 10784 3596
rect 10744 3587 10784 3593
rect 10744 3553 10756 3587
rect 10744 3547 10784 3553
rect 10778 3544 10784 3547
rect 10836 3544 10842 3596
rect 1946 3476 1952 3528
rect 2004 3516 2010 3528
rect 7101 3519 7159 3525
rect 7101 3516 7113 3519
rect 2004 3488 7113 3516
rect 2004 3476 2010 3488
rect 7101 3485 7113 3488
rect 7147 3485 7159 3519
rect 7282 3516 7288 3528
rect 7243 3488 7288 3516
rect 7101 3479 7159 3485
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7561 3519 7619 3525
rect 7561 3485 7573 3519
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 7576 3448 7604 3479
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 9456 3488 10977 3516
rect 9456 3476 9462 3488
rect 10965 3485 10977 3488
rect 11011 3516 11023 3519
rect 11330 3516 11336 3528
rect 11011 3488 11336 3516
rect 11011 3485 11023 3488
rect 10965 3479 11023 3485
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 6972 3420 7604 3448
rect 6972 3408 6978 3420
rect 9858 3408 9864 3460
rect 9916 3448 9922 3460
rect 11992 3457 12020 3692
rect 12437 3689 12449 3692
rect 12483 3689 12495 3723
rect 12437 3683 12495 3689
rect 14274 3680 14280 3732
rect 14332 3720 14338 3732
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 14332 3692 14657 3720
rect 14332 3680 14338 3692
rect 14645 3689 14657 3692
rect 14691 3689 14703 3723
rect 14645 3683 14703 3689
rect 16485 3723 16543 3729
rect 16485 3689 16497 3723
rect 16531 3720 16543 3723
rect 16574 3720 16580 3732
rect 16531 3692 16580 3720
rect 16531 3689 16543 3692
rect 16485 3683 16543 3689
rect 16574 3680 16580 3692
rect 16632 3720 16638 3732
rect 19978 3720 19984 3732
rect 16632 3692 18460 3720
rect 19939 3692 19984 3720
rect 16632 3680 16638 3692
rect 18432 3664 18460 3692
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 20070 3680 20076 3732
rect 20128 3720 20134 3732
rect 20257 3723 20315 3729
rect 20257 3720 20269 3723
rect 20128 3692 20269 3720
rect 20128 3680 20134 3692
rect 20257 3689 20269 3692
rect 20303 3689 20315 3723
rect 21174 3720 21180 3732
rect 21135 3692 21180 3720
rect 20257 3683 20315 3689
rect 21174 3680 21180 3692
rect 21232 3680 21238 3732
rect 22646 3720 22652 3732
rect 22607 3692 22652 3720
rect 22646 3680 22652 3692
rect 22704 3680 22710 3732
rect 23474 3720 23480 3732
rect 23435 3692 23480 3720
rect 23474 3680 23480 3692
rect 23532 3680 23538 3732
rect 24854 3720 24860 3732
rect 24815 3692 24860 3720
rect 24854 3680 24860 3692
rect 24912 3680 24918 3732
rect 12158 3652 12164 3664
rect 12119 3624 12164 3652
rect 12158 3612 12164 3624
rect 12216 3612 12222 3664
rect 13814 3652 13820 3664
rect 13775 3624 13820 3652
rect 13814 3612 13820 3624
rect 13872 3612 13878 3664
rect 14366 3652 14372 3664
rect 14327 3624 14372 3652
rect 14366 3612 14372 3624
rect 14424 3612 14430 3664
rect 15470 3652 15476 3664
rect 15431 3624 15476 3652
rect 15470 3612 15476 3624
rect 15528 3612 15534 3664
rect 16025 3655 16083 3661
rect 16025 3621 16037 3655
rect 16071 3652 16083 3655
rect 16206 3652 16212 3664
rect 16071 3624 16212 3652
rect 16071 3621 16083 3624
rect 16025 3615 16083 3621
rect 16206 3612 16212 3624
rect 16264 3612 16270 3664
rect 16850 3652 16856 3664
rect 16811 3624 16856 3652
rect 16850 3612 16856 3624
rect 16908 3612 16914 3664
rect 18414 3652 18420 3664
rect 18375 3624 18420 3652
rect 18414 3612 18420 3624
rect 18472 3612 18478 3664
rect 18966 3652 18972 3664
rect 18927 3624 18972 3652
rect 18966 3612 18972 3624
rect 19024 3652 19030 3664
rect 21450 3652 21456 3664
rect 19024 3624 21456 3652
rect 19024 3612 19030 3624
rect 21450 3612 21456 3624
rect 21508 3612 21514 3664
rect 21726 3612 21732 3664
rect 21784 3652 21790 3664
rect 21821 3655 21879 3661
rect 21821 3652 21833 3655
rect 21784 3624 21833 3652
rect 21784 3612 21790 3624
rect 21821 3621 21833 3624
rect 21867 3621 21879 3655
rect 21821 3615 21879 3621
rect 22186 3612 22192 3664
rect 22244 3652 22250 3664
rect 23017 3655 23075 3661
rect 23017 3652 23029 3655
rect 22244 3624 23029 3652
rect 22244 3612 22250 3624
rect 23017 3621 23029 3624
rect 23063 3652 23075 3655
rect 23063 3624 23704 3652
rect 23063 3621 23075 3624
rect 23017 3615 23075 3621
rect 12176 3516 12204 3612
rect 12250 3544 12256 3596
rect 12308 3584 12314 3596
rect 12345 3587 12403 3593
rect 12345 3584 12357 3587
rect 12308 3556 12357 3584
rect 12308 3544 12314 3556
rect 12345 3553 12357 3556
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 16942 3544 16948 3596
rect 17000 3584 17006 3596
rect 17129 3587 17187 3593
rect 17129 3584 17141 3587
rect 17000 3556 17141 3584
rect 17000 3544 17006 3556
rect 17129 3553 17141 3556
rect 17175 3553 17187 3587
rect 17129 3547 17187 3553
rect 19797 3587 19855 3593
rect 19797 3553 19809 3587
rect 19843 3584 19855 3587
rect 20162 3584 20168 3596
rect 19843 3556 20168 3584
rect 19843 3553 19855 3556
rect 19797 3547 19855 3553
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 20806 3544 20812 3596
rect 20864 3544 20870 3596
rect 22738 3544 22744 3596
rect 22796 3584 22802 3596
rect 23676 3593 23704 3624
rect 24946 3612 24952 3664
rect 25004 3652 25010 3664
rect 25004 3624 25268 3652
rect 25004 3612 25010 3624
rect 23201 3587 23259 3593
rect 23201 3584 23213 3587
rect 22796 3556 23213 3584
rect 22796 3544 22802 3556
rect 23201 3553 23213 3556
rect 23247 3553 23259 3587
rect 23201 3547 23259 3553
rect 23661 3587 23719 3593
rect 23661 3553 23673 3587
rect 23707 3553 23719 3587
rect 25038 3584 25044 3596
rect 24999 3556 25044 3584
rect 23661 3547 23719 3553
rect 25038 3544 25044 3556
rect 25096 3544 25102 3596
rect 25240 3593 25268 3624
rect 25225 3587 25283 3593
rect 25225 3553 25237 3587
rect 25271 3584 25283 3587
rect 25314 3584 25320 3596
rect 25271 3556 25320 3584
rect 25271 3553 25283 3556
rect 25225 3547 25283 3553
rect 25314 3544 25320 3556
rect 25372 3544 25378 3596
rect 12989 3519 13047 3525
rect 12989 3516 13001 3519
rect 12176 3488 13001 3516
rect 12989 3485 13001 3488
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3516 13783 3519
rect 14182 3516 14188 3528
rect 13771 3488 14188 3516
rect 13771 3485 13783 3488
rect 13725 3479 13783 3485
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3516 15163 3519
rect 15378 3516 15384 3528
rect 15151 3488 15384 3516
rect 15151 3485 15163 3488
rect 15105 3479 15163 3485
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3516 17831 3519
rect 18322 3516 18328 3528
rect 17819 3488 18328 3516
rect 17819 3485 17831 3488
rect 17773 3479 17831 3485
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 18782 3476 18788 3528
rect 18840 3516 18846 3528
rect 19337 3519 19395 3525
rect 19337 3516 19349 3519
rect 18840 3488 19349 3516
rect 18840 3476 18846 3488
rect 19337 3485 19349 3488
rect 19383 3516 19395 3519
rect 20824 3516 20852 3544
rect 19383 3488 20852 3516
rect 21729 3519 21787 3525
rect 19383 3485 19395 3488
rect 19337 3479 19395 3485
rect 21729 3485 21741 3519
rect 21775 3516 21787 3519
rect 21910 3516 21916 3528
rect 21775 3488 21916 3516
rect 21775 3485 21787 3488
rect 21729 3479 21787 3485
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 22373 3519 22431 3525
rect 22373 3485 22385 3519
rect 22419 3516 22431 3519
rect 23014 3516 23020 3528
rect 22419 3488 23020 3516
rect 22419 3485 22431 3488
rect 22373 3479 22431 3485
rect 23014 3476 23020 3488
rect 23072 3516 23078 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 23072 3488 24593 3516
rect 23072 3476 23078 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 11977 3451 12035 3457
rect 11977 3448 11989 3451
rect 9916 3420 11989 3448
rect 9916 3408 9922 3420
rect 11977 3417 11989 3420
rect 12023 3417 12035 3451
rect 11977 3411 12035 3417
rect 1535 3383 1593 3389
rect 1535 3349 1547 3383
rect 1581 3380 1593 3383
rect 1762 3380 1768 3392
rect 1581 3352 1768 3380
rect 1581 3349 1593 3352
rect 1535 3343 1593 3349
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 1946 3380 1952 3392
rect 1907 3352 1952 3380
rect 1946 3340 1952 3352
rect 2004 3340 2010 3392
rect 7006 3380 7012 3392
rect 6967 3352 7012 3380
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7101 3383 7159 3389
rect 7101 3349 7113 3383
rect 7147 3380 7159 3383
rect 9030 3380 9036 3392
rect 7147 3352 9036 3380
rect 7147 3349 7159 3352
rect 7101 3343 7159 3349
rect 9030 3340 9036 3352
rect 9088 3340 9094 3392
rect 10502 3340 10508 3392
rect 10560 3380 10566 3392
rect 10873 3383 10931 3389
rect 10873 3380 10885 3383
rect 10560 3352 10885 3380
rect 10560 3340 10566 3352
rect 10873 3349 10885 3352
rect 10919 3380 10931 3383
rect 10962 3380 10968 3392
rect 10919 3352 10968 3380
rect 10919 3349 10931 3352
rect 10873 3343 10931 3349
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11238 3380 11244 3392
rect 11199 3352 11244 3380
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 12802 3340 12808 3392
rect 12860 3380 12866 3392
rect 13357 3383 13415 3389
rect 13357 3380 13369 3383
rect 12860 3352 13369 3380
rect 12860 3340 12866 3352
rect 13357 3349 13369 3352
rect 13403 3349 13415 3383
rect 17310 3380 17316 3392
rect 17271 3352 17316 3380
rect 13357 3343 13415 3349
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 18138 3380 18144 3392
rect 18099 3352 18144 3380
rect 18138 3340 18144 3352
rect 18196 3340 18202 3392
rect 24210 3380 24216 3392
rect 24171 3352 24216 3380
rect 24210 3340 24216 3352
rect 24268 3340 24274 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1486 3136 1492 3188
rect 1544 3176 1550 3188
rect 1581 3179 1639 3185
rect 1581 3176 1593 3179
rect 1544 3148 1593 3176
rect 1544 3136 1550 3148
rect 1581 3145 1593 3148
rect 1627 3145 1639 3179
rect 2866 3176 2872 3188
rect 2827 3148 2872 3176
rect 1581 3139 1639 3145
rect 2866 3136 2872 3148
rect 2924 3176 2930 3188
rect 6178 3176 6184 3188
rect 2924 3148 6184 3176
rect 2924 3136 2930 3148
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 6641 3179 6699 3185
rect 6641 3145 6653 3179
rect 6687 3176 6699 3179
rect 6822 3176 6828 3188
rect 6687 3148 6828 3176
rect 6687 3145 6699 3148
rect 6641 3139 6699 3145
rect 5534 3108 5540 3120
rect 5495 3080 5540 3108
rect 5534 3068 5540 3080
rect 5592 3068 5598 3120
rect 2590 3000 2596 3052
rect 2648 3040 2654 3052
rect 3145 3043 3203 3049
rect 3145 3040 3157 3043
rect 2648 3012 3157 3040
rect 2648 3000 2654 3012
rect 3145 3009 3157 3012
rect 3191 3040 3203 3043
rect 3234 3040 3240 3052
rect 3191 3012 3240 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3040 4583 3043
rect 4798 3040 4804 3052
rect 4571 3012 4804 3040
rect 4571 3009 4583 3012
rect 4525 3003 4583 3009
rect 4798 3000 4804 3012
rect 4856 3040 4862 3052
rect 6656 3040 6684 3139
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7432 3148 7849 3176
rect 7432 3136 7438 3148
rect 7837 3145 7849 3148
rect 7883 3176 7895 3179
rect 8113 3179 8171 3185
rect 8113 3176 8125 3179
rect 7883 3148 8125 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 8113 3145 8125 3148
rect 8159 3145 8171 3179
rect 9766 3176 9772 3188
rect 9727 3148 9772 3176
rect 8113 3139 8171 3145
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 10045 3179 10103 3185
rect 10045 3176 10057 3179
rect 10008 3148 10057 3176
rect 10008 3136 10014 3148
rect 10045 3145 10057 3148
rect 10091 3145 10103 3179
rect 10045 3139 10103 3145
rect 10394 3179 10452 3185
rect 10394 3145 10406 3179
rect 10440 3176 10452 3179
rect 10778 3176 10784 3188
rect 10440 3148 10784 3176
rect 10440 3145 10452 3148
rect 10394 3139 10452 3145
rect 8570 3040 8576 3052
rect 4856 3012 6684 3040
rect 8483 3012 8576 3040
rect 4856 3000 4862 3012
rect 1946 2972 1952 2984
rect 1907 2944 1952 2972
rect 1946 2932 1952 2944
rect 2004 2972 2010 2984
rect 2314 2972 2320 2984
rect 2004 2944 2320 2972
rect 2004 2932 2010 2944
rect 2314 2932 2320 2944
rect 2372 2932 2378 2984
rect 3418 2972 3424 2984
rect 3379 2944 3424 2972
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 3786 2972 3792 2984
rect 3747 2944 3792 2972
rect 3786 2932 3792 2944
rect 3844 2932 3850 2984
rect 2498 2904 2504 2916
rect 2459 2876 2504 2904
rect 2498 2864 2504 2876
rect 2556 2864 2562 2916
rect 3970 2864 3976 2916
rect 4028 2904 4034 2916
rect 4065 2907 4123 2913
rect 4065 2904 4077 2907
rect 4028 2876 4077 2904
rect 4028 2864 4034 2876
rect 4065 2873 4077 2876
rect 4111 2873 4123 2907
rect 4982 2904 4988 2916
rect 4943 2876 4988 2904
rect 4065 2867 4123 2873
rect 4982 2864 4988 2876
rect 5040 2864 5046 2916
rect 5074 2864 5080 2916
rect 5132 2904 5138 2916
rect 6656 2904 6684 3012
rect 8570 3000 8576 3012
rect 8628 3040 8634 3052
rect 9306 3040 9312 3052
rect 8628 3012 9312 3040
rect 8628 3000 8634 3012
rect 6917 2975 6975 2981
rect 6917 2941 6929 2975
rect 6963 2972 6975 2975
rect 7006 2972 7012 2984
rect 6963 2944 7012 2972
rect 6963 2941 6975 2944
rect 6917 2935 6975 2941
rect 7006 2932 7012 2944
rect 7064 2972 7070 2984
rect 8956 2981 8984 3012
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 10060 3040 10088 3139
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 10962 3136 10968 3188
rect 11020 3176 11026 3188
rect 11241 3179 11299 3185
rect 11241 3176 11253 3179
rect 11020 3148 11253 3176
rect 11020 3136 11026 3148
rect 11241 3145 11253 3148
rect 11287 3145 11299 3179
rect 12158 3176 12164 3188
rect 12119 3148 12164 3176
rect 11241 3139 11299 3145
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 13725 3179 13783 3185
rect 13725 3145 13737 3179
rect 13771 3176 13783 3179
rect 13814 3176 13820 3188
rect 13771 3148 13820 3176
rect 13771 3145 13783 3148
rect 13725 3139 13783 3145
rect 13814 3136 13820 3148
rect 13872 3176 13878 3188
rect 14001 3179 14059 3185
rect 14001 3176 14013 3179
rect 13872 3148 14013 3176
rect 13872 3136 13878 3148
rect 14001 3145 14013 3148
rect 14047 3145 14059 3179
rect 15470 3176 15476 3188
rect 15431 3148 15476 3176
rect 14001 3139 14059 3145
rect 15470 3136 15476 3148
rect 15528 3176 15534 3188
rect 15749 3179 15807 3185
rect 15749 3176 15761 3179
rect 15528 3148 15761 3176
rect 15528 3136 15534 3148
rect 15749 3145 15761 3148
rect 15795 3176 15807 3179
rect 16025 3179 16083 3185
rect 16025 3176 16037 3179
rect 15795 3148 16037 3176
rect 15795 3145 15807 3148
rect 15749 3139 15807 3145
rect 16025 3145 16037 3148
rect 16071 3176 16083 3179
rect 16117 3179 16175 3185
rect 16117 3176 16129 3179
rect 16071 3148 16129 3176
rect 16071 3145 16083 3148
rect 16025 3139 16083 3145
rect 16117 3145 16129 3148
rect 16163 3145 16175 3179
rect 16117 3139 16175 3145
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 17313 3179 17371 3185
rect 17313 3176 17325 3179
rect 17000 3148 17325 3176
rect 17000 3136 17006 3148
rect 17313 3145 17325 3148
rect 17359 3145 17371 3179
rect 17313 3139 17371 3145
rect 19889 3179 19947 3185
rect 19889 3145 19901 3179
rect 19935 3176 19947 3179
rect 20162 3176 20168 3188
rect 19935 3148 20168 3176
rect 19935 3145 19947 3148
rect 19889 3139 19947 3145
rect 20162 3136 20168 3148
rect 20220 3136 20226 3188
rect 22370 3136 22376 3188
rect 22428 3176 22434 3188
rect 22695 3179 22753 3185
rect 22695 3176 22707 3179
rect 22428 3148 22707 3176
rect 22428 3136 22434 3148
rect 22695 3145 22707 3148
rect 22741 3145 22753 3179
rect 22695 3139 22753 3145
rect 23109 3179 23167 3185
rect 23109 3145 23121 3179
rect 23155 3176 23167 3179
rect 23198 3176 23204 3188
rect 23155 3148 23204 3176
rect 23155 3145 23167 3148
rect 23109 3139 23167 3145
rect 10502 3108 10508 3120
rect 10463 3080 10508 3108
rect 10502 3068 10508 3080
rect 10560 3068 10566 3120
rect 10686 3108 10692 3120
rect 10647 3080 10692 3108
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 10597 3043 10655 3049
rect 10597 3040 10609 3043
rect 10060 3012 10609 3040
rect 10597 3009 10609 3012
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 12802 3040 12808 3052
rect 12492 3012 12808 3040
rect 12492 3000 12498 3012
rect 12802 3000 12808 3012
rect 12860 3000 12866 3052
rect 16393 3043 16451 3049
rect 16393 3009 16405 3043
rect 16439 3040 16451 3043
rect 16850 3040 16856 3052
rect 16439 3012 16856 3040
rect 16439 3009 16451 3012
rect 16393 3003 16451 3009
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 17034 3040 17040 3052
rect 16995 3012 17040 3040
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 18782 3040 18788 3052
rect 18743 3012 18788 3040
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 18966 3000 18972 3052
rect 19024 3040 19030 3052
rect 19061 3043 19119 3049
rect 19061 3040 19073 3043
rect 19024 3012 19073 3040
rect 19024 3000 19030 3012
rect 19061 3009 19073 3012
rect 19107 3009 19119 3043
rect 19061 3003 19119 3009
rect 20349 3043 20407 3049
rect 20349 3009 20361 3043
rect 20395 3040 20407 3043
rect 20806 3040 20812 3052
rect 20395 3012 20812 3040
rect 20395 3009 20407 3012
rect 20349 3003 20407 3009
rect 20806 3000 20812 3012
rect 20864 3000 20870 3052
rect 22465 3043 22523 3049
rect 22465 3009 22477 3043
rect 22511 3040 22523 3043
rect 22738 3040 22744 3052
rect 22511 3012 22744 3040
rect 22511 3009 22523 3012
rect 22465 3003 22523 3009
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 8941 2975 8999 2981
rect 7064 2944 7604 2972
rect 7064 2932 7070 2944
rect 7238 2907 7296 2913
rect 7238 2904 7250 2907
rect 5132 2876 5177 2904
rect 6656 2876 7250 2904
rect 5132 2864 5138 2876
rect 7238 2873 7250 2876
rect 7284 2873 7296 2907
rect 7576 2904 7604 2944
rect 8941 2941 8953 2975
rect 8987 2941 8999 2975
rect 9214 2972 9220 2984
rect 9175 2944 9220 2972
rect 8941 2935 8999 2941
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 10229 2975 10287 2981
rect 10229 2972 10241 2975
rect 9916 2944 10241 2972
rect 9916 2932 9922 2944
rect 10229 2941 10241 2944
rect 10275 2941 10287 2975
rect 10229 2935 10287 2941
rect 11330 2932 11336 2984
rect 11388 2972 11394 2984
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 11388 2944 11713 2972
rect 11388 2932 11394 2944
rect 11701 2941 11713 2944
rect 11747 2972 11759 2975
rect 12894 2972 12900 2984
rect 11747 2944 12900 2972
rect 11747 2941 11759 2944
rect 11701 2935 11759 2941
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 14550 2972 14556 2984
rect 14511 2944 14556 2972
rect 14550 2932 14556 2944
rect 14608 2932 14614 2984
rect 22624 2975 22682 2981
rect 22624 2941 22636 2975
rect 22670 2972 22682 2975
rect 23124 2972 23152 3139
rect 23198 3136 23204 3148
rect 23256 3136 23262 3188
rect 23477 3179 23535 3185
rect 23477 3145 23489 3179
rect 23523 3176 23535 3179
rect 23566 3176 23572 3188
rect 23523 3148 23572 3176
rect 23523 3145 23535 3148
rect 23477 3139 23535 3145
rect 23566 3136 23572 3148
rect 23624 3136 23630 3188
rect 23750 3136 23756 3188
rect 23808 3185 23814 3188
rect 23808 3179 23857 3185
rect 23808 3145 23811 3179
rect 23845 3176 23857 3179
rect 24673 3179 24731 3185
rect 24673 3176 24685 3179
rect 23845 3148 24685 3176
rect 23845 3145 23857 3148
rect 23808 3139 23857 3145
rect 24673 3145 24685 3148
rect 24719 3145 24731 3179
rect 25038 3176 25044 3188
rect 24999 3148 25044 3176
rect 24673 3139 24731 3145
rect 23808 3136 23814 3139
rect 25038 3136 25044 3148
rect 25096 3136 25102 3188
rect 25314 3136 25320 3188
rect 25372 3176 25378 3188
rect 25777 3179 25835 3185
rect 25777 3176 25789 3179
rect 25372 3148 25789 3176
rect 25372 3136 25378 3148
rect 25777 3145 25789 3148
rect 25823 3145 25835 3179
rect 25777 3139 25835 3145
rect 23382 3068 23388 3120
rect 23440 3108 23446 3120
rect 23937 3111 23995 3117
rect 23937 3108 23949 3111
rect 23440 3080 23949 3108
rect 23440 3068 23446 3080
rect 23937 3077 23949 3080
rect 23983 3077 23995 3111
rect 23937 3071 23995 3077
rect 24026 3040 24032 3052
rect 23939 3012 24032 3040
rect 24026 3000 24032 3012
rect 24084 3040 24090 3052
rect 24210 3040 24216 3052
rect 24084 3012 24216 3040
rect 24084 3000 24090 3012
rect 24210 3000 24216 3012
rect 24268 3000 24274 3052
rect 22670 2944 23152 2972
rect 22670 2941 22682 2944
rect 22624 2935 22682 2941
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23624 2944 23673 2972
rect 23624 2932 23630 2944
rect 23661 2941 23673 2944
rect 23707 2941 23719 2975
rect 25222 2972 25228 2984
rect 25135 2944 25228 2972
rect 23661 2935 23719 2941
rect 25222 2932 25228 2944
rect 25280 2972 25286 2984
rect 26145 2975 26203 2981
rect 26145 2972 26157 2975
rect 25280 2944 26157 2972
rect 25280 2932 25286 2944
rect 26145 2941 26157 2944
rect 26191 2941 26203 2975
rect 26145 2935 26203 2941
rect 13126 2907 13184 2913
rect 13126 2904 13138 2907
rect 7576 2876 8800 2904
rect 7238 2867 7296 2873
rect 8772 2845 8800 2876
rect 12636 2876 13138 2904
rect 12636 2848 12664 2876
rect 13126 2873 13138 2876
rect 13172 2904 13184 2907
rect 14369 2907 14427 2913
rect 14369 2904 14381 2907
rect 13172 2876 14381 2904
rect 13172 2873 13184 2876
rect 13126 2867 13184 2873
rect 14369 2873 14381 2876
rect 14415 2904 14427 2907
rect 14874 2907 14932 2913
rect 14874 2904 14886 2907
rect 14415 2876 14886 2904
rect 14415 2873 14427 2876
rect 14369 2867 14427 2873
rect 14874 2873 14886 2876
rect 14920 2904 14932 2907
rect 15654 2904 15660 2916
rect 14920 2876 15660 2904
rect 14920 2873 14932 2876
rect 14874 2867 14932 2873
rect 15654 2864 15660 2876
rect 15712 2904 15718 2916
rect 16206 2904 16212 2916
rect 15712 2876 16212 2904
rect 15712 2864 15718 2876
rect 16206 2864 16212 2876
rect 16264 2864 16270 2916
rect 16485 2907 16543 2913
rect 16485 2873 16497 2907
rect 16531 2873 16543 2907
rect 16485 2867 16543 2873
rect 18325 2907 18383 2913
rect 18325 2873 18337 2907
rect 18371 2904 18383 2907
rect 18414 2904 18420 2916
rect 18371 2876 18420 2904
rect 18371 2873 18383 2876
rect 18325 2867 18383 2873
rect 8757 2839 8815 2845
rect 8757 2805 8769 2839
rect 8803 2805 8815 2839
rect 12618 2836 12624 2848
rect 12579 2808 12624 2836
rect 8757 2799 8815 2805
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 16025 2839 16083 2845
rect 16025 2805 16037 2839
rect 16071 2836 16083 2839
rect 16500 2836 16528 2867
rect 18414 2864 18420 2876
rect 18472 2864 18478 2916
rect 18877 2907 18935 2913
rect 18877 2873 18889 2907
rect 18923 2904 18935 2907
rect 19242 2904 19248 2916
rect 18923 2876 19248 2904
rect 18923 2873 18935 2876
rect 18877 2867 18935 2873
rect 16071 2808 16528 2836
rect 16071 2805 16083 2808
rect 16025 2799 16083 2805
rect 17402 2796 17408 2848
rect 17460 2836 17466 2848
rect 17773 2839 17831 2845
rect 17773 2836 17785 2839
rect 17460 2808 17785 2836
rect 17460 2796 17466 2808
rect 17773 2805 17785 2808
rect 17819 2836 17831 2839
rect 18892 2836 18920 2867
rect 19242 2864 19248 2876
rect 19300 2864 19306 2916
rect 20717 2907 20775 2913
rect 20717 2873 20729 2907
rect 20763 2904 20775 2907
rect 21082 2904 21088 2916
rect 20763 2876 21088 2904
rect 20763 2873 20775 2876
rect 20717 2867 20775 2873
rect 21082 2864 21088 2876
rect 21140 2913 21146 2916
rect 21140 2907 21188 2913
rect 21140 2873 21142 2907
rect 21176 2873 21188 2907
rect 21140 2867 21188 2873
rect 23768 2876 25452 2904
rect 21140 2864 21146 2867
rect 21726 2836 21732 2848
rect 17819 2808 18920 2836
rect 21687 2808 21732 2836
rect 17819 2805 17831 2808
rect 17773 2799 17831 2805
rect 21726 2796 21732 2808
rect 21784 2836 21790 2848
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 21784 2808 22017 2836
rect 21784 2796 21790 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22005 2799 22063 2805
rect 23566 2796 23572 2848
rect 23624 2836 23630 2848
rect 23768 2836 23796 2876
rect 23624 2808 23796 2836
rect 23624 2796 23630 2808
rect 23842 2796 23848 2848
rect 23900 2836 23906 2848
rect 25424 2845 25452 2876
rect 24305 2839 24363 2845
rect 24305 2836 24317 2839
rect 23900 2808 24317 2836
rect 23900 2796 23906 2808
rect 24305 2805 24317 2808
rect 24351 2805 24363 2839
rect 24305 2799 24363 2805
rect 25409 2839 25467 2845
rect 25409 2805 25421 2839
rect 25455 2805 25467 2839
rect 25409 2799 25467 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 3786 2632 3792 2644
rect 3747 2604 3792 2632
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 4798 2592 4804 2644
rect 4856 2632 4862 2644
rect 4985 2635 5043 2641
rect 4985 2632 4997 2635
rect 4856 2604 4997 2632
rect 4856 2592 4862 2604
rect 4985 2601 4997 2604
rect 5031 2601 5043 2635
rect 4985 2595 5043 2601
rect 5997 2635 6055 2641
rect 5997 2601 6009 2635
rect 6043 2632 6055 2635
rect 6086 2632 6092 2644
rect 6043 2604 6092 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 4522 2564 4528 2576
rect 2976 2536 4528 2564
rect 1486 2505 1492 2508
rect 1464 2499 1492 2505
rect 1464 2465 1476 2499
rect 1544 2496 1550 2508
rect 2976 2505 3004 2536
rect 4522 2524 4528 2536
rect 4580 2524 4586 2576
rect 5000 2564 5028 2595
rect 6086 2592 6092 2604
rect 6144 2632 6150 2644
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 6144 2604 6653 2632
rect 6144 2592 6150 2604
rect 6641 2601 6653 2604
rect 6687 2632 6699 2635
rect 6687 2604 7144 2632
rect 6687 2601 6699 2604
rect 6641 2595 6699 2601
rect 7116 2573 7144 2604
rect 7834 2592 7840 2644
rect 7892 2632 7898 2644
rect 7929 2635 7987 2641
rect 7929 2632 7941 2635
rect 7892 2604 7941 2632
rect 7892 2592 7898 2604
rect 7929 2601 7941 2604
rect 7975 2601 7987 2635
rect 7929 2595 7987 2601
rect 8662 2592 8668 2644
rect 8720 2632 8726 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8720 2604 9137 2632
rect 8720 2592 8726 2604
rect 9125 2601 9137 2604
rect 9171 2632 9183 2635
rect 9582 2632 9588 2644
rect 9171 2604 9588 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 11146 2632 11152 2644
rect 9784 2604 11152 2632
rect 5439 2567 5497 2573
rect 5439 2564 5451 2567
rect 5000 2536 5451 2564
rect 5439 2533 5451 2536
rect 5485 2533 5497 2567
rect 5439 2527 5497 2533
rect 7101 2567 7159 2573
rect 7101 2533 7113 2567
rect 7147 2533 7159 2567
rect 7650 2564 7656 2576
rect 7611 2536 7656 2564
rect 7101 2527 7159 2533
rect 7650 2524 7656 2536
rect 7708 2524 7714 2576
rect 8294 2564 8300 2576
rect 8255 2536 8300 2564
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1544 2468 1869 2496
rect 1464 2459 1492 2465
rect 1486 2456 1492 2459
rect 1544 2456 1550 2468
rect 1857 2465 1869 2468
rect 1903 2465 1915 2499
rect 1857 2459 1915 2465
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2496 2375 2499
rect 2685 2499 2743 2505
rect 2685 2496 2697 2499
rect 2363 2468 2697 2496
rect 2363 2465 2375 2468
rect 2317 2459 2375 2465
rect 2685 2465 2697 2468
rect 2731 2496 2743 2499
rect 2961 2499 3019 2505
rect 2731 2468 2820 2496
rect 2731 2465 2743 2468
rect 2685 2459 2743 2465
rect 2792 2428 2820 2468
rect 2961 2465 2973 2499
rect 3007 2465 3019 2499
rect 3418 2496 3424 2508
rect 2961 2459 3019 2465
rect 3068 2468 3424 2496
rect 3068 2428 3096 2468
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 4132 2499 4190 2505
rect 4132 2465 4144 2499
rect 4178 2496 4190 2499
rect 5166 2496 5172 2508
rect 4178 2468 5172 2496
rect 4178 2465 4190 2468
rect 4132 2459 4190 2465
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 8680 2505 8708 2592
rect 9784 2508 9812 2604
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 12526 2632 12532 2644
rect 11440 2604 12532 2632
rect 11440 2508 11468 2604
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 13630 2632 13636 2644
rect 13591 2604 13636 2632
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 14550 2632 14556 2644
rect 14511 2604 14556 2632
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 15654 2632 15660 2644
rect 15615 2604 15660 2632
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 16206 2592 16212 2644
rect 16264 2632 16270 2644
rect 16301 2635 16359 2641
rect 16301 2632 16313 2635
rect 16264 2604 16313 2632
rect 16264 2592 16270 2604
rect 16301 2601 16313 2604
rect 16347 2632 16359 2635
rect 17402 2632 17408 2644
rect 16347 2604 16849 2632
rect 17363 2604 17408 2632
rect 16347 2601 16359 2604
rect 16301 2595 16359 2601
rect 11701 2567 11759 2573
rect 11701 2533 11713 2567
rect 11747 2564 11759 2567
rect 12342 2564 12348 2576
rect 11747 2536 12348 2564
rect 11747 2533 11759 2536
rect 11701 2527 11759 2533
rect 12342 2524 12348 2536
rect 12400 2524 12406 2576
rect 12618 2524 12624 2576
rect 12676 2564 12682 2576
rect 16821 2573 16849 2604
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 18414 2592 18420 2644
rect 18472 2632 18478 2644
rect 19245 2635 19303 2641
rect 19245 2632 19257 2635
rect 18472 2604 19257 2632
rect 18472 2592 18478 2604
rect 19245 2601 19257 2604
rect 19291 2601 19303 2635
rect 19245 2595 19303 2601
rect 20211 2635 20269 2641
rect 20211 2601 20223 2635
rect 20257 2632 20269 2635
rect 20622 2632 20628 2644
rect 20257 2604 20628 2632
rect 20257 2601 20269 2604
rect 20211 2595 20269 2601
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 21910 2592 21916 2644
rect 21968 2632 21974 2644
rect 22281 2635 22339 2641
rect 22281 2632 22293 2635
rect 21968 2604 22293 2632
rect 21968 2592 21974 2604
rect 22281 2601 22293 2604
rect 22327 2601 22339 2635
rect 22281 2595 22339 2601
rect 22741 2635 22799 2641
rect 22741 2601 22753 2635
rect 22787 2632 22799 2635
rect 23106 2632 23112 2644
rect 22787 2604 23112 2632
rect 22787 2601 22799 2604
rect 22741 2595 22799 2601
rect 13034 2567 13092 2573
rect 13034 2564 13046 2567
rect 12676 2536 13046 2564
rect 12676 2524 12682 2536
rect 13034 2533 13046 2536
rect 13080 2533 13092 2567
rect 13034 2527 13092 2533
rect 16806 2567 16864 2573
rect 16806 2533 16818 2567
rect 16852 2564 16864 2567
rect 17862 2564 17868 2576
rect 16852 2536 17868 2564
rect 16852 2533 16864 2536
rect 16806 2527 16864 2533
rect 17862 2524 17868 2536
rect 17920 2564 17926 2576
rect 18049 2567 18107 2573
rect 18049 2564 18061 2567
rect 17920 2536 18061 2564
rect 17920 2524 17926 2536
rect 18049 2533 18061 2536
rect 18095 2564 18107 2567
rect 18646 2567 18704 2573
rect 18646 2564 18658 2567
rect 18095 2536 18658 2564
rect 18095 2533 18107 2536
rect 18049 2527 18107 2533
rect 18646 2533 18658 2536
rect 18692 2533 18704 2567
rect 18646 2527 18704 2533
rect 20993 2567 21051 2573
rect 20993 2533 21005 2567
rect 21039 2564 21051 2567
rect 21453 2567 21511 2573
rect 21453 2564 21465 2567
rect 21039 2536 21465 2564
rect 21039 2533 21051 2536
rect 20993 2527 21051 2533
rect 21453 2533 21465 2536
rect 21499 2564 21511 2567
rect 21726 2564 21732 2576
rect 21499 2536 21732 2564
rect 21499 2533 21511 2536
rect 21453 2527 21511 2533
rect 21726 2524 21732 2536
rect 21784 2524 21790 2576
rect 8665 2499 8723 2505
rect 8665 2465 8677 2499
rect 8711 2465 8723 2499
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 8665 2459 8723 2465
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 11146 2496 11152 2508
rect 11107 2468 11152 2496
rect 11146 2456 11152 2468
rect 11204 2456 11210 2508
rect 11422 2496 11428 2508
rect 11383 2468 11428 2496
rect 11422 2456 11428 2468
rect 11480 2456 11486 2508
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 15470 2456 15476 2468
rect 15528 2496 15534 2508
rect 15933 2499 15991 2505
rect 15933 2496 15945 2499
rect 15528 2468 15945 2496
rect 15528 2456 15534 2468
rect 15933 2465 15945 2468
rect 15979 2465 15991 2499
rect 15933 2459 15991 2465
rect 19978 2456 19984 2508
rect 20036 2496 20042 2508
rect 20140 2499 20198 2505
rect 20140 2496 20152 2499
rect 20036 2468 20152 2496
rect 20036 2456 20042 2468
rect 20140 2465 20152 2468
rect 20186 2496 20198 2499
rect 20533 2499 20591 2505
rect 20533 2496 20545 2499
rect 20186 2468 20545 2496
rect 20186 2465 20198 2468
rect 20140 2459 20198 2465
rect 20533 2465 20545 2468
rect 20579 2465 20591 2499
rect 20533 2459 20591 2465
rect 2792 2400 3096 2428
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2428 3203 2431
rect 3878 2428 3884 2440
rect 3191 2400 3884 2428
rect 3191 2397 3203 2400
rect 3145 2391 3203 2397
rect 3878 2388 3884 2400
rect 3936 2388 3942 2440
rect 3970 2388 3976 2440
rect 4028 2428 4034 2440
rect 5077 2431 5135 2437
rect 5077 2428 5089 2431
rect 4028 2400 5089 2428
rect 4028 2388 4034 2400
rect 5077 2397 5089 2400
rect 5123 2428 5135 2431
rect 6273 2431 6331 2437
rect 6273 2428 6285 2431
rect 5123 2400 6285 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 6273 2397 6285 2400
rect 6319 2397 6331 2431
rect 6273 2391 6331 2397
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 7834 2428 7840 2440
rect 7055 2400 7840 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 9490 2428 9496 2440
rect 9451 2400 9496 2428
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 9600 2400 10333 2428
rect 9600 2360 9628 2400
rect 10321 2397 10333 2400
rect 10367 2428 10379 2431
rect 10689 2431 10747 2437
rect 10689 2428 10701 2431
rect 10367 2400 10701 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 10689 2397 10701 2400
rect 10735 2428 10747 2431
rect 10778 2428 10784 2440
rect 10735 2400 10784 2428
rect 10735 2397 10747 2400
rect 10689 2391 10747 2397
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 11164 2428 11192 2456
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11164 2400 11989 2428
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 12710 2428 12716 2440
rect 12671 2400 12716 2428
rect 11977 2391 12035 2397
rect 12710 2388 12716 2400
rect 12768 2428 12774 2440
rect 13909 2431 13967 2437
rect 13909 2428 13921 2431
rect 12768 2400 13921 2428
rect 12768 2388 12774 2400
rect 13909 2397 13921 2400
rect 13955 2397 13967 2431
rect 13909 2391 13967 2397
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 16482 2428 16488 2440
rect 15335 2400 16488 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 16482 2388 16488 2400
rect 16540 2388 16546 2440
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2428 17831 2431
rect 18322 2428 18328 2440
rect 17819 2400 18328 2428
rect 17819 2397 17831 2400
rect 17773 2391 17831 2397
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 21361 2431 21419 2437
rect 21361 2397 21373 2431
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 8864 2332 9628 2360
rect 21376 2360 21404 2391
rect 21450 2388 21456 2440
rect 21508 2428 21514 2440
rect 21637 2431 21695 2437
rect 21637 2428 21649 2431
rect 21508 2400 21649 2428
rect 21508 2388 21514 2400
rect 21637 2397 21649 2400
rect 21683 2397 21695 2431
rect 22756 2428 22784 2595
rect 23106 2592 23112 2604
rect 23164 2592 23170 2644
rect 23382 2592 23388 2644
rect 23440 2632 23446 2644
rect 23753 2635 23811 2641
rect 23753 2632 23765 2635
rect 23440 2604 23765 2632
rect 23440 2592 23446 2604
rect 23753 2601 23765 2604
rect 23799 2601 23811 2635
rect 24118 2632 24124 2644
rect 24079 2604 24124 2632
rect 23753 2595 23811 2601
rect 24118 2592 24124 2604
rect 24176 2592 24182 2644
rect 25314 2592 25320 2644
rect 25372 2632 25378 2644
rect 25409 2635 25467 2641
rect 25409 2632 25421 2635
rect 25372 2604 25421 2632
rect 25372 2592 25378 2604
rect 25409 2601 25421 2604
rect 25455 2601 25467 2635
rect 25409 2595 25467 2601
rect 23477 2567 23535 2573
rect 23477 2533 23489 2567
rect 23523 2564 23535 2567
rect 23658 2564 23664 2576
rect 23523 2536 23664 2564
rect 23523 2533 23535 2536
rect 23477 2527 23535 2533
rect 22833 2499 22891 2505
rect 22833 2465 22845 2499
rect 22879 2496 22891 2499
rect 23492 2496 23520 2527
rect 23658 2524 23664 2536
rect 23716 2524 23722 2576
rect 24029 2499 24087 2505
rect 24029 2496 24041 2499
rect 22879 2468 23520 2496
rect 23952 2468 24041 2496
rect 22879 2465 22891 2468
rect 22833 2459 22891 2465
rect 21637 2391 21695 2397
rect 21744 2400 22784 2428
rect 23952 2428 23980 2468
rect 24029 2465 24041 2468
rect 24075 2465 24087 2499
rect 24029 2459 24087 2465
rect 24581 2499 24639 2505
rect 24581 2465 24593 2499
rect 24627 2496 24639 2499
rect 25332 2496 25360 2592
rect 24627 2468 25360 2496
rect 25660 2499 25718 2505
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 25660 2465 25672 2499
rect 25706 2496 25718 2499
rect 26142 2496 26148 2508
rect 25706 2468 26148 2496
rect 25706 2465 25718 2468
rect 25660 2459 25718 2465
rect 26142 2456 26148 2468
rect 26200 2456 26206 2508
rect 25041 2431 25099 2437
rect 25041 2428 25053 2431
rect 23952 2400 25053 2428
rect 21744 2360 21772 2400
rect 21376 2332 21772 2360
rect 8864 2304 8892 2332
rect 22738 2320 22744 2372
rect 22796 2360 22802 2372
rect 23952 2360 23980 2400
rect 25041 2397 25053 2400
rect 25087 2397 25099 2431
rect 25041 2391 25099 2397
rect 22796 2332 23980 2360
rect 22796 2320 22802 2332
rect 1535 2295 1593 2301
rect 1535 2261 1547 2295
rect 1581 2292 1593 2295
rect 2130 2292 2136 2304
rect 1581 2264 2136 2292
rect 1581 2261 1593 2264
rect 1535 2255 1593 2261
rect 2130 2252 2136 2264
rect 2188 2252 2194 2304
rect 4203 2295 4261 2301
rect 4203 2261 4215 2295
rect 4249 2292 4261 2295
rect 5442 2292 5448 2304
rect 4249 2264 5448 2292
rect 4249 2261 4261 2264
rect 4203 2255 4261 2261
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 8846 2292 8852 2304
rect 8807 2264 8852 2292
rect 8846 2252 8852 2264
rect 8904 2252 8910 2304
rect 9950 2292 9956 2304
rect 9911 2264 9956 2292
rect 9950 2252 9956 2264
rect 10008 2252 10014 2304
rect 10042 2252 10048 2304
rect 10100 2292 10106 2304
rect 12345 2295 12403 2301
rect 12345 2292 12357 2295
rect 10100 2264 12357 2292
rect 10100 2252 10106 2264
rect 12345 2261 12357 2264
rect 12391 2292 12403 2295
rect 12618 2292 12624 2304
rect 12391 2264 12624 2292
rect 12391 2261 12403 2264
rect 12345 2255 12403 2261
rect 12618 2252 12624 2264
rect 12676 2252 12682 2304
rect 21634 2252 21640 2304
rect 21692 2292 21698 2304
rect 23017 2295 23075 2301
rect 23017 2292 23029 2295
rect 21692 2264 23029 2292
rect 21692 2252 21698 2264
rect 23017 2261 23029 2264
rect 23063 2261 23075 2295
rect 23017 2255 23075 2261
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25731 2295 25789 2301
rect 25731 2292 25743 2295
rect 25188 2264 25743 2292
rect 25188 2252 25194 2264
rect 25731 2261 25743 2264
rect 25777 2261 25789 2295
rect 26142 2292 26148 2304
rect 26103 2264 26148 2292
rect 25731 2255 25789 2261
rect 26142 2252 26148 2264
rect 26200 2252 26206 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 20254 2048 20260 2100
rect 20312 2088 20318 2100
rect 22646 2088 22652 2100
rect 20312 2060 22652 2088
rect 20312 2048 20318 2060
rect 22646 2048 22652 2060
rect 22704 2048 22710 2100
rect 14458 1980 14464 2032
rect 14516 2020 14522 2032
rect 14918 2020 14924 2032
rect 14516 1992 14924 2020
rect 14516 1980 14522 1992
rect 14918 1980 14924 1992
rect 14976 1980 14982 2032
rect 24578 1980 24584 2032
rect 24636 2020 24642 2032
rect 25590 2020 25596 2032
rect 24636 1992 25596 2020
rect 24636 1980 24642 1992
rect 25590 1980 25596 1992
rect 25648 1980 25654 2032
rect 16850 552 16856 604
rect 16908 592 16914 604
rect 18046 592 18052 604
rect 16908 564 18052 592
rect 16908 552 16914 564
rect 18046 552 18052 564
rect 18104 552 18110 604
<< via1 >>
rect 18328 26596 18380 26648
rect 23480 26596 23532 26648
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 17132 24395 17184 24404
rect 17132 24361 17141 24395
rect 17141 24361 17175 24395
rect 17175 24361 17184 24395
rect 17132 24352 17184 24361
rect 18236 24395 18288 24404
rect 18236 24361 18245 24395
rect 18245 24361 18279 24395
rect 18279 24361 18288 24395
rect 18236 24352 18288 24361
rect 10692 24259 10744 24268
rect 10692 24225 10710 24259
rect 10710 24225 10744 24259
rect 10692 24216 10744 24225
rect 11612 24259 11664 24268
rect 11612 24225 11656 24259
rect 11656 24225 11664 24259
rect 11612 24216 11664 24225
rect 17316 24216 17368 24268
rect 18696 24216 18748 24268
rect 10048 24012 10100 24064
rect 11888 24012 11940 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 10692 23851 10744 23860
rect 10692 23817 10701 23851
rect 10701 23817 10735 23851
rect 10735 23817 10744 23851
rect 10692 23808 10744 23817
rect 14556 23851 14608 23860
rect 14556 23817 14565 23851
rect 14565 23817 14599 23851
rect 14599 23817 14608 23851
rect 14556 23808 14608 23817
rect 16212 23851 16264 23860
rect 16212 23817 16221 23851
rect 16221 23817 16255 23851
rect 16255 23817 16264 23851
rect 16212 23808 16264 23817
rect 18236 23851 18288 23860
rect 18236 23817 18245 23851
rect 18245 23817 18279 23851
rect 18279 23817 18288 23851
rect 18236 23808 18288 23817
rect 20352 23851 20404 23860
rect 20352 23817 20361 23851
rect 20361 23817 20395 23851
rect 20395 23817 20404 23851
rect 20352 23808 20404 23817
rect 21456 23851 21508 23860
rect 21456 23817 21465 23851
rect 21465 23817 21499 23851
rect 21499 23817 21508 23851
rect 21456 23808 21508 23817
rect 22560 23851 22612 23860
rect 22560 23817 22569 23851
rect 22569 23817 22603 23851
rect 22603 23817 22612 23851
rect 22560 23808 22612 23817
rect 24768 23851 24820 23860
rect 24768 23817 24777 23851
rect 24777 23817 24811 23851
rect 24811 23817 24820 23851
rect 24768 23808 24820 23817
rect 8944 23647 8996 23656
rect 8944 23613 8953 23647
rect 8953 23613 8987 23647
rect 8987 23613 8996 23647
rect 8944 23604 8996 23613
rect 11152 23647 11204 23656
rect 11152 23613 11170 23647
rect 11170 23613 11204 23647
rect 11152 23604 11204 23613
rect 12440 23647 12492 23656
rect 12440 23613 12484 23647
rect 12484 23613 12492 23647
rect 12440 23604 12492 23613
rect 13820 23604 13872 23656
rect 16028 23647 16080 23656
rect 16028 23613 16037 23647
rect 16037 23613 16071 23647
rect 16071 23613 16080 23647
rect 16028 23604 16080 23613
rect 18144 23604 18196 23656
rect 21272 23647 21324 23656
rect 2044 23511 2096 23520
rect 2044 23477 2053 23511
rect 2053 23477 2087 23511
rect 2087 23477 2096 23511
rect 2044 23468 2096 23477
rect 9128 23511 9180 23520
rect 9128 23477 9137 23511
rect 9137 23477 9171 23511
rect 9171 23477 9180 23511
rect 9128 23468 9180 23477
rect 9956 23511 10008 23520
rect 9956 23477 9965 23511
rect 9965 23477 9999 23511
rect 9999 23477 10008 23511
rect 9956 23468 10008 23477
rect 10968 23468 11020 23520
rect 11612 23511 11664 23520
rect 11612 23477 11621 23511
rect 11621 23477 11655 23511
rect 11655 23477 11664 23511
rect 11612 23468 11664 23477
rect 13360 23468 13412 23520
rect 17316 23468 17368 23520
rect 18696 23511 18748 23520
rect 18696 23477 18705 23511
rect 18705 23477 18739 23511
rect 18739 23477 18748 23511
rect 18696 23468 18748 23477
rect 21272 23613 21281 23647
rect 21281 23613 21315 23647
rect 21315 23613 21324 23647
rect 21272 23604 21324 23613
rect 22192 23604 22244 23656
rect 24584 23647 24636 23656
rect 24584 23613 24593 23647
rect 24593 23613 24627 23647
rect 24627 23613 24636 23647
rect 24584 23604 24636 23613
rect 21272 23468 21324 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1400 23264 1452 23316
rect 11152 23307 11204 23316
rect 11152 23273 11161 23307
rect 11161 23273 11195 23307
rect 11195 23273 11204 23307
rect 11152 23264 11204 23273
rect 13728 23264 13780 23316
rect 18328 23264 18380 23316
rect 24676 23264 24728 23316
rect 9864 23239 9916 23248
rect 9864 23205 9873 23239
rect 9873 23205 9907 23239
rect 9907 23205 9916 23239
rect 9864 23196 9916 23205
rect 1676 23128 1728 23180
rect 7288 23171 7340 23180
rect 7288 23137 7332 23171
rect 7332 23137 7340 23171
rect 7288 23128 7340 23137
rect 8576 23171 8628 23180
rect 8576 23137 8620 23171
rect 8620 23137 8628 23171
rect 8576 23128 8628 23137
rect 11336 23171 11388 23180
rect 11336 23137 11354 23171
rect 11354 23137 11388 23171
rect 11336 23128 11388 23137
rect 12256 23171 12308 23180
rect 12256 23137 12300 23171
rect 12300 23137 12308 23171
rect 12256 23128 12308 23137
rect 13544 23171 13596 23180
rect 13544 23137 13588 23171
rect 13588 23137 13596 23171
rect 13544 23128 13596 23137
rect 15568 23171 15620 23180
rect 15568 23137 15586 23171
rect 15586 23137 15620 23171
rect 15568 23128 15620 23137
rect 16764 23171 16816 23180
rect 16764 23137 16808 23171
rect 16808 23137 16816 23171
rect 18052 23171 18104 23180
rect 16764 23128 16816 23137
rect 18052 23137 18061 23171
rect 18061 23137 18095 23171
rect 18095 23137 18104 23171
rect 18052 23128 18104 23137
rect 24124 23128 24176 23180
rect 7472 23060 7524 23112
rect 9772 23103 9824 23112
rect 9772 23069 9781 23103
rect 9781 23069 9815 23103
rect 9815 23069 9824 23103
rect 9772 23060 9824 23069
rect 10140 23103 10192 23112
rect 10140 23069 10149 23103
rect 10149 23069 10183 23103
rect 10183 23069 10192 23103
rect 10140 23060 10192 23069
rect 7656 22924 7708 22976
rect 8760 22924 8812 22976
rect 11152 22924 11204 22976
rect 12348 22924 12400 22976
rect 15936 22924 15988 22976
rect 17408 22924 17460 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1492 22720 1544 22772
rect 6276 22763 6328 22772
rect 6276 22729 6285 22763
rect 6285 22729 6319 22763
rect 6319 22729 6328 22763
rect 6276 22720 6328 22729
rect 8576 22763 8628 22772
rect 8576 22729 8585 22763
rect 8585 22729 8619 22763
rect 8619 22729 8628 22763
rect 8576 22720 8628 22729
rect 9588 22720 9640 22772
rect 9772 22720 9824 22772
rect 13544 22720 13596 22772
rect 15568 22763 15620 22772
rect 15568 22729 15577 22763
rect 15577 22729 15611 22763
rect 15611 22729 15620 22763
rect 15568 22720 15620 22729
rect 16764 22763 16816 22772
rect 16764 22729 16773 22763
rect 16773 22729 16807 22763
rect 16807 22729 16816 22763
rect 16764 22720 16816 22729
rect 7288 22652 7340 22704
rect 7840 22652 7892 22704
rect 13820 22652 13872 22704
rect 18052 22652 18104 22704
rect 7472 22584 7524 22636
rect 7564 22584 7616 22636
rect 9680 22584 9732 22636
rect 10140 22584 10192 22636
rect 5540 22516 5592 22568
rect 6276 22516 6328 22568
rect 6736 22448 6788 22500
rect 2228 22380 2280 22432
rect 10784 22559 10836 22568
rect 12256 22584 12308 22636
rect 10784 22525 10828 22559
rect 10828 22525 10836 22559
rect 10784 22516 10836 22525
rect 12440 22559 12492 22568
rect 12440 22525 12449 22559
rect 12449 22525 12483 22559
rect 12483 22525 12492 22559
rect 12440 22516 12492 22525
rect 14464 22516 14516 22568
rect 16672 22516 16724 22568
rect 9312 22491 9364 22500
rect 9312 22457 9321 22491
rect 9321 22457 9355 22491
rect 9355 22457 9364 22491
rect 9312 22448 9364 22457
rect 7748 22380 7800 22432
rect 8668 22380 8720 22432
rect 12808 22448 12860 22500
rect 14004 22491 14056 22500
rect 14004 22457 14013 22491
rect 14013 22457 14047 22491
rect 14047 22457 14056 22491
rect 14004 22448 14056 22457
rect 9864 22380 9916 22432
rect 10692 22380 10744 22432
rect 11336 22423 11388 22432
rect 11336 22389 11345 22423
rect 11345 22389 11379 22423
rect 11379 22389 11388 22423
rect 11336 22380 11388 22389
rect 13084 22380 13136 22432
rect 15660 22423 15712 22432
rect 15660 22389 15669 22423
rect 15669 22389 15703 22423
rect 15703 22389 15712 22423
rect 15660 22380 15712 22389
rect 24124 22380 24176 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 7472 22176 7524 22228
rect 8760 22219 8812 22228
rect 5172 22151 5224 22160
rect 5172 22117 5181 22151
rect 5181 22117 5215 22151
rect 5215 22117 5224 22151
rect 5172 22108 5224 22117
rect 6920 22108 6972 22160
rect 6184 22083 6236 22092
rect 6184 22049 6228 22083
rect 6228 22049 6236 22083
rect 8760 22185 8769 22219
rect 8769 22185 8803 22219
rect 8803 22185 8812 22219
rect 8760 22176 8812 22185
rect 11152 22176 11204 22228
rect 12348 22219 12400 22228
rect 12348 22185 12357 22219
rect 12357 22185 12391 22219
rect 12391 22185 12400 22219
rect 12348 22176 12400 22185
rect 10140 22151 10192 22160
rect 10140 22117 10149 22151
rect 10149 22117 10183 22151
rect 10183 22117 10192 22151
rect 10140 22108 10192 22117
rect 13636 22108 13688 22160
rect 15568 22108 15620 22160
rect 6184 22040 6236 22049
rect 9128 22040 9180 22092
rect 11520 22083 11572 22092
rect 11520 22049 11564 22083
rect 11564 22049 11572 22083
rect 11520 22040 11572 22049
rect 1676 22015 1728 22024
rect 1676 21981 1685 22015
rect 1685 21981 1719 22015
rect 1719 21981 1728 22015
rect 1676 21972 1728 21981
rect 5540 21972 5592 22024
rect 7564 22015 7616 22024
rect 7564 21981 7573 22015
rect 7573 21981 7607 22015
rect 7607 21981 7616 22015
rect 7564 21972 7616 21981
rect 9496 21972 9548 22024
rect 10692 21972 10744 22024
rect 13452 22015 13504 22024
rect 13452 21981 13461 22015
rect 13461 21981 13495 22015
rect 13495 21981 13504 22015
rect 13452 21972 13504 21981
rect 16948 21972 17000 22024
rect 8024 21904 8076 21956
rect 9680 21904 9732 21956
rect 15752 21904 15804 21956
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 12900 21836 12952 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 6184 21632 6236 21684
rect 7288 21632 7340 21684
rect 9680 21632 9732 21684
rect 9864 21632 9916 21684
rect 10692 21632 10744 21684
rect 11520 21675 11572 21684
rect 11520 21641 11529 21675
rect 11529 21641 11563 21675
rect 11563 21641 11572 21675
rect 11520 21632 11572 21641
rect 13636 21632 13688 21684
rect 15844 21632 15896 21684
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 8760 21564 8812 21616
rect 7564 21539 7616 21548
rect 7564 21505 7573 21539
rect 7573 21505 7607 21539
rect 7607 21505 7616 21539
rect 7564 21496 7616 21505
rect 13912 21564 13964 21616
rect 9128 21539 9180 21548
rect 9128 21505 9137 21539
rect 9137 21505 9171 21539
rect 9171 21505 9180 21539
rect 9128 21496 9180 21505
rect 9864 21496 9916 21548
rect 10048 21496 10100 21548
rect 11152 21496 11204 21548
rect 12808 21539 12860 21548
rect 12808 21505 12817 21539
rect 12817 21505 12851 21539
rect 12851 21505 12860 21539
rect 12808 21496 12860 21505
rect 13452 21539 13504 21548
rect 13452 21505 13461 21539
rect 13461 21505 13495 21539
rect 13495 21505 13504 21539
rect 14372 21539 14424 21548
rect 13452 21496 13504 21505
rect 14372 21505 14381 21539
rect 14381 21505 14415 21539
rect 14415 21505 14424 21539
rect 14372 21496 14424 21505
rect 2044 21471 2096 21480
rect 2044 21437 2053 21471
rect 2053 21437 2087 21471
rect 2087 21437 2096 21471
rect 2044 21428 2096 21437
rect 6276 21403 6328 21412
rect 6276 21369 6285 21403
rect 6285 21369 6319 21403
rect 6319 21369 6328 21403
rect 6276 21360 6328 21369
rect 7288 21403 7340 21412
rect 7288 21369 7297 21403
rect 7297 21369 7331 21403
rect 7331 21369 7340 21403
rect 7288 21360 7340 21369
rect 7380 21403 7432 21412
rect 7380 21369 7389 21403
rect 7389 21369 7423 21403
rect 7423 21369 7432 21403
rect 7380 21360 7432 21369
rect 4436 21292 4488 21344
rect 5080 21335 5132 21344
rect 5080 21301 5089 21335
rect 5089 21301 5123 21335
rect 5123 21301 5132 21335
rect 5080 21292 5132 21301
rect 6000 21292 6052 21344
rect 6828 21292 6880 21344
rect 8668 21335 8720 21344
rect 8668 21301 8677 21335
rect 8677 21301 8711 21335
rect 8711 21301 8720 21335
rect 8668 21292 8720 21301
rect 10048 21292 10100 21344
rect 12900 21403 12952 21412
rect 12900 21369 12909 21403
rect 12909 21369 12943 21403
rect 12943 21369 12952 21403
rect 12900 21360 12952 21369
rect 13544 21360 13596 21412
rect 15016 21403 15068 21412
rect 14188 21335 14240 21344
rect 14188 21301 14197 21335
rect 14197 21301 14231 21335
rect 14231 21301 14240 21335
rect 15016 21369 15025 21403
rect 15025 21369 15059 21403
rect 15059 21369 15068 21403
rect 15016 21360 15068 21369
rect 16120 21564 16172 21616
rect 15936 21539 15988 21548
rect 15936 21505 15945 21539
rect 15945 21505 15979 21539
rect 15979 21505 15988 21539
rect 15936 21496 15988 21505
rect 18144 21471 18196 21480
rect 18144 21437 18162 21471
rect 18162 21437 18196 21471
rect 18144 21428 18196 21437
rect 16764 21360 16816 21412
rect 16948 21403 17000 21412
rect 16948 21369 16957 21403
rect 16957 21369 16991 21403
rect 16991 21369 17000 21403
rect 16948 21360 17000 21369
rect 17868 21360 17920 21412
rect 14188 21292 14240 21301
rect 15568 21292 15620 21344
rect 16856 21292 16908 21344
rect 17500 21292 17552 21344
rect 18788 21292 18840 21344
rect 24216 21292 24268 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 5264 21131 5316 21140
rect 5264 21097 5273 21131
rect 5273 21097 5307 21131
rect 5307 21097 5316 21131
rect 5264 21088 5316 21097
rect 7380 21131 7432 21140
rect 7380 21097 7389 21131
rect 7389 21097 7423 21131
rect 7423 21097 7432 21131
rect 7380 21088 7432 21097
rect 8024 21131 8076 21140
rect 8024 21097 8033 21131
rect 8033 21097 8067 21131
rect 8067 21097 8076 21131
rect 8024 21088 8076 21097
rect 9772 21088 9824 21140
rect 15844 21088 15896 21140
rect 6644 21020 6696 21072
rect 9496 21063 9548 21072
rect 9496 21029 9505 21063
rect 9505 21029 9539 21063
rect 9539 21029 9548 21063
rect 9496 21020 9548 21029
rect 10692 21020 10744 21072
rect 13912 21020 13964 21072
rect 14372 21063 14424 21072
rect 14372 21029 14381 21063
rect 14381 21029 14415 21063
rect 14415 21029 14424 21063
rect 14372 21020 14424 21029
rect 15660 21020 15712 21072
rect 16764 21088 16816 21140
rect 17500 21063 17552 21072
rect 17500 21029 17509 21063
rect 17509 21029 17543 21063
rect 17543 21029 17552 21063
rect 17500 21020 17552 21029
rect 4712 20952 4764 21004
rect 5080 20952 5132 21004
rect 6092 20952 6144 21004
rect 8852 20952 8904 21004
rect 11152 20995 11204 21004
rect 11152 20961 11161 20995
rect 11161 20961 11195 20995
rect 11195 20961 11204 20995
rect 12072 20995 12124 21004
rect 11152 20952 11204 20961
rect 12072 20961 12081 20995
rect 12081 20961 12115 20995
rect 12115 20961 12124 20995
rect 12072 20952 12124 20961
rect 12624 20995 12676 21004
rect 12624 20961 12633 20995
rect 12633 20961 12667 20995
rect 12667 20961 12676 20995
rect 12624 20952 12676 20961
rect 5632 20884 5684 20936
rect 10692 20884 10744 20936
rect 13268 20927 13320 20936
rect 13268 20893 13277 20927
rect 13277 20893 13311 20927
rect 13311 20893 13320 20927
rect 13268 20884 13320 20893
rect 13728 20927 13780 20936
rect 13728 20893 13737 20927
rect 13737 20893 13771 20927
rect 13771 20893 13780 20927
rect 13728 20884 13780 20893
rect 16120 20884 16172 20936
rect 4160 20748 4212 20800
rect 6552 20748 6604 20800
rect 7012 20748 7064 20800
rect 9036 20791 9088 20800
rect 9036 20757 9045 20791
rect 9045 20757 9079 20791
rect 9079 20757 9088 20791
rect 9036 20748 9088 20757
rect 10048 20748 10100 20800
rect 15752 20791 15804 20800
rect 15752 20757 15761 20791
rect 15761 20757 15795 20791
rect 15795 20757 15804 20791
rect 15752 20748 15804 20757
rect 16580 20748 16632 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2412 20476 2464 20528
rect 6368 20544 6420 20596
rect 7748 20587 7800 20596
rect 7748 20553 7757 20587
rect 7757 20553 7791 20587
rect 7791 20553 7800 20587
rect 7748 20544 7800 20553
rect 8852 20544 8904 20596
rect 9956 20587 10008 20596
rect 9956 20553 9965 20587
rect 9965 20553 9999 20587
rect 9999 20553 10008 20587
rect 9956 20544 10008 20553
rect 10784 20544 10836 20596
rect 12072 20587 12124 20596
rect 12072 20553 12081 20587
rect 12081 20553 12115 20587
rect 12115 20553 12124 20587
rect 12072 20544 12124 20553
rect 12624 20587 12676 20596
rect 12624 20553 12633 20587
rect 12633 20553 12667 20587
rect 12667 20553 12676 20587
rect 12624 20544 12676 20553
rect 14188 20587 14240 20596
rect 14188 20553 14197 20587
rect 14197 20553 14231 20587
rect 14231 20553 14240 20587
rect 14188 20544 14240 20553
rect 15660 20544 15712 20596
rect 16764 20544 16816 20596
rect 17500 20544 17552 20596
rect 17960 20544 18012 20596
rect 6092 20476 6144 20528
rect 6828 20476 6880 20528
rect 9036 20408 9088 20460
rect 9128 20451 9180 20460
rect 9128 20417 9137 20451
rect 9137 20417 9171 20451
rect 9171 20417 9180 20451
rect 9128 20408 9180 20417
rect 10508 20451 10560 20460
rect 10508 20417 10517 20451
rect 10517 20417 10551 20451
rect 10551 20417 10560 20451
rect 10508 20408 10560 20417
rect 10876 20408 10928 20460
rect 13268 20451 13320 20460
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 15568 20451 15620 20460
rect 15568 20417 15577 20451
rect 15577 20417 15611 20451
rect 15611 20417 15620 20451
rect 15568 20408 15620 20417
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 3792 20383 3844 20392
rect 3792 20349 3836 20383
rect 3836 20349 3844 20383
rect 3792 20340 3844 20349
rect 4896 20340 4948 20392
rect 5264 20340 5316 20392
rect 6092 20340 6144 20392
rect 7012 20340 7064 20392
rect 14740 20340 14792 20392
rect 5908 20315 5960 20324
rect 5908 20281 5917 20315
rect 5917 20281 5951 20315
rect 5951 20281 5960 20315
rect 5908 20272 5960 20281
rect 8760 20315 8812 20324
rect 8760 20281 8769 20315
rect 8769 20281 8803 20315
rect 8803 20281 8812 20315
rect 8760 20272 8812 20281
rect 10048 20272 10100 20324
rect 15752 20272 15804 20324
rect 1952 20204 2004 20256
rect 3148 20204 3200 20256
rect 3884 20204 3936 20256
rect 4712 20247 4764 20256
rect 4712 20213 4721 20247
rect 4721 20213 4755 20247
rect 4755 20213 4764 20247
rect 4712 20204 4764 20213
rect 5448 20204 5500 20256
rect 6644 20247 6696 20256
rect 6644 20213 6653 20247
rect 6653 20213 6687 20247
rect 6687 20213 6696 20247
rect 6644 20204 6696 20213
rect 10692 20204 10744 20256
rect 13452 20204 13504 20256
rect 14464 20247 14516 20256
rect 14464 20213 14473 20247
rect 14473 20213 14507 20247
rect 14507 20213 14516 20247
rect 14464 20204 14516 20213
rect 14832 20204 14884 20256
rect 16488 20272 16540 20324
rect 18696 20340 18748 20392
rect 19064 20383 19116 20392
rect 19064 20349 19108 20383
rect 19108 20349 19116 20383
rect 19064 20340 19116 20349
rect 16580 20204 16632 20256
rect 18512 20247 18564 20256
rect 18512 20213 18521 20247
rect 18521 20213 18555 20247
rect 18555 20213 18564 20247
rect 18512 20204 18564 20213
rect 19984 20204 20036 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 6920 20000 6972 20052
rect 9036 20000 9088 20052
rect 10692 20000 10744 20052
rect 13820 20000 13872 20052
rect 15844 20043 15896 20052
rect 15844 20009 15853 20043
rect 15853 20009 15887 20043
rect 15887 20009 15896 20043
rect 15844 20000 15896 20009
rect 5540 19975 5592 19984
rect 5540 19941 5549 19975
rect 5549 19941 5583 19975
rect 5583 19941 5592 19975
rect 5540 19932 5592 19941
rect 6644 19932 6696 19984
rect 9956 19932 10008 19984
rect 13452 19932 13504 19984
rect 16212 19975 16264 19984
rect 16212 19941 16221 19975
rect 16221 19941 16255 19975
rect 16255 19941 16264 19975
rect 16212 19932 16264 19941
rect 16856 19932 16908 19984
rect 17868 19932 17920 19984
rect 1860 19864 1912 19916
rect 3056 19864 3108 19916
rect 4160 19864 4212 19916
rect 5080 19907 5132 19916
rect 5080 19873 5089 19907
rect 5089 19873 5123 19907
rect 5123 19873 5132 19907
rect 5080 19864 5132 19873
rect 5264 19907 5316 19916
rect 5264 19873 5273 19907
rect 5273 19873 5307 19907
rect 5307 19873 5316 19907
rect 5264 19864 5316 19873
rect 9404 19864 9456 19916
rect 9680 19907 9732 19916
rect 9680 19873 9689 19907
rect 9689 19873 9723 19907
rect 9723 19873 9732 19907
rect 9680 19864 9732 19873
rect 6184 19796 6236 19848
rect 8760 19796 8812 19848
rect 10784 19864 10836 19916
rect 11980 19864 12032 19916
rect 13912 19864 13964 19916
rect 14464 19864 14516 19916
rect 19248 19907 19300 19916
rect 19248 19873 19266 19907
rect 19266 19873 19300 19907
rect 19248 19864 19300 19873
rect 12440 19796 12492 19848
rect 16120 19839 16172 19848
rect 16120 19805 16129 19839
rect 16129 19805 16163 19839
rect 16163 19805 16172 19839
rect 16120 19796 16172 19805
rect 17684 19839 17736 19848
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 17776 19796 17828 19848
rect 16672 19771 16724 19780
rect 16672 19737 16681 19771
rect 16681 19737 16715 19771
rect 16715 19737 16724 19771
rect 16672 19728 16724 19737
rect 2596 19660 2648 19712
rect 3516 19660 3568 19712
rect 7748 19703 7800 19712
rect 7748 19669 7757 19703
rect 7757 19669 7791 19703
rect 7791 19669 7800 19703
rect 7748 19660 7800 19669
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 17960 19660 18012 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 3056 19456 3108 19508
rect 4620 19456 4672 19508
rect 5080 19456 5132 19508
rect 10048 19456 10100 19508
rect 16212 19499 16264 19508
rect 16212 19465 16221 19499
rect 16221 19465 16255 19499
rect 16255 19465 16264 19499
rect 16212 19456 16264 19465
rect 17868 19456 17920 19508
rect 24768 19499 24820 19508
rect 24768 19465 24777 19499
rect 24777 19465 24811 19499
rect 24811 19465 24820 19499
rect 24768 19456 24820 19465
rect 9680 19388 9732 19440
rect 2320 19320 2372 19372
rect 6184 19320 6236 19372
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 2136 19116 2188 19168
rect 3608 19295 3660 19304
rect 3608 19261 3617 19295
rect 3617 19261 3651 19295
rect 3651 19261 3660 19295
rect 3608 19252 3660 19261
rect 5172 19295 5224 19304
rect 5172 19261 5181 19295
rect 5181 19261 5215 19295
rect 5215 19261 5224 19295
rect 5172 19252 5224 19261
rect 5264 19252 5316 19304
rect 5816 19252 5868 19304
rect 9404 19320 9456 19372
rect 12440 19320 12492 19372
rect 14740 19388 14792 19440
rect 7748 19295 7800 19304
rect 7748 19261 7757 19295
rect 7757 19261 7791 19295
rect 7791 19261 7800 19295
rect 7748 19252 7800 19261
rect 8668 19295 8720 19304
rect 8668 19261 8677 19295
rect 8677 19261 8711 19295
rect 8711 19261 8720 19295
rect 8668 19252 8720 19261
rect 9496 19295 9548 19304
rect 9496 19261 9505 19295
rect 9505 19261 9539 19295
rect 9539 19261 9548 19295
rect 9496 19252 9548 19261
rect 3240 19116 3292 19168
rect 3884 19159 3936 19168
rect 3884 19125 3893 19159
rect 3893 19125 3927 19159
rect 3927 19125 3936 19159
rect 3884 19116 3936 19125
rect 6184 19116 6236 19168
rect 6644 19116 6696 19168
rect 9312 19159 9364 19168
rect 9312 19125 9321 19159
rect 9321 19125 9355 19159
rect 9355 19125 9364 19159
rect 9312 19116 9364 19125
rect 9956 19184 10008 19236
rect 12532 19295 12584 19304
rect 12532 19261 12541 19295
rect 12541 19261 12575 19295
rect 12575 19261 12584 19295
rect 12532 19252 12584 19261
rect 13636 19252 13688 19304
rect 14372 19320 14424 19372
rect 16120 19320 16172 19372
rect 14740 19252 14792 19304
rect 18328 19320 18380 19372
rect 19248 19320 19300 19372
rect 10140 19116 10192 19168
rect 11152 19159 11204 19168
rect 11152 19125 11161 19159
rect 11161 19125 11195 19159
rect 11195 19125 11204 19159
rect 11152 19116 11204 19125
rect 11428 19116 11480 19168
rect 11980 19116 12032 19168
rect 13452 19116 13504 19168
rect 17776 19252 17828 19304
rect 18052 19295 18104 19304
rect 18052 19261 18096 19295
rect 18096 19261 18104 19295
rect 18052 19252 18104 19261
rect 19064 19295 19116 19304
rect 19064 19261 19073 19295
rect 19073 19261 19107 19295
rect 19107 19261 19116 19295
rect 19064 19252 19116 19261
rect 19892 19295 19944 19304
rect 19892 19261 19901 19295
rect 19901 19261 19935 19295
rect 19935 19261 19944 19295
rect 19892 19252 19944 19261
rect 24584 19295 24636 19304
rect 24584 19261 24593 19295
rect 24593 19261 24627 19295
rect 24627 19261 24636 19295
rect 24584 19252 24636 19261
rect 17684 19184 17736 19236
rect 19340 19184 19392 19236
rect 17224 19159 17276 19168
rect 17224 19125 17233 19159
rect 17233 19125 17267 19159
rect 17267 19125 17276 19159
rect 17224 19116 17276 19125
rect 17960 19116 18012 19168
rect 19248 19159 19300 19168
rect 19248 19125 19257 19159
rect 19257 19125 19291 19159
rect 19291 19125 19300 19159
rect 19248 19116 19300 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 4160 18912 4212 18964
rect 5264 18912 5316 18964
rect 9496 18955 9548 18964
rect 9496 18921 9505 18955
rect 9505 18921 9539 18955
rect 9539 18921 9548 18955
rect 9496 18912 9548 18921
rect 11244 18955 11296 18964
rect 6092 18887 6144 18896
rect 6092 18853 6101 18887
rect 6101 18853 6135 18887
rect 6135 18853 6144 18887
rect 6092 18844 6144 18853
rect 8944 18844 8996 18896
rect 9312 18844 9364 18896
rect 9956 18887 10008 18896
rect 9956 18853 9965 18887
rect 9965 18853 9999 18887
rect 9999 18853 10008 18887
rect 9956 18844 10008 18853
rect 11244 18921 11253 18955
rect 11253 18921 11287 18955
rect 11287 18921 11296 18955
rect 11244 18912 11296 18921
rect 12624 18912 12676 18964
rect 16488 18912 16540 18964
rect 17132 18955 17184 18964
rect 17132 18921 17141 18955
rect 17141 18921 17175 18955
rect 17175 18921 17184 18955
rect 17132 18912 17184 18921
rect 17684 18912 17736 18964
rect 24676 18912 24728 18964
rect 10324 18887 10376 18896
rect 10324 18853 10333 18887
rect 10333 18853 10367 18887
rect 10367 18853 10376 18887
rect 10876 18887 10928 18896
rect 10324 18844 10376 18853
rect 10876 18853 10885 18887
rect 10885 18853 10919 18887
rect 10919 18853 10928 18887
rect 10876 18844 10928 18853
rect 13452 18844 13504 18896
rect 15568 18844 15620 18896
rect 16028 18844 16080 18896
rect 17868 18844 17920 18896
rect 2228 18776 2280 18828
rect 3148 18776 3200 18828
rect 2688 18708 2740 18760
rect 3884 18708 3936 18760
rect 5540 18776 5592 18828
rect 5816 18819 5868 18828
rect 5816 18785 5825 18819
rect 5825 18785 5859 18819
rect 5859 18785 5868 18819
rect 5816 18776 5868 18785
rect 7012 18819 7064 18828
rect 7012 18785 7021 18819
rect 7021 18785 7055 18819
rect 7055 18785 7064 18819
rect 7012 18776 7064 18785
rect 7748 18776 7800 18828
rect 8668 18819 8720 18828
rect 8668 18785 8686 18819
rect 8686 18785 8720 18819
rect 8668 18776 8720 18785
rect 11796 18819 11848 18828
rect 11796 18785 11814 18819
rect 11814 18785 11848 18819
rect 11796 18776 11848 18785
rect 13544 18776 13596 18828
rect 17040 18819 17092 18828
rect 17040 18785 17049 18819
rect 17049 18785 17083 18819
rect 17083 18785 17092 18819
rect 17040 18776 17092 18785
rect 17776 18776 17828 18828
rect 18696 18819 18748 18828
rect 18696 18785 18714 18819
rect 18714 18785 18748 18819
rect 18696 18776 18748 18785
rect 6368 18708 6420 18760
rect 8024 18708 8076 18760
rect 13176 18708 13228 18760
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 18052 18708 18104 18760
rect 20076 18776 20128 18828
rect 24676 18776 24728 18828
rect 20904 18751 20956 18760
rect 20904 18717 20913 18751
rect 20913 18717 20947 18751
rect 20947 18717 20956 18751
rect 20904 18708 20956 18717
rect 2228 18640 2280 18692
rect 4896 18640 4948 18692
rect 9036 18640 9088 18692
rect 1860 18572 1912 18624
rect 2688 18572 2740 18624
rect 3424 18572 3476 18624
rect 5264 18615 5316 18624
rect 5264 18581 5273 18615
rect 5273 18581 5307 18615
rect 5307 18581 5316 18615
rect 5264 18572 5316 18581
rect 8116 18572 8168 18624
rect 9588 18572 9640 18624
rect 12072 18572 12124 18624
rect 14740 18572 14792 18624
rect 18604 18572 18656 18624
rect 20352 18572 20404 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2504 18411 2556 18420
rect 2504 18377 2513 18411
rect 2513 18377 2547 18411
rect 2547 18377 2556 18411
rect 2504 18368 2556 18377
rect 7012 18411 7064 18420
rect 7012 18377 7021 18411
rect 7021 18377 7055 18411
rect 7055 18377 7064 18411
rect 7012 18368 7064 18377
rect 9036 18411 9088 18420
rect 9036 18377 9045 18411
rect 9045 18377 9079 18411
rect 9079 18377 9088 18411
rect 9036 18368 9088 18377
rect 11520 18368 11572 18420
rect 11796 18411 11848 18420
rect 11796 18377 11805 18411
rect 11805 18377 11839 18411
rect 11839 18377 11848 18411
rect 11796 18368 11848 18377
rect 15844 18411 15896 18420
rect 15844 18377 15853 18411
rect 15853 18377 15887 18411
rect 15887 18377 15896 18411
rect 15844 18368 15896 18377
rect 20076 18411 20128 18420
rect 20076 18377 20085 18411
rect 20085 18377 20119 18411
rect 20119 18377 20128 18411
rect 20076 18368 20128 18377
rect 3148 18164 3200 18216
rect 7104 18300 7156 18352
rect 7748 18300 7800 18352
rect 12256 18300 12308 18352
rect 16580 18343 16632 18352
rect 5264 18232 5316 18284
rect 4160 18207 4212 18216
rect 4160 18173 4169 18207
rect 4169 18173 4203 18207
rect 4203 18173 4212 18207
rect 4160 18164 4212 18173
rect 4712 18164 4764 18216
rect 5356 18207 5408 18216
rect 5356 18173 5365 18207
rect 5365 18173 5399 18207
rect 5399 18173 5408 18207
rect 5356 18164 5408 18173
rect 6920 18232 6972 18284
rect 8208 18232 8260 18284
rect 6276 18164 6328 18216
rect 8668 18207 8720 18216
rect 8668 18173 8677 18207
rect 8677 18173 8711 18207
rect 8711 18173 8720 18207
rect 8668 18164 8720 18173
rect 9036 18164 9088 18216
rect 9220 18207 9272 18216
rect 9220 18173 9229 18207
rect 9229 18173 9263 18207
rect 9263 18173 9272 18207
rect 9220 18164 9272 18173
rect 9772 18207 9824 18216
rect 9772 18173 9781 18207
rect 9781 18173 9815 18207
rect 9815 18173 9824 18207
rect 9772 18164 9824 18173
rect 11428 18232 11480 18284
rect 12348 18232 12400 18284
rect 16580 18309 16589 18343
rect 16589 18309 16623 18343
rect 16623 18309 16632 18343
rect 16580 18300 16632 18309
rect 24584 18343 24636 18352
rect 24584 18309 24593 18343
rect 24593 18309 24627 18343
rect 24627 18309 24636 18343
rect 24584 18300 24636 18309
rect 14740 18275 14792 18284
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 16028 18275 16080 18284
rect 16028 18241 16037 18275
rect 16037 18241 16071 18275
rect 16071 18241 16080 18275
rect 16028 18232 16080 18241
rect 19248 18232 19300 18284
rect 21916 18232 21968 18284
rect 6644 18096 6696 18148
rect 1768 18028 1820 18080
rect 2596 18071 2648 18080
rect 2596 18037 2605 18071
rect 2605 18037 2639 18071
rect 2639 18037 2648 18071
rect 2596 18028 2648 18037
rect 3148 18071 3200 18080
rect 3148 18037 3157 18071
rect 3157 18037 3191 18071
rect 3191 18037 3200 18071
rect 3148 18028 3200 18037
rect 4068 18028 4120 18080
rect 6368 18028 6420 18080
rect 7472 18139 7524 18148
rect 7472 18105 7481 18139
rect 7481 18105 7515 18139
rect 7515 18105 7524 18139
rect 7472 18096 7524 18105
rect 10876 18096 10928 18148
rect 8116 18028 8168 18080
rect 10048 18028 10100 18080
rect 12624 18096 12676 18148
rect 13176 18139 13228 18148
rect 13176 18105 13185 18139
rect 13185 18105 13219 18139
rect 13219 18105 13228 18139
rect 13176 18096 13228 18105
rect 14188 18164 14240 18216
rect 18420 18164 18472 18216
rect 19651 18207 19703 18216
rect 19651 18173 19660 18207
rect 19660 18173 19694 18207
rect 19694 18173 19703 18207
rect 19651 18164 19703 18173
rect 15844 18096 15896 18148
rect 11704 18028 11756 18080
rect 12256 18071 12308 18080
rect 12256 18037 12265 18071
rect 12265 18037 12299 18071
rect 12299 18037 12308 18071
rect 12256 18028 12308 18037
rect 13452 18071 13504 18080
rect 13452 18037 13461 18071
rect 13461 18037 13495 18071
rect 13495 18037 13504 18071
rect 13452 18028 13504 18037
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 14740 18028 14792 18080
rect 15568 18028 15620 18080
rect 17040 18071 17092 18080
rect 17040 18037 17049 18071
rect 17049 18037 17083 18071
rect 17083 18037 17092 18071
rect 17040 18028 17092 18037
rect 17776 18028 17828 18080
rect 18696 18028 18748 18080
rect 19248 18028 19300 18080
rect 20260 18028 20312 18080
rect 20628 18071 20680 18080
rect 20628 18037 20637 18071
rect 20637 18037 20671 18071
rect 20671 18037 20680 18071
rect 20628 18028 20680 18037
rect 21180 18028 21232 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 4068 17824 4120 17876
rect 5540 17867 5592 17876
rect 5540 17833 5549 17867
rect 5549 17833 5583 17867
rect 5583 17833 5592 17867
rect 5540 17824 5592 17833
rect 7472 17824 7524 17876
rect 9772 17824 9824 17876
rect 10140 17867 10192 17876
rect 10140 17833 10149 17867
rect 10149 17833 10183 17867
rect 10183 17833 10192 17867
rect 10140 17824 10192 17833
rect 13176 17824 13228 17876
rect 16120 17824 16172 17876
rect 6184 17756 6236 17808
rect 7932 17799 7984 17808
rect 7932 17765 7941 17799
rect 7941 17765 7975 17799
rect 7975 17765 7984 17799
rect 7932 17756 7984 17765
rect 8300 17756 8352 17808
rect 10784 17756 10836 17808
rect 2136 17688 2188 17740
rect 4712 17731 4764 17740
rect 4712 17697 4721 17731
rect 4721 17697 4755 17731
rect 4755 17697 4764 17731
rect 4712 17688 4764 17697
rect 5264 17688 5316 17740
rect 11428 17688 11480 17740
rect 12624 17688 12676 17740
rect 12900 17688 12952 17740
rect 13544 17731 13596 17740
rect 13544 17697 13553 17731
rect 13553 17697 13587 17731
rect 13587 17697 13596 17731
rect 13544 17688 13596 17697
rect 14188 17756 14240 17808
rect 15292 17756 15344 17808
rect 16948 17799 17000 17808
rect 16948 17765 16951 17799
rect 16951 17765 16985 17799
rect 16985 17765 17000 17799
rect 16948 17756 17000 17765
rect 17776 17756 17828 17808
rect 15752 17688 15804 17740
rect 16672 17688 16724 17740
rect 17132 17688 17184 17740
rect 18696 17688 18748 17740
rect 20812 17688 20864 17740
rect 22836 17688 22888 17740
rect 23388 17688 23440 17740
rect 3240 17620 3292 17672
rect 6828 17620 6880 17672
rect 8668 17620 8720 17672
rect 10968 17620 11020 17672
rect 12532 17663 12584 17672
rect 12532 17629 12541 17663
rect 12541 17629 12575 17663
rect 12575 17629 12584 17663
rect 12532 17620 12584 17629
rect 11060 17595 11112 17604
rect 11060 17561 11069 17595
rect 11069 17561 11103 17595
rect 11103 17561 11112 17595
rect 11060 17552 11112 17561
rect 11704 17552 11756 17604
rect 1492 17484 1544 17536
rect 4804 17484 4856 17536
rect 14556 17527 14608 17536
rect 14556 17493 14565 17527
rect 14565 17493 14599 17527
rect 14599 17493 14608 17527
rect 14556 17484 14608 17493
rect 16488 17484 16540 17536
rect 17500 17527 17552 17536
rect 17500 17493 17509 17527
rect 17509 17493 17543 17527
rect 17543 17493 17552 17527
rect 17500 17484 17552 17493
rect 18236 17484 18288 17536
rect 21364 17484 21416 17536
rect 22376 17484 22428 17536
rect 22468 17484 22520 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 4712 17280 4764 17332
rect 5080 17280 5132 17332
rect 5264 17280 5316 17332
rect 5540 17280 5592 17332
rect 6368 17280 6420 17332
rect 7932 17280 7984 17332
rect 8024 17323 8076 17332
rect 8024 17289 8033 17323
rect 8033 17289 8067 17323
rect 8067 17289 8076 17323
rect 8024 17280 8076 17289
rect 20812 17280 20864 17332
rect 24768 17323 24820 17332
rect 24768 17289 24777 17323
rect 24777 17289 24811 17323
rect 24811 17289 24820 17323
rect 24768 17280 24820 17289
rect 1584 17144 1636 17196
rect 2044 17144 2096 17196
rect 3792 17144 3844 17196
rect 4712 17187 4764 17196
rect 4712 17153 4721 17187
rect 4721 17153 4755 17187
rect 4755 17153 4764 17187
rect 4712 17144 4764 17153
rect 6644 17144 6696 17196
rect 10140 17212 10192 17264
rect 12624 17212 12676 17264
rect 11060 17144 11112 17196
rect 2044 16983 2096 16992
rect 2044 16949 2053 16983
rect 2053 16949 2087 16983
rect 2087 16949 2096 16983
rect 2044 16940 2096 16949
rect 2136 16940 2188 16992
rect 2596 16940 2648 16992
rect 2780 16983 2832 16992
rect 2780 16949 2789 16983
rect 2789 16949 2823 16983
rect 2823 16949 2832 16983
rect 2780 16940 2832 16949
rect 3976 16940 4028 16992
rect 9772 17076 9824 17128
rect 13820 17212 13872 17264
rect 18236 17212 18288 17264
rect 14556 17144 14608 17196
rect 16120 17187 16172 17196
rect 16120 17153 16129 17187
rect 16129 17153 16163 17187
rect 16163 17153 16172 17187
rect 16120 17144 16172 17153
rect 18420 17187 18472 17196
rect 18420 17153 18429 17187
rect 18429 17153 18463 17187
rect 18463 17153 18472 17187
rect 18420 17144 18472 17153
rect 4804 17051 4856 17060
rect 4804 17017 4813 17051
rect 4813 17017 4847 17051
rect 4847 17017 4856 17051
rect 5356 17051 5408 17060
rect 4804 17008 4856 17017
rect 5356 17017 5365 17051
rect 5365 17017 5399 17051
rect 5399 17017 5408 17051
rect 5356 17008 5408 17017
rect 4988 16940 5040 16992
rect 6184 16940 6236 16992
rect 6368 16940 6420 16992
rect 8944 17008 8996 17060
rect 10784 17008 10836 17060
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 9496 16940 9548 16949
rect 9772 16940 9824 16992
rect 9956 16983 10008 16992
rect 9956 16949 9965 16983
rect 9965 16949 9999 16983
rect 9999 16949 10008 16983
rect 9956 16940 10008 16949
rect 11428 16940 11480 16992
rect 12532 16940 12584 16992
rect 13268 17119 13320 17128
rect 13268 17085 13277 17119
rect 13277 17085 13311 17119
rect 13311 17085 13320 17119
rect 13268 17076 13320 17085
rect 17776 17119 17828 17128
rect 17776 17085 17785 17119
rect 17785 17085 17819 17119
rect 17819 17085 17828 17119
rect 17776 17076 17828 17085
rect 18880 17076 18932 17128
rect 20720 17119 20772 17128
rect 13452 17008 13504 17060
rect 14740 17008 14792 17060
rect 16948 17008 17000 17060
rect 18144 17051 18196 17060
rect 18144 17017 18153 17051
rect 18153 17017 18187 17051
rect 18187 17017 18196 17051
rect 18144 17008 18196 17017
rect 18236 17051 18288 17060
rect 18236 17017 18245 17051
rect 18245 17017 18279 17051
rect 18279 17017 18288 17051
rect 20720 17085 20738 17119
rect 20738 17085 20772 17119
rect 20720 17076 20772 17085
rect 22192 17076 22244 17128
rect 24124 17076 24176 17128
rect 18236 17008 18288 17017
rect 25044 17008 25096 17060
rect 12900 16940 12952 16992
rect 15292 16983 15344 16992
rect 15292 16949 15301 16983
rect 15301 16949 15335 16983
rect 15335 16949 15344 16983
rect 15292 16940 15344 16949
rect 15752 16940 15804 16992
rect 18696 16940 18748 16992
rect 19524 16940 19576 16992
rect 20720 16940 20772 16992
rect 21548 16940 21600 16992
rect 22836 16940 22888 16992
rect 23388 16940 23440 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 4068 16736 4120 16788
rect 6828 16779 6880 16788
rect 6828 16745 6837 16779
rect 6837 16745 6871 16779
rect 6871 16745 6880 16779
rect 6828 16736 6880 16745
rect 7932 16736 7984 16788
rect 8668 16779 8720 16788
rect 8668 16745 8677 16779
rect 8677 16745 8711 16779
rect 8711 16745 8720 16779
rect 8668 16736 8720 16745
rect 11060 16779 11112 16788
rect 11060 16745 11069 16779
rect 11069 16745 11103 16779
rect 11103 16745 11112 16779
rect 11060 16736 11112 16745
rect 12440 16736 12492 16788
rect 14188 16736 14240 16788
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 18144 16736 18196 16788
rect 21272 16736 21324 16788
rect 4252 16668 4304 16720
rect 4712 16668 4764 16720
rect 6000 16711 6052 16720
rect 6000 16677 6009 16711
rect 6009 16677 6043 16711
rect 6043 16677 6052 16711
rect 6000 16668 6052 16677
rect 7840 16711 7892 16720
rect 7840 16677 7849 16711
rect 7849 16677 7883 16711
rect 7883 16677 7892 16711
rect 7840 16668 7892 16677
rect 9588 16668 9640 16720
rect 9864 16711 9916 16720
rect 9864 16677 9873 16711
rect 9873 16677 9907 16711
rect 9907 16677 9916 16711
rect 9864 16668 9916 16677
rect 2136 16600 2188 16652
rect 2780 16600 2832 16652
rect 3700 16600 3752 16652
rect 5356 16600 5408 16652
rect 10968 16668 11020 16720
rect 11336 16668 11388 16720
rect 12348 16668 12400 16720
rect 13268 16668 13320 16720
rect 13452 16668 13504 16720
rect 15292 16668 15344 16720
rect 15844 16668 15896 16720
rect 17500 16668 17552 16720
rect 4344 16532 4396 16584
rect 5908 16575 5960 16584
rect 3332 16464 3384 16516
rect 4068 16464 4120 16516
rect 5908 16541 5917 16575
rect 5917 16541 5951 16575
rect 5951 16541 5960 16575
rect 5908 16532 5960 16541
rect 6184 16532 6236 16584
rect 6828 16532 6880 16584
rect 7748 16575 7800 16584
rect 7748 16541 7757 16575
rect 7757 16541 7791 16575
rect 7791 16541 7800 16575
rect 7748 16532 7800 16541
rect 8024 16575 8076 16584
rect 8024 16541 8033 16575
rect 8033 16541 8067 16575
rect 8067 16541 8076 16575
rect 8024 16532 8076 16541
rect 8668 16532 8720 16584
rect 10140 16532 10192 16584
rect 11520 16532 11572 16584
rect 11704 16575 11756 16584
rect 11704 16541 11713 16575
rect 11713 16541 11747 16575
rect 11747 16541 11756 16575
rect 11704 16532 11756 16541
rect 13176 16575 13228 16584
rect 13176 16541 13185 16575
rect 13185 16541 13219 16575
rect 13219 16541 13228 16575
rect 13176 16532 13228 16541
rect 18972 16600 19024 16652
rect 15476 16532 15528 16584
rect 17684 16575 17736 16584
rect 17684 16541 17693 16575
rect 17693 16541 17727 16575
rect 17727 16541 17736 16575
rect 17684 16532 17736 16541
rect 14740 16464 14792 16516
rect 18420 16532 18472 16584
rect 19892 16711 19944 16720
rect 19892 16677 19901 16711
rect 19901 16677 19935 16711
rect 19935 16677 19944 16711
rect 19892 16668 19944 16677
rect 24676 16668 24728 16720
rect 21088 16600 21140 16652
rect 19064 16532 19116 16584
rect 22928 16643 22980 16652
rect 22928 16609 22972 16643
rect 22972 16609 22980 16643
rect 22928 16600 22980 16609
rect 23112 16600 23164 16652
rect 22284 16532 22336 16584
rect 22652 16532 22704 16584
rect 25504 16600 25556 16652
rect 20720 16464 20772 16516
rect 1768 16396 1820 16448
rect 1952 16396 2004 16448
rect 2044 16396 2096 16448
rect 3148 16396 3200 16448
rect 8392 16396 8444 16448
rect 25412 16396 25464 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1400 16192 1452 16244
rect 4804 16192 4856 16244
rect 6000 16192 6052 16244
rect 6184 16235 6236 16244
rect 6184 16201 6193 16235
rect 6193 16201 6227 16235
rect 6227 16201 6236 16235
rect 6184 16192 6236 16201
rect 6644 16235 6696 16244
rect 6644 16201 6653 16235
rect 6653 16201 6687 16235
rect 6687 16201 6696 16235
rect 6644 16192 6696 16201
rect 7840 16192 7892 16244
rect 9496 16192 9548 16244
rect 10784 16235 10836 16244
rect 10784 16201 10793 16235
rect 10793 16201 10827 16235
rect 10827 16201 10836 16235
rect 10784 16192 10836 16201
rect 11336 16235 11388 16244
rect 11336 16201 11345 16235
rect 11345 16201 11379 16235
rect 11379 16201 11388 16235
rect 11336 16192 11388 16201
rect 15844 16235 15896 16244
rect 15844 16201 15853 16235
rect 15853 16201 15887 16235
rect 15887 16201 15896 16235
rect 15844 16192 15896 16201
rect 17500 16235 17552 16244
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 24768 16235 24820 16244
rect 24768 16201 24777 16235
rect 24777 16201 24811 16235
rect 24811 16201 24820 16235
rect 24768 16192 24820 16201
rect 2320 16124 2372 16176
rect 9128 16124 9180 16176
rect 15476 16167 15528 16176
rect 15476 16133 15485 16167
rect 15485 16133 15519 16167
rect 15519 16133 15528 16167
rect 15476 16124 15528 16133
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 2872 16031 2924 16040
rect 2872 15997 2881 16031
rect 2881 15997 2915 16031
rect 2915 15997 2924 16031
rect 2872 15988 2924 15997
rect 3608 15988 3660 16040
rect 3332 15963 3384 15972
rect 3332 15929 3341 15963
rect 3341 15929 3375 15963
rect 3375 15929 3384 15963
rect 3332 15920 3384 15929
rect 3700 15963 3752 15972
rect 3700 15929 3709 15963
rect 3709 15929 3743 15963
rect 3743 15929 3752 15963
rect 3700 15920 3752 15929
rect 7472 16056 7524 16108
rect 8116 16056 8168 16108
rect 8668 16056 8720 16108
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 15200 16056 15252 16108
rect 16488 16099 16540 16108
rect 16488 16065 16497 16099
rect 16497 16065 16531 16099
rect 16531 16065 16540 16099
rect 16488 16056 16540 16065
rect 19432 16124 19484 16176
rect 18604 16056 18656 16108
rect 19524 16056 19576 16108
rect 19892 16056 19944 16108
rect 21088 16099 21140 16108
rect 21088 16065 21097 16099
rect 21097 16065 21131 16099
rect 21131 16065 21140 16099
rect 21088 16056 21140 16065
rect 21732 16056 21784 16108
rect 4252 15920 4304 15972
rect 6368 15920 6420 15972
rect 7840 15963 7892 15972
rect 7840 15929 7849 15963
rect 7849 15929 7883 15963
rect 7883 15929 7892 15963
rect 7840 15920 7892 15929
rect 13084 16031 13136 16040
rect 13084 15997 13093 16031
rect 13093 15997 13127 16031
rect 13127 15997 13136 16031
rect 13084 15988 13136 15997
rect 16304 15988 16356 16040
rect 13452 15920 13504 15972
rect 16580 15963 16632 15972
rect 5356 15895 5408 15904
rect 5356 15861 5365 15895
rect 5365 15861 5399 15895
rect 5399 15861 5408 15895
rect 5356 15852 5408 15861
rect 9312 15895 9364 15904
rect 9312 15861 9321 15895
rect 9321 15861 9355 15895
rect 9355 15861 9364 15895
rect 9312 15852 9364 15861
rect 9864 15852 9916 15904
rect 11520 15852 11572 15904
rect 13268 15852 13320 15904
rect 14740 15852 14792 15904
rect 16580 15929 16589 15963
rect 16589 15929 16623 15963
rect 16623 15929 16632 15963
rect 16580 15920 16632 15929
rect 18788 15963 18840 15972
rect 18788 15929 18797 15963
rect 18797 15929 18831 15963
rect 18831 15929 18840 15963
rect 18788 15920 18840 15929
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 19064 15852 19116 15861
rect 19248 15852 19300 15904
rect 20720 15920 20772 15972
rect 22100 15963 22152 15972
rect 22100 15929 22109 15963
rect 22109 15929 22143 15963
rect 22143 15929 22152 15963
rect 22928 15988 22980 16040
rect 22100 15920 22152 15929
rect 22560 15920 22612 15972
rect 21824 15852 21876 15904
rect 22192 15852 22244 15904
rect 25504 15895 25556 15904
rect 25504 15861 25513 15895
rect 25513 15861 25547 15895
rect 25547 15861 25556 15895
rect 25504 15852 25556 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1676 15648 1728 15700
rect 4252 15691 4304 15700
rect 4252 15657 4261 15691
rect 4261 15657 4295 15691
rect 4295 15657 4304 15691
rect 4252 15648 4304 15657
rect 5264 15691 5316 15700
rect 5264 15657 5273 15691
rect 5273 15657 5307 15691
rect 5307 15657 5316 15691
rect 5264 15648 5316 15657
rect 7840 15648 7892 15700
rect 8116 15691 8168 15700
rect 8116 15657 8125 15691
rect 8125 15657 8159 15691
rect 8159 15657 8168 15691
rect 8116 15648 8168 15657
rect 9588 15648 9640 15700
rect 4896 15580 4948 15632
rect 2412 15512 2464 15564
rect 2964 15555 3016 15564
rect 2964 15521 2973 15555
rect 2973 15521 3007 15555
rect 3007 15521 3016 15555
rect 2964 15512 3016 15521
rect 5172 15555 5224 15564
rect 5172 15521 5181 15555
rect 5181 15521 5215 15555
rect 5215 15521 5224 15555
rect 5172 15512 5224 15521
rect 5264 15512 5316 15564
rect 6368 15580 6420 15632
rect 6828 15580 6880 15632
rect 6552 15555 6604 15564
rect 6552 15521 6561 15555
rect 6561 15521 6595 15555
rect 6595 15521 6604 15555
rect 6552 15512 6604 15521
rect 7012 15512 7064 15564
rect 8484 15512 8536 15564
rect 9588 15512 9640 15564
rect 9772 15512 9824 15564
rect 9956 15512 10008 15564
rect 11336 15512 11388 15564
rect 12256 15648 12308 15700
rect 13176 15648 13228 15700
rect 14832 15691 14884 15700
rect 14832 15657 14841 15691
rect 14841 15657 14875 15691
rect 14875 15657 14884 15691
rect 14832 15648 14884 15657
rect 16488 15691 16540 15700
rect 16488 15657 16497 15691
rect 16497 15657 16531 15691
rect 16531 15657 16540 15691
rect 16488 15648 16540 15657
rect 18236 15691 18288 15700
rect 18236 15657 18245 15691
rect 18245 15657 18279 15691
rect 18279 15657 18288 15691
rect 18236 15648 18288 15657
rect 18604 15691 18656 15700
rect 18604 15657 18613 15691
rect 18613 15657 18647 15691
rect 18647 15657 18656 15691
rect 18604 15648 18656 15657
rect 19524 15648 19576 15700
rect 13084 15580 13136 15632
rect 13268 15580 13320 15632
rect 14740 15580 14792 15632
rect 16764 15580 16816 15632
rect 17684 15580 17736 15632
rect 18788 15580 18840 15632
rect 18880 15623 18932 15632
rect 18880 15589 18889 15623
rect 18889 15589 18923 15623
rect 18923 15589 18932 15623
rect 19432 15623 19484 15632
rect 18880 15580 18932 15589
rect 19432 15589 19441 15623
rect 19441 15589 19475 15623
rect 19475 15589 19484 15623
rect 19432 15580 19484 15589
rect 21180 15623 21232 15632
rect 21180 15589 21189 15623
rect 21189 15589 21223 15623
rect 21223 15589 21232 15623
rect 21180 15580 21232 15589
rect 21456 15580 21508 15632
rect 11980 15555 12032 15564
rect 11980 15521 11989 15555
rect 11989 15521 12023 15555
rect 12023 15521 12032 15555
rect 11980 15512 12032 15521
rect 12348 15512 12400 15564
rect 22928 15512 22980 15564
rect 23756 15555 23808 15564
rect 23756 15521 23774 15555
rect 23774 15521 23808 15555
rect 23756 15512 23808 15521
rect 23940 15512 23992 15564
rect 24216 15512 24268 15564
rect 25136 15512 25188 15564
rect 1676 15376 1728 15428
rect 3608 15444 3660 15496
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 12256 15444 12308 15496
rect 15476 15444 15528 15496
rect 17224 15487 17276 15496
rect 17224 15453 17233 15487
rect 17233 15453 17267 15487
rect 17267 15453 17276 15487
rect 17224 15444 17276 15453
rect 18604 15444 18656 15496
rect 22100 15487 22152 15496
rect 22100 15453 22109 15487
rect 22109 15453 22143 15487
rect 22143 15453 22152 15487
rect 22100 15444 22152 15453
rect 22284 15444 22336 15496
rect 2872 15376 2924 15428
rect 3700 15376 3752 15428
rect 15292 15376 15344 15428
rect 21732 15419 21784 15428
rect 21732 15385 21741 15419
rect 21741 15385 21775 15419
rect 21775 15385 21784 15419
rect 21732 15376 21784 15385
rect 1308 15308 1360 15360
rect 2136 15308 2188 15360
rect 3608 15351 3660 15360
rect 3608 15317 3617 15351
rect 3617 15317 3651 15351
rect 3651 15317 3660 15351
rect 3608 15308 3660 15317
rect 4344 15308 4396 15360
rect 6368 15351 6420 15360
rect 6368 15317 6377 15351
rect 6377 15317 6411 15351
rect 6411 15317 6420 15351
rect 6368 15308 6420 15317
rect 7748 15308 7800 15360
rect 8208 15308 8260 15360
rect 12348 15308 12400 15360
rect 14740 15308 14792 15360
rect 22468 15308 22520 15360
rect 23480 15308 23532 15360
rect 25228 15308 25280 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1952 15147 2004 15156
rect 1952 15113 1961 15147
rect 1961 15113 1995 15147
rect 1995 15113 2004 15147
rect 1952 15104 2004 15113
rect 2412 15147 2464 15156
rect 2412 15113 2421 15147
rect 2421 15113 2455 15147
rect 2455 15113 2464 15147
rect 2412 15104 2464 15113
rect 4620 15147 4672 15156
rect 4620 15113 4629 15147
rect 4629 15113 4663 15147
rect 4663 15113 4672 15147
rect 4620 15104 4672 15113
rect 2320 14900 2372 14952
rect 3148 14943 3200 14952
rect 3148 14909 3157 14943
rect 3157 14909 3191 14943
rect 3191 14909 3200 14943
rect 3148 14900 3200 14909
rect 3700 14900 3752 14952
rect 5080 15036 5132 15088
rect 4344 15011 4396 15020
rect 4344 14977 4353 15011
rect 4353 14977 4387 15011
rect 4387 14977 4396 15011
rect 4344 14968 4396 14977
rect 4160 14943 4212 14952
rect 4160 14909 4169 14943
rect 4169 14909 4203 14943
rect 4203 14909 4212 14943
rect 4160 14900 4212 14909
rect 5080 14900 5132 14952
rect 7012 15104 7064 15156
rect 9772 15104 9824 15156
rect 9956 15036 10008 15088
rect 6368 14968 6420 15020
rect 8668 14968 8720 15020
rect 7012 14900 7064 14952
rect 11428 15104 11480 15156
rect 11980 15104 12032 15156
rect 12440 15104 12492 15156
rect 12716 15104 12768 15156
rect 14740 15147 14792 15156
rect 14740 15113 14749 15147
rect 14749 15113 14783 15147
rect 14783 15113 14792 15147
rect 14740 15104 14792 15113
rect 16764 15147 16816 15156
rect 16764 15113 16773 15147
rect 16773 15113 16807 15147
rect 16807 15113 16816 15147
rect 16764 15104 16816 15113
rect 18880 15104 18932 15156
rect 21180 15104 21232 15156
rect 22928 15104 22980 15156
rect 15936 15079 15988 15088
rect 15936 15045 15945 15079
rect 15945 15045 15979 15079
rect 15979 15045 15988 15079
rect 15936 15036 15988 15045
rect 16580 15036 16632 15088
rect 12348 14968 12400 15020
rect 13912 14968 13964 15020
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 16396 15011 16448 15020
rect 16396 14977 16405 15011
rect 16405 14977 16439 15011
rect 16439 14977 16448 15011
rect 16396 14968 16448 14977
rect 17132 14968 17184 15020
rect 18236 14968 18288 15020
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 11336 14943 11388 14952
rect 11336 14909 11345 14943
rect 11345 14909 11379 14943
rect 11379 14909 11388 14943
rect 11336 14900 11388 14909
rect 11980 14900 12032 14952
rect 12716 14900 12768 14952
rect 16304 14900 16356 14952
rect 20536 14943 20588 14952
rect 20536 14909 20545 14943
rect 20545 14909 20579 14943
rect 20579 14909 20588 14943
rect 20536 14900 20588 14909
rect 21456 14943 21508 14952
rect 21456 14909 21465 14943
rect 21465 14909 21499 14943
rect 21499 14909 21508 14943
rect 21456 14900 21508 14909
rect 21640 14900 21692 14952
rect 24032 14900 24084 14952
rect 2136 14764 2188 14816
rect 2964 14832 3016 14884
rect 4344 14764 4396 14816
rect 6828 14832 6880 14884
rect 8668 14875 8720 14884
rect 8668 14841 8677 14875
rect 8677 14841 8711 14875
rect 8711 14841 8720 14875
rect 8668 14832 8720 14841
rect 8760 14875 8812 14884
rect 8760 14841 8769 14875
rect 8769 14841 8803 14875
rect 8803 14841 8812 14875
rect 8760 14832 8812 14841
rect 11428 14832 11480 14884
rect 13912 14875 13964 14884
rect 13912 14841 13921 14875
rect 13921 14841 13955 14875
rect 13955 14841 13964 14875
rect 13912 14832 13964 14841
rect 15384 14832 15436 14884
rect 17960 14832 18012 14884
rect 5172 14764 5224 14816
rect 6552 14807 6604 14816
rect 6552 14773 6561 14807
rect 6561 14773 6595 14807
rect 6595 14773 6604 14807
rect 6552 14764 6604 14773
rect 7748 14807 7800 14816
rect 7748 14773 7757 14807
rect 7757 14773 7791 14807
rect 7791 14773 7800 14807
rect 7748 14764 7800 14773
rect 8484 14807 8536 14816
rect 8484 14773 8493 14807
rect 8493 14773 8527 14807
rect 8527 14773 8536 14807
rect 8484 14764 8536 14773
rect 12716 14764 12768 14816
rect 12900 14764 12952 14816
rect 13084 14764 13136 14816
rect 13268 14807 13320 14816
rect 13268 14773 13277 14807
rect 13277 14773 13311 14807
rect 13311 14773 13320 14807
rect 13268 14764 13320 14773
rect 19248 14832 19300 14884
rect 19340 14764 19392 14816
rect 19524 14764 19576 14816
rect 23572 14832 23624 14884
rect 20996 14764 21048 14816
rect 23480 14764 23532 14816
rect 23940 14764 23992 14816
rect 25136 14807 25188 14816
rect 25136 14773 25145 14807
rect 25145 14773 25179 14807
rect 25179 14773 25188 14807
rect 25136 14764 25188 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 3148 14560 3200 14612
rect 3332 14560 3384 14612
rect 5080 14560 5132 14612
rect 5264 14560 5316 14612
rect 8668 14560 8720 14612
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 11336 14560 11388 14612
rect 13820 14603 13872 14612
rect 13820 14569 13829 14603
rect 13829 14569 13863 14603
rect 13863 14569 13872 14603
rect 13820 14560 13872 14569
rect 17224 14603 17276 14612
rect 17224 14569 17233 14603
rect 17233 14569 17267 14603
rect 17267 14569 17276 14603
rect 17224 14560 17276 14569
rect 3700 14535 3752 14544
rect 3700 14501 3709 14535
rect 3709 14501 3743 14535
rect 3743 14501 3752 14535
rect 3700 14492 3752 14501
rect 4068 14492 4120 14544
rect 7748 14535 7800 14544
rect 1584 14424 1636 14476
rect 3148 14424 3200 14476
rect 3608 14424 3660 14476
rect 4160 14467 4212 14476
rect 4160 14433 4169 14467
rect 4169 14433 4203 14467
rect 4203 14433 4212 14467
rect 4160 14424 4212 14433
rect 7748 14501 7757 14535
rect 7757 14501 7791 14535
rect 7791 14501 7800 14535
rect 7748 14492 7800 14501
rect 8116 14492 8168 14544
rect 8760 14492 8812 14544
rect 6276 14467 6328 14476
rect 6276 14433 6285 14467
rect 6285 14433 6319 14467
rect 6319 14433 6328 14467
rect 6276 14424 6328 14433
rect 9772 14467 9824 14476
rect 9772 14433 9781 14467
rect 9781 14433 9815 14467
rect 9815 14433 9824 14467
rect 9772 14424 9824 14433
rect 6184 14356 6236 14408
rect 6368 14399 6420 14408
rect 6368 14365 6377 14399
rect 6377 14365 6411 14399
rect 6411 14365 6420 14399
rect 6368 14356 6420 14365
rect 7932 14356 7984 14408
rect 8024 14399 8076 14408
rect 8024 14365 8033 14399
rect 8033 14365 8067 14399
rect 8067 14365 8076 14399
rect 8024 14356 8076 14365
rect 9588 14356 9640 14408
rect 11060 14424 11112 14476
rect 12256 14492 12308 14544
rect 12992 14535 13044 14544
rect 12992 14501 13001 14535
rect 13001 14501 13035 14535
rect 13035 14501 13044 14535
rect 12992 14492 13044 14501
rect 14096 14492 14148 14544
rect 11704 14467 11756 14476
rect 11704 14433 11713 14467
rect 11713 14433 11747 14467
rect 11747 14433 11756 14467
rect 11704 14424 11756 14433
rect 11796 14356 11848 14408
rect 12072 14356 12124 14408
rect 12900 14399 12952 14408
rect 12900 14365 12909 14399
rect 12909 14365 12943 14399
rect 12943 14365 12952 14399
rect 12900 14356 12952 14365
rect 13820 14356 13872 14408
rect 17408 14492 17460 14544
rect 17868 14560 17920 14612
rect 20536 14560 20588 14612
rect 24768 14603 24820 14612
rect 24768 14569 24777 14603
rect 24777 14569 24811 14603
rect 24811 14569 24820 14603
rect 24768 14560 24820 14569
rect 18052 14492 18104 14544
rect 18972 14492 19024 14544
rect 19524 14492 19576 14544
rect 20168 14492 20220 14544
rect 21088 14535 21140 14544
rect 21088 14501 21097 14535
rect 21097 14501 21131 14535
rect 21131 14501 21140 14535
rect 21088 14492 21140 14501
rect 22744 14467 22796 14476
rect 22744 14433 22753 14467
rect 22753 14433 22787 14467
rect 22787 14433 22796 14467
rect 22744 14424 22796 14433
rect 22928 14467 22980 14476
rect 22928 14433 22937 14467
rect 22937 14433 22971 14467
rect 22971 14433 22980 14467
rect 22928 14424 22980 14433
rect 24676 14424 24728 14476
rect 14832 14356 14884 14408
rect 15476 14356 15528 14408
rect 16028 14399 16080 14408
rect 16028 14365 16037 14399
rect 16037 14365 16071 14399
rect 16071 14365 16080 14399
rect 16028 14356 16080 14365
rect 18788 14356 18840 14408
rect 19248 14356 19300 14408
rect 20996 14399 21048 14408
rect 20996 14365 21005 14399
rect 21005 14365 21039 14399
rect 21039 14365 21048 14399
rect 20996 14356 21048 14365
rect 21456 14399 21508 14408
rect 21456 14365 21465 14399
rect 21465 14365 21499 14399
rect 21499 14365 21508 14399
rect 21456 14356 21508 14365
rect 3056 14288 3108 14340
rect 3700 14288 3752 14340
rect 13544 14288 13596 14340
rect 15292 14288 15344 14340
rect 7288 14220 7340 14272
rect 10140 14220 10192 14272
rect 21640 14220 21692 14272
rect 22284 14263 22336 14272
rect 22284 14229 22293 14263
rect 22293 14229 22327 14263
rect 22327 14229 22336 14263
rect 22284 14220 22336 14229
rect 23756 14263 23808 14272
rect 23756 14229 23765 14263
rect 23765 14229 23799 14263
rect 23799 14229 23808 14263
rect 23756 14220 23808 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1492 14016 1544 14068
rect 2780 14016 2832 14068
rect 4160 14016 4212 14068
rect 6184 14016 6236 14068
rect 6276 14016 6328 14068
rect 8116 14059 8168 14068
rect 8116 14025 8125 14059
rect 8125 14025 8159 14059
rect 8159 14025 8168 14059
rect 8116 14016 8168 14025
rect 8300 14016 8352 14068
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 11060 14016 11112 14068
rect 11704 14059 11756 14068
rect 11704 14025 11713 14059
rect 11713 14025 11747 14059
rect 11747 14025 11756 14059
rect 11704 14016 11756 14025
rect 12900 14016 12952 14068
rect 18972 14016 19024 14068
rect 21088 14016 21140 14068
rect 24676 14059 24728 14068
rect 24676 14025 24685 14059
rect 24685 14025 24719 14059
rect 24719 14025 24728 14059
rect 24676 14016 24728 14025
rect 24860 14016 24912 14068
rect 2688 13948 2740 14000
rect 3148 13880 3200 13932
rect 5540 13880 5592 13932
rect 6276 13880 6328 13932
rect 7472 13948 7524 14000
rect 8668 13948 8720 14000
rect 3332 13812 3384 13864
rect 4712 13855 4764 13864
rect 4712 13821 4721 13855
rect 4721 13821 4755 13855
rect 4755 13821 4764 13855
rect 4712 13812 4764 13821
rect 5172 13855 5224 13864
rect 5172 13821 5181 13855
rect 5181 13821 5215 13855
rect 5215 13821 5224 13855
rect 5172 13812 5224 13821
rect 8208 13812 8260 13864
rect 8392 13812 8444 13864
rect 9220 13812 9272 13864
rect 12992 13948 13044 14000
rect 13636 13991 13688 14000
rect 13636 13957 13645 13991
rect 13645 13957 13679 13991
rect 13679 13957 13688 13991
rect 13636 13948 13688 13957
rect 13820 13948 13872 14000
rect 18052 13948 18104 14000
rect 18788 13948 18840 14000
rect 12440 13923 12492 13932
rect 12440 13889 12449 13923
rect 12449 13889 12483 13923
rect 12483 13889 12492 13923
rect 12440 13880 12492 13889
rect 15200 13923 15252 13932
rect 15200 13889 15209 13923
rect 15209 13889 15243 13923
rect 15243 13889 15252 13923
rect 15200 13880 15252 13889
rect 15936 13880 15988 13932
rect 18236 13880 18288 13932
rect 20076 13880 20128 13932
rect 20628 13880 20680 13932
rect 22284 13948 22336 14000
rect 23020 13948 23072 14000
rect 21732 13923 21784 13932
rect 21732 13889 21741 13923
rect 21741 13889 21775 13923
rect 21775 13889 21784 13923
rect 21732 13880 21784 13889
rect 3976 13744 4028 13796
rect 5356 13787 5408 13796
rect 5356 13753 5365 13787
rect 5365 13753 5399 13787
rect 5399 13753 5408 13787
rect 5356 13744 5408 13753
rect 7288 13787 7340 13796
rect 7288 13753 7297 13787
rect 7297 13753 7331 13787
rect 7331 13753 7340 13787
rect 7288 13744 7340 13753
rect 9128 13744 9180 13796
rect 10968 13812 11020 13864
rect 10140 13787 10192 13796
rect 10140 13753 10149 13787
rect 10149 13753 10183 13787
rect 10183 13753 10192 13787
rect 10140 13744 10192 13753
rect 5540 13676 5592 13728
rect 9220 13719 9272 13728
rect 9220 13685 9229 13719
rect 9229 13685 9263 13719
rect 9263 13685 9272 13719
rect 9220 13676 9272 13685
rect 9312 13676 9364 13728
rect 11336 13676 11388 13728
rect 12072 13676 12124 13728
rect 16856 13812 16908 13864
rect 17224 13812 17276 13864
rect 22744 13812 22796 13864
rect 23756 13855 23808 13864
rect 23756 13821 23765 13855
rect 23765 13821 23799 13855
rect 23799 13821 23808 13855
rect 23756 13812 23808 13821
rect 17316 13744 17368 13796
rect 18144 13744 18196 13796
rect 18880 13744 18932 13796
rect 20168 13744 20220 13796
rect 21640 13744 21692 13796
rect 22192 13744 22244 13796
rect 22928 13787 22980 13796
rect 22928 13753 22937 13787
rect 22937 13753 22971 13787
rect 22971 13753 22980 13787
rect 22928 13744 22980 13753
rect 23848 13744 23900 13796
rect 24952 13812 25004 13864
rect 23480 13676 23532 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 3332 13515 3384 13524
rect 3332 13481 3341 13515
rect 3341 13481 3375 13515
rect 3375 13481 3384 13515
rect 3332 13472 3384 13481
rect 2688 13404 2740 13456
rect 2780 13404 2832 13456
rect 4068 13472 4120 13524
rect 3976 13404 4028 13456
rect 4896 13404 4948 13456
rect 6368 13472 6420 13524
rect 7288 13472 7340 13524
rect 7472 13515 7524 13524
rect 7472 13481 7481 13515
rect 7481 13481 7515 13515
rect 7515 13481 7524 13515
rect 7472 13472 7524 13481
rect 9128 13515 9180 13524
rect 9128 13481 9137 13515
rect 9137 13481 9171 13515
rect 9171 13481 9180 13515
rect 9128 13472 9180 13481
rect 9588 13472 9640 13524
rect 10140 13472 10192 13524
rect 11060 13472 11112 13524
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 13728 13472 13780 13524
rect 14832 13472 14884 13524
rect 17868 13472 17920 13524
rect 18236 13515 18288 13524
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 20076 13472 20128 13524
rect 20996 13472 21048 13524
rect 6552 13404 6604 13456
rect 8208 13447 8260 13456
rect 8208 13413 8217 13447
rect 8217 13413 8251 13447
rect 8251 13413 8260 13447
rect 8208 13404 8260 13413
rect 9864 13404 9916 13456
rect 12072 13404 12124 13456
rect 12992 13404 13044 13456
rect 15384 13404 15436 13456
rect 16028 13447 16080 13456
rect 16028 13413 16037 13447
rect 16037 13413 16071 13447
rect 16071 13413 16080 13447
rect 16028 13404 16080 13413
rect 17040 13447 17092 13456
rect 17040 13413 17049 13447
rect 17049 13413 17083 13447
rect 17083 13413 17092 13447
rect 17040 13404 17092 13413
rect 18604 13447 18656 13456
rect 18604 13413 18613 13447
rect 18613 13413 18647 13447
rect 18647 13413 18656 13447
rect 18604 13404 18656 13413
rect 19248 13404 19300 13456
rect 20168 13404 20220 13456
rect 21548 13447 21600 13456
rect 21548 13413 21557 13447
rect 21557 13413 21591 13447
rect 21591 13413 21600 13447
rect 21548 13404 21600 13413
rect 23388 13404 23440 13456
rect 11428 13379 11480 13388
rect 11428 13345 11437 13379
rect 11437 13345 11471 13379
rect 11471 13345 11480 13379
rect 11428 13336 11480 13345
rect 12624 13379 12676 13388
rect 12624 13345 12633 13379
rect 12633 13345 12667 13379
rect 12667 13345 12676 13379
rect 12624 13336 12676 13345
rect 24216 13336 24268 13388
rect 2504 13268 2556 13320
rect 4068 13311 4120 13320
rect 4068 13277 4077 13311
rect 4077 13277 4111 13311
rect 4111 13277 4120 13311
rect 4068 13268 4120 13277
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 8300 13268 8352 13320
rect 9772 13268 9824 13320
rect 10784 13268 10836 13320
rect 14556 13268 14608 13320
rect 17224 13268 17276 13320
rect 17316 13311 17368 13320
rect 17316 13277 17325 13311
rect 17325 13277 17359 13311
rect 17359 13277 17368 13311
rect 18512 13311 18564 13320
rect 17316 13268 17368 13277
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 18788 13311 18840 13320
rect 18788 13277 18797 13311
rect 18797 13277 18831 13311
rect 18831 13277 18840 13311
rect 18788 13268 18840 13277
rect 21456 13311 21508 13320
rect 21456 13277 21465 13311
rect 21465 13277 21499 13311
rect 21499 13277 21508 13311
rect 21456 13268 21508 13277
rect 22468 13268 22520 13320
rect 2872 13243 2924 13252
rect 2872 13209 2881 13243
rect 2881 13209 2915 13243
rect 2915 13209 2924 13243
rect 2872 13200 2924 13209
rect 4620 13200 4672 13252
rect 9404 13200 9456 13252
rect 11060 13200 11112 13252
rect 20720 13200 20772 13252
rect 21732 13200 21784 13252
rect 22100 13200 22152 13252
rect 1676 13175 1728 13184
rect 1676 13141 1685 13175
rect 1685 13141 1719 13175
rect 1719 13141 1728 13175
rect 1676 13132 1728 13141
rect 3976 13132 4028 13184
rect 7932 13175 7984 13184
rect 7932 13141 7941 13175
rect 7941 13141 7975 13175
rect 7975 13141 7984 13175
rect 7932 13132 7984 13141
rect 9680 13132 9732 13184
rect 11796 13132 11848 13184
rect 13820 13175 13872 13184
rect 13820 13141 13829 13175
rect 13829 13141 13863 13175
rect 13863 13141 13872 13175
rect 13820 13132 13872 13141
rect 21088 13175 21140 13184
rect 21088 13141 21097 13175
rect 21097 13141 21131 13175
rect 21131 13141 21140 13175
rect 21088 13132 21140 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2504 12928 2556 12980
rect 2688 12971 2740 12980
rect 2688 12937 2697 12971
rect 2697 12937 2731 12971
rect 2731 12937 2740 12971
rect 2688 12928 2740 12937
rect 4068 12928 4120 12980
rect 8116 12928 8168 12980
rect 8484 12928 8536 12980
rect 8760 12971 8812 12980
rect 8760 12937 8769 12971
rect 8769 12937 8803 12971
rect 8803 12937 8812 12971
rect 8760 12928 8812 12937
rect 10784 12971 10836 12980
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 11428 12928 11480 12980
rect 11980 12928 12032 12980
rect 13544 12928 13596 12980
rect 15384 12971 15436 12980
rect 15384 12937 15393 12971
rect 15393 12937 15427 12971
rect 15427 12937 15436 12971
rect 15384 12928 15436 12937
rect 21548 12928 21600 12980
rect 22468 12971 22520 12980
rect 22468 12937 22477 12971
rect 22477 12937 22511 12971
rect 22511 12937 22520 12971
rect 22468 12928 22520 12937
rect 23388 12971 23440 12980
rect 23388 12937 23397 12971
rect 23397 12937 23431 12971
rect 23431 12937 23440 12971
rect 23388 12928 23440 12937
rect 24768 12928 24820 12980
rect 25596 12971 25648 12980
rect 25596 12937 25605 12971
rect 25605 12937 25639 12971
rect 25639 12937 25648 12971
rect 25596 12928 25648 12937
rect 1768 12860 1820 12912
rect 6644 12860 6696 12912
rect 4068 12792 4120 12844
rect 4620 12792 4672 12844
rect 12992 12860 13044 12912
rect 8208 12792 8260 12844
rect 10324 12792 10376 12844
rect 11060 12792 11112 12844
rect 12440 12792 12492 12844
rect 13820 12792 13872 12844
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 6828 12767 6880 12776
rect 3884 12699 3936 12708
rect 3884 12665 3893 12699
rect 3893 12665 3927 12699
rect 3927 12665 3936 12699
rect 3884 12656 3936 12665
rect 3976 12699 4028 12708
rect 3976 12665 3985 12699
rect 3985 12665 4019 12699
rect 4019 12665 4028 12699
rect 3976 12656 4028 12665
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 7288 12724 7340 12776
rect 11244 12724 11296 12776
rect 12072 12724 12124 12776
rect 12716 12724 12768 12776
rect 6000 12656 6052 12708
rect 2780 12588 2832 12640
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 6552 12656 6604 12708
rect 7104 12656 7156 12708
rect 9864 12656 9916 12708
rect 10140 12656 10192 12708
rect 11060 12656 11112 12708
rect 13728 12699 13780 12708
rect 13728 12665 13737 12699
rect 13737 12665 13771 12699
rect 13771 12665 13780 12699
rect 15936 12860 15988 12912
rect 18880 12903 18932 12912
rect 18880 12869 18889 12903
rect 18889 12869 18923 12903
rect 18923 12869 18932 12903
rect 18880 12860 18932 12869
rect 22284 12860 22336 12912
rect 24216 12860 24268 12912
rect 15568 12792 15620 12844
rect 16028 12792 16080 12844
rect 17960 12792 18012 12844
rect 18144 12792 18196 12844
rect 20628 12792 20680 12844
rect 21088 12792 21140 12844
rect 21456 12792 21508 12844
rect 22008 12792 22060 12844
rect 22468 12792 22520 12844
rect 22744 12792 22796 12844
rect 19800 12767 19852 12776
rect 19800 12733 19844 12767
rect 19844 12733 19852 12767
rect 19800 12724 19852 12733
rect 24860 12792 24912 12844
rect 25228 12792 25280 12844
rect 25596 12724 25648 12776
rect 13728 12656 13780 12665
rect 4896 12588 4948 12597
rect 9772 12588 9824 12640
rect 10048 12588 10100 12640
rect 14556 12631 14608 12640
rect 14556 12597 14565 12631
rect 14565 12597 14599 12631
rect 14599 12597 14608 12631
rect 14556 12588 14608 12597
rect 15936 12699 15988 12708
rect 15936 12665 15945 12699
rect 15945 12665 15979 12699
rect 15979 12665 15988 12699
rect 15936 12656 15988 12665
rect 17040 12656 17092 12708
rect 18420 12699 18472 12708
rect 18420 12665 18429 12699
rect 18429 12665 18463 12699
rect 18463 12665 18472 12699
rect 18420 12656 18472 12665
rect 18604 12656 18656 12708
rect 21180 12656 21232 12708
rect 22008 12656 22060 12708
rect 22192 12656 22244 12708
rect 24952 12656 25004 12708
rect 16396 12588 16448 12640
rect 17224 12631 17276 12640
rect 17224 12597 17233 12631
rect 17233 12597 17267 12631
rect 17267 12597 17276 12631
rect 17224 12588 17276 12597
rect 18512 12588 18564 12640
rect 22284 12588 22336 12640
rect 22744 12588 22796 12640
rect 23296 12588 23348 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 3976 12384 4028 12436
rect 4160 12427 4212 12436
rect 4160 12393 4169 12427
rect 4169 12393 4203 12427
rect 4203 12393 4212 12427
rect 4160 12384 4212 12393
rect 4344 12384 4396 12436
rect 9036 12384 9088 12436
rect 9956 12427 10008 12436
rect 9956 12393 9965 12427
rect 9965 12393 9999 12427
rect 9999 12393 10008 12427
rect 9956 12384 10008 12393
rect 10140 12384 10192 12436
rect 12624 12384 12676 12436
rect 13728 12427 13780 12436
rect 13728 12393 13737 12427
rect 13737 12393 13771 12427
rect 13771 12393 13780 12427
rect 13728 12384 13780 12393
rect 16396 12427 16448 12436
rect 16396 12393 16405 12427
rect 16405 12393 16439 12427
rect 16439 12393 16448 12427
rect 16396 12384 16448 12393
rect 18052 12384 18104 12436
rect 18512 12427 18564 12436
rect 18512 12393 18521 12427
rect 18521 12393 18555 12427
rect 18555 12393 18564 12427
rect 18512 12384 18564 12393
rect 22008 12384 22060 12436
rect 22192 12384 22244 12436
rect 22468 12384 22520 12436
rect 24124 12384 24176 12436
rect 3332 12316 3384 12368
rect 1492 12248 1544 12300
rect 2320 12248 2372 12300
rect 2872 12291 2924 12300
rect 2872 12257 2881 12291
rect 2881 12257 2915 12291
rect 2915 12257 2924 12291
rect 2872 12248 2924 12257
rect 2964 12248 3016 12300
rect 3884 12248 3936 12300
rect 4252 12248 4304 12300
rect 6276 12316 6328 12368
rect 9680 12316 9732 12368
rect 9772 12316 9824 12368
rect 10600 12359 10652 12368
rect 10600 12325 10609 12359
rect 10609 12325 10643 12359
rect 10643 12325 10652 12359
rect 10600 12316 10652 12325
rect 10876 12316 10928 12368
rect 12992 12316 13044 12368
rect 15384 12316 15436 12368
rect 16028 12359 16080 12368
rect 16028 12325 16037 12359
rect 16037 12325 16071 12359
rect 16071 12325 16080 12359
rect 16028 12316 16080 12325
rect 16212 12316 16264 12368
rect 16856 12316 16908 12368
rect 17408 12316 17460 12368
rect 18880 12316 18932 12368
rect 19616 12316 19668 12368
rect 20536 12316 20588 12368
rect 21180 12316 21232 12368
rect 22284 12316 22336 12368
rect 23204 12316 23256 12368
rect 6092 12291 6144 12300
rect 6092 12257 6101 12291
rect 6101 12257 6135 12291
rect 6135 12257 6144 12291
rect 6092 12248 6144 12257
rect 7012 12248 7064 12300
rect 8576 12291 8628 12300
rect 6828 12180 6880 12232
rect 8576 12257 8585 12291
rect 8585 12257 8619 12291
rect 8619 12257 8628 12291
rect 8576 12248 8628 12257
rect 9588 12248 9640 12300
rect 18144 12248 18196 12300
rect 22100 12291 22152 12300
rect 22100 12257 22109 12291
rect 22109 12257 22143 12291
rect 22143 12257 22152 12291
rect 22100 12248 22152 12257
rect 24584 12248 24636 12300
rect 25136 12248 25188 12300
rect 8944 12180 8996 12232
rect 12440 12180 12492 12232
rect 13084 12180 13136 12232
rect 14096 12180 14148 12232
rect 14740 12180 14792 12232
rect 17684 12180 17736 12232
rect 19340 12223 19392 12232
rect 19340 12189 19349 12223
rect 19349 12189 19383 12223
rect 19383 12189 19392 12223
rect 19340 12180 19392 12189
rect 20996 12180 21048 12232
rect 22744 12223 22796 12232
rect 22744 12189 22753 12223
rect 22753 12189 22787 12223
rect 22787 12189 22796 12223
rect 22744 12180 22796 12189
rect 23020 12223 23072 12232
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 23756 12180 23808 12232
rect 4712 12112 4764 12164
rect 10784 12112 10836 12164
rect 11060 12112 11112 12164
rect 20536 12112 20588 12164
rect 21180 12112 21232 12164
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 2412 12044 2464 12096
rect 4620 12044 4672 12096
rect 7104 12044 7156 12096
rect 8024 12044 8076 12096
rect 14096 12087 14148 12096
rect 14096 12053 14105 12087
rect 14105 12053 14139 12087
rect 14139 12053 14148 12087
rect 14096 12044 14148 12053
rect 19156 12044 19208 12096
rect 20260 12044 20312 12096
rect 20720 12087 20772 12096
rect 20720 12053 20729 12087
rect 20729 12053 20763 12087
rect 20763 12053 20772 12087
rect 20720 12044 20772 12053
rect 22100 12044 22152 12096
rect 23020 12044 23072 12096
rect 23664 12087 23716 12096
rect 23664 12053 23673 12087
rect 23673 12053 23707 12087
rect 23707 12053 23716 12087
rect 23664 12044 23716 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1492 11840 1544 11892
rect 2964 11840 3016 11892
rect 2044 11772 2096 11824
rect 1308 11704 1360 11756
rect 1492 11704 1544 11756
rect 1584 11704 1636 11756
rect 3608 11840 3660 11892
rect 3884 11883 3936 11892
rect 3884 11849 3893 11883
rect 3893 11849 3927 11883
rect 3927 11849 3936 11883
rect 3884 11840 3936 11849
rect 6276 11840 6328 11892
rect 6092 11815 6144 11824
rect 6092 11781 6101 11815
rect 6101 11781 6135 11815
rect 6135 11781 6144 11815
rect 8576 11840 8628 11892
rect 10600 11840 10652 11892
rect 8944 11815 8996 11824
rect 6092 11772 6144 11781
rect 8944 11781 8953 11815
rect 8953 11781 8987 11815
rect 8987 11781 8996 11815
rect 8944 11772 8996 11781
rect 17316 11840 17368 11892
rect 18880 11840 18932 11892
rect 21548 11840 21600 11892
rect 22284 11840 22336 11892
rect 25412 11883 25464 11892
rect 25412 11849 25421 11883
rect 25421 11849 25455 11883
rect 25455 11849 25464 11883
rect 25412 11840 25464 11849
rect 4528 11704 4580 11756
rect 7196 11704 7248 11756
rect 8668 11704 8720 11756
rect 9956 11704 10008 11756
rect 2320 11500 2372 11552
rect 4068 11636 4120 11688
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 11060 11636 11112 11688
rect 12532 11679 12584 11688
rect 12532 11645 12541 11679
rect 12541 11645 12575 11679
rect 12575 11645 12584 11679
rect 12532 11636 12584 11645
rect 12992 11679 13044 11688
rect 12992 11645 13001 11679
rect 13001 11645 13035 11679
rect 13035 11645 13044 11679
rect 15384 11704 15436 11756
rect 19616 11772 19668 11824
rect 23204 11772 23256 11824
rect 16028 11704 16080 11756
rect 17408 11704 17460 11756
rect 20720 11747 20772 11756
rect 20720 11713 20729 11747
rect 20729 11713 20763 11747
rect 20763 11713 20772 11747
rect 20720 11704 20772 11713
rect 20996 11704 21048 11756
rect 12992 11636 13044 11645
rect 14096 11679 14148 11688
rect 14096 11645 14105 11679
rect 14105 11645 14139 11679
rect 14139 11645 14148 11679
rect 14096 11636 14148 11645
rect 18880 11679 18932 11688
rect 5080 11611 5132 11620
rect 5080 11577 5089 11611
rect 5089 11577 5123 11611
rect 5123 11577 5132 11611
rect 5080 11568 5132 11577
rect 8024 11611 8076 11620
rect 8024 11577 8033 11611
rect 8033 11577 8067 11611
rect 8067 11577 8076 11611
rect 8024 11568 8076 11577
rect 9864 11568 9916 11620
rect 13268 11611 13320 11620
rect 3976 11500 4028 11552
rect 7012 11543 7064 11552
rect 7012 11509 7021 11543
rect 7021 11509 7055 11543
rect 7055 11509 7064 11543
rect 7012 11500 7064 11509
rect 7564 11500 7616 11552
rect 7748 11500 7800 11552
rect 9404 11543 9456 11552
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 10876 11543 10928 11552
rect 10876 11509 10885 11543
rect 10885 11509 10919 11543
rect 10919 11509 10928 11543
rect 10876 11500 10928 11509
rect 11520 11543 11572 11552
rect 11520 11509 11529 11543
rect 11529 11509 11563 11543
rect 11563 11509 11572 11543
rect 11520 11500 11572 11509
rect 13268 11577 13277 11611
rect 13277 11577 13311 11611
rect 13311 11577 13320 11611
rect 13268 11568 13320 11577
rect 13728 11500 13780 11552
rect 15292 11543 15344 11552
rect 15292 11509 15301 11543
rect 15301 11509 15335 11543
rect 15335 11509 15344 11543
rect 15292 11500 15344 11509
rect 18880 11645 18889 11679
rect 18889 11645 18923 11679
rect 18923 11645 18932 11679
rect 18880 11636 18932 11645
rect 22468 11679 22520 11688
rect 22468 11645 22512 11679
rect 22512 11645 22520 11679
rect 22468 11636 22520 11645
rect 23664 11636 23716 11688
rect 23848 11636 23900 11688
rect 25320 11636 25372 11688
rect 18972 11568 19024 11620
rect 20536 11611 20588 11620
rect 20536 11577 20545 11611
rect 20545 11577 20579 11611
rect 20579 11577 20588 11611
rect 20536 11568 20588 11577
rect 23296 11568 23348 11620
rect 24676 11611 24728 11620
rect 24676 11577 24685 11611
rect 24685 11577 24719 11611
rect 24719 11577 24728 11611
rect 24676 11568 24728 11577
rect 17684 11543 17736 11552
rect 17684 11509 17693 11543
rect 17693 11509 17727 11543
rect 17727 11509 17736 11543
rect 17684 11500 17736 11509
rect 20812 11500 20864 11552
rect 21364 11500 21416 11552
rect 22008 11500 22060 11552
rect 23204 11500 23256 11552
rect 23756 11543 23808 11552
rect 23756 11509 23765 11543
rect 23765 11509 23799 11543
rect 23799 11509 23808 11543
rect 23756 11500 23808 11509
rect 25136 11543 25188 11552
rect 25136 11509 25145 11543
rect 25145 11509 25179 11543
rect 25179 11509 25188 11543
rect 25136 11500 25188 11509
rect 25872 11500 25924 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 2872 11296 2924 11348
rect 4160 11296 4212 11348
rect 7196 11296 7248 11348
rect 8024 11296 8076 11348
rect 2504 11228 2556 11280
rect 4068 11228 4120 11280
rect 4252 11271 4304 11280
rect 4252 11237 4261 11271
rect 4261 11237 4295 11271
rect 4295 11237 4304 11271
rect 4252 11228 4304 11237
rect 1584 11160 1636 11212
rect 1768 11160 1820 11212
rect 2596 11160 2648 11212
rect 7104 11228 7156 11280
rect 7656 11228 7708 11280
rect 9404 11228 9456 11280
rect 10876 11271 10928 11280
rect 10876 11237 10885 11271
rect 10885 11237 10919 11271
rect 10919 11237 10928 11271
rect 10876 11228 10928 11237
rect 12532 11296 12584 11348
rect 13084 11339 13136 11348
rect 13084 11305 13093 11339
rect 13093 11305 13127 11339
rect 13127 11305 13136 11339
rect 13084 11296 13136 11305
rect 15292 11296 15344 11348
rect 18420 11296 18472 11348
rect 18880 11339 18932 11348
rect 18880 11305 18889 11339
rect 18889 11305 18923 11339
rect 18923 11305 18932 11339
rect 18880 11296 18932 11305
rect 20996 11339 21048 11348
rect 20996 11305 21005 11339
rect 21005 11305 21039 11339
rect 21039 11305 21048 11339
rect 20996 11296 21048 11305
rect 22744 11339 22796 11348
rect 22744 11305 22753 11339
rect 22753 11305 22787 11339
rect 22787 11305 22796 11339
rect 22744 11296 22796 11305
rect 23204 11296 23256 11348
rect 23848 11296 23900 11348
rect 24952 11339 25004 11348
rect 24952 11305 24961 11339
rect 24961 11305 24995 11339
rect 24995 11305 25004 11339
rect 24952 11296 25004 11305
rect 12808 11228 12860 11280
rect 13728 11271 13780 11280
rect 13728 11237 13731 11271
rect 13731 11237 13765 11271
rect 13765 11237 13780 11271
rect 13728 11228 13780 11237
rect 14832 11228 14884 11280
rect 15568 11271 15620 11280
rect 15568 11237 15577 11271
rect 15577 11237 15611 11271
rect 15611 11237 15620 11271
rect 15568 11228 15620 11237
rect 15660 11271 15712 11280
rect 15660 11237 15669 11271
rect 15669 11237 15703 11271
rect 15703 11237 15712 11271
rect 15660 11228 15712 11237
rect 17408 11228 17460 11280
rect 19340 11228 19392 11280
rect 20628 11228 20680 11280
rect 23388 11271 23440 11280
rect 23388 11237 23397 11271
rect 23397 11237 23431 11271
rect 23431 11237 23440 11271
rect 23388 11228 23440 11237
rect 23480 11271 23532 11280
rect 23480 11237 23489 11271
rect 23489 11237 23523 11271
rect 23523 11237 23532 11271
rect 23480 11228 23532 11237
rect 2320 11092 2372 11144
rect 2872 11135 2924 11144
rect 1584 11024 1636 11076
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 3700 11092 3752 11144
rect 4068 11092 4120 11144
rect 4620 11160 4672 11212
rect 5264 11160 5316 11212
rect 6368 11160 6420 11212
rect 4804 11092 4856 11144
rect 5540 11092 5592 11144
rect 8392 11160 8444 11212
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 12072 11160 12124 11212
rect 13268 11160 13320 11212
rect 14740 11160 14792 11212
rect 17316 11203 17368 11212
rect 17316 11169 17325 11203
rect 17325 11169 17359 11203
rect 17359 11169 17368 11203
rect 17316 11160 17368 11169
rect 19432 11203 19484 11212
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 19432 11160 19484 11169
rect 7196 11092 7248 11144
rect 11060 11135 11112 11144
rect 4528 11067 4580 11076
rect 4528 11033 4537 11067
rect 4537 11033 4571 11067
rect 4571 11033 4580 11067
rect 4528 11024 4580 11033
rect 9956 11024 10008 11076
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 11244 11092 11296 11144
rect 11428 11092 11480 11144
rect 12532 11092 12584 11144
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 19340 11092 19392 11144
rect 20536 11160 20588 11212
rect 23664 11135 23716 11144
rect 23664 11101 23673 11135
rect 23673 11101 23707 11135
rect 23707 11101 23716 11135
rect 23664 11092 23716 11101
rect 3700 10956 3752 11008
rect 21548 11024 21600 11076
rect 21916 11024 21968 11076
rect 23848 11024 23900 11076
rect 24952 11092 25004 11144
rect 25596 11024 25648 11076
rect 11244 10956 11296 11008
rect 11888 10956 11940 11008
rect 20444 10956 20496 11008
rect 20996 10956 21048 11008
rect 22284 10956 22336 11008
rect 23756 10956 23808 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1768 10752 1820 10804
rect 2596 10752 2648 10804
rect 2872 10752 2924 10804
rect 4804 10795 4856 10804
rect 4804 10761 4813 10795
rect 4813 10761 4847 10795
rect 4847 10761 4856 10795
rect 4804 10752 4856 10761
rect 5540 10795 5592 10804
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 6368 10752 6420 10804
rect 7196 10795 7248 10804
rect 7196 10761 7205 10795
rect 7205 10761 7239 10795
rect 7239 10761 7248 10795
rect 7196 10752 7248 10761
rect 7656 10795 7708 10804
rect 7656 10761 7665 10795
rect 7665 10761 7699 10795
rect 7699 10761 7708 10795
rect 7656 10752 7708 10761
rect 10876 10795 10928 10804
rect 10876 10761 10885 10795
rect 10885 10761 10919 10795
rect 10919 10761 10928 10795
rect 10876 10752 10928 10761
rect 11336 10752 11388 10804
rect 12808 10752 12860 10804
rect 13728 10752 13780 10804
rect 2320 10727 2372 10736
rect 2320 10693 2329 10727
rect 2329 10693 2363 10727
rect 2363 10693 2372 10727
rect 2320 10684 2372 10693
rect 2412 10616 2464 10668
rect 2504 10591 2556 10600
rect 2504 10557 2513 10591
rect 2513 10557 2547 10591
rect 2547 10557 2556 10591
rect 2504 10548 2556 10557
rect 4528 10548 4580 10600
rect 7288 10616 7340 10668
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 9680 10616 9732 10668
rect 12532 10659 12584 10668
rect 8484 10591 8536 10600
rect 8484 10557 8493 10591
rect 8493 10557 8527 10591
rect 8527 10557 8536 10591
rect 9312 10591 9364 10600
rect 8484 10548 8536 10557
rect 9312 10557 9321 10591
rect 9321 10557 9355 10591
rect 9355 10557 9364 10591
rect 9312 10548 9364 10557
rect 12532 10625 12541 10659
rect 12541 10625 12575 10659
rect 12575 10625 12584 10659
rect 12532 10616 12584 10625
rect 13360 10616 13412 10668
rect 13544 10616 13596 10668
rect 8024 10480 8076 10532
rect 9404 10480 9456 10532
rect 12624 10523 12676 10532
rect 12624 10489 12633 10523
rect 12633 10489 12667 10523
rect 12667 10489 12676 10523
rect 12624 10480 12676 10489
rect 13360 10480 13412 10532
rect 15384 10752 15436 10804
rect 15844 10795 15896 10804
rect 15844 10761 15853 10795
rect 15853 10761 15887 10795
rect 15887 10761 15896 10795
rect 15844 10752 15896 10761
rect 17040 10752 17092 10804
rect 18052 10752 18104 10804
rect 18696 10752 18748 10804
rect 21548 10795 21600 10804
rect 21548 10761 21557 10795
rect 21557 10761 21591 10795
rect 21591 10761 21600 10795
rect 21548 10752 21600 10761
rect 25320 10752 25372 10804
rect 17408 10727 17460 10736
rect 17408 10693 17417 10727
rect 17417 10693 17451 10727
rect 17451 10693 17460 10727
rect 17408 10684 17460 10693
rect 17960 10684 18012 10736
rect 14372 10548 14424 10600
rect 15844 10548 15896 10600
rect 18328 10616 18380 10668
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 21180 10616 21232 10668
rect 21364 10616 21416 10668
rect 20996 10591 21048 10600
rect 4252 10455 4304 10464
rect 4252 10421 4261 10455
rect 4261 10421 4295 10455
rect 4295 10421 4304 10455
rect 4252 10412 4304 10421
rect 4896 10412 4948 10464
rect 6092 10412 6144 10464
rect 10140 10412 10192 10464
rect 12072 10412 12124 10464
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 19432 10480 19484 10532
rect 20996 10557 21005 10591
rect 21005 10557 21039 10591
rect 21039 10557 21048 10591
rect 20996 10548 21048 10557
rect 20628 10480 20680 10532
rect 21180 10523 21232 10532
rect 21180 10489 21189 10523
rect 21189 10489 21223 10523
rect 21223 10489 21232 10523
rect 21180 10480 21232 10489
rect 22284 10591 22336 10600
rect 22284 10557 22293 10591
rect 22293 10557 22327 10591
rect 22327 10557 22336 10591
rect 22284 10548 22336 10557
rect 24492 10548 24544 10600
rect 23204 10480 23256 10532
rect 23756 10523 23808 10532
rect 23756 10489 23765 10523
rect 23765 10489 23799 10523
rect 23799 10489 23808 10523
rect 23756 10480 23808 10489
rect 18144 10455 18196 10464
rect 18144 10421 18153 10455
rect 18153 10421 18187 10455
rect 18187 10421 18196 10455
rect 18144 10412 18196 10421
rect 19340 10455 19392 10464
rect 19340 10421 19349 10455
rect 19349 10421 19383 10455
rect 19383 10421 19392 10455
rect 19340 10412 19392 10421
rect 20444 10412 20496 10464
rect 22100 10455 22152 10464
rect 22100 10421 22109 10455
rect 22109 10421 22143 10455
rect 22143 10421 22152 10455
rect 22100 10412 22152 10421
rect 22744 10412 22796 10464
rect 23480 10412 23532 10464
rect 24308 10412 24360 10464
rect 24676 10480 24728 10532
rect 24860 10480 24912 10532
rect 24952 10455 25004 10464
rect 24952 10421 24961 10455
rect 24961 10421 24995 10455
rect 24995 10421 25004 10455
rect 24952 10412 25004 10421
rect 25596 10412 25648 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 4620 10208 4672 10260
rect 5264 10251 5316 10260
rect 5264 10217 5273 10251
rect 5273 10217 5307 10251
rect 5307 10217 5316 10251
rect 5264 10208 5316 10217
rect 8024 10208 8076 10260
rect 11244 10251 11296 10260
rect 11244 10217 11253 10251
rect 11253 10217 11287 10251
rect 11287 10217 11296 10251
rect 11244 10208 11296 10217
rect 12348 10208 12400 10260
rect 12440 10208 12492 10260
rect 12624 10208 12676 10260
rect 13268 10208 13320 10260
rect 14372 10251 14424 10260
rect 14372 10217 14381 10251
rect 14381 10217 14415 10251
rect 14415 10217 14424 10251
rect 14372 10208 14424 10217
rect 14832 10208 14884 10260
rect 15200 10208 15252 10260
rect 15660 10208 15712 10260
rect 17316 10208 17368 10260
rect 18328 10251 18380 10260
rect 18328 10217 18337 10251
rect 18337 10217 18371 10251
rect 18371 10217 18380 10251
rect 18328 10208 18380 10217
rect 21088 10208 21140 10260
rect 21180 10208 21232 10260
rect 21824 10208 21876 10260
rect 23388 10251 23440 10260
rect 1768 10140 1820 10192
rect 2596 10140 2648 10192
rect 2320 10072 2372 10124
rect 2412 10115 2464 10124
rect 2412 10081 2421 10115
rect 2421 10081 2455 10115
rect 2455 10081 2464 10115
rect 2412 10072 2464 10081
rect 3884 10072 3936 10124
rect 4620 10072 4672 10124
rect 4804 10115 4856 10124
rect 4804 10081 4813 10115
rect 4813 10081 4847 10115
rect 4847 10081 4856 10115
rect 4804 10072 4856 10081
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 6368 10115 6420 10124
rect 9312 10183 9364 10192
rect 9312 10149 9321 10183
rect 9321 10149 9355 10183
rect 9355 10149 9364 10183
rect 9312 10140 9364 10149
rect 10140 10140 10192 10192
rect 10968 10183 11020 10192
rect 10968 10149 10977 10183
rect 10977 10149 11011 10183
rect 11011 10149 11020 10183
rect 10968 10140 11020 10149
rect 13176 10183 13228 10192
rect 13176 10149 13185 10183
rect 13185 10149 13219 10183
rect 13219 10149 13228 10183
rect 13176 10140 13228 10149
rect 17500 10183 17552 10192
rect 17500 10149 17509 10183
rect 17509 10149 17543 10183
rect 17543 10149 17552 10183
rect 17500 10140 17552 10149
rect 22008 10140 22060 10192
rect 22100 10140 22152 10192
rect 23388 10217 23397 10251
rect 23397 10217 23431 10251
rect 23431 10217 23440 10251
rect 23388 10208 23440 10217
rect 24860 10208 24912 10260
rect 24216 10140 24268 10192
rect 24492 10140 24544 10192
rect 6368 10081 6382 10115
rect 6382 10081 6416 10115
rect 6416 10081 6420 10115
rect 6368 10072 6420 10081
rect 7012 10072 7064 10124
rect 8024 10115 8076 10124
rect 8024 10081 8033 10115
rect 8033 10081 8067 10115
rect 8067 10081 8076 10115
rect 8024 10072 8076 10081
rect 8392 10072 8444 10124
rect 11796 10072 11848 10124
rect 12716 10072 12768 10124
rect 15752 10115 15804 10124
rect 1308 10004 1360 10056
rect 1584 10004 1636 10056
rect 1952 10004 2004 10056
rect 2596 10004 2648 10056
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 10048 10004 10100 10056
rect 13360 10047 13412 10056
rect 2412 9936 2464 9988
rect 4896 9979 4948 9988
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 1952 9911 2004 9920
rect 1952 9877 1961 9911
rect 1961 9877 1995 9911
rect 1995 9877 2004 9911
rect 1952 9868 2004 9877
rect 4896 9945 4905 9979
rect 4905 9945 4939 9979
rect 4939 9945 4948 9979
rect 4896 9936 4948 9945
rect 13360 10013 13369 10047
rect 13369 10013 13403 10047
rect 13403 10013 13412 10047
rect 13360 10004 13412 10013
rect 15752 10081 15761 10115
rect 15761 10081 15795 10115
rect 15795 10081 15804 10115
rect 15752 10072 15804 10081
rect 18880 10115 18932 10124
rect 18880 10081 18889 10115
rect 18889 10081 18923 10115
rect 18923 10081 18932 10115
rect 18880 10072 18932 10081
rect 20260 10072 20312 10124
rect 21456 10072 21508 10124
rect 21640 10072 21692 10124
rect 25228 10115 25280 10124
rect 25228 10081 25237 10115
rect 25237 10081 25271 10115
rect 25271 10081 25280 10115
rect 25228 10072 25280 10081
rect 15660 10004 15712 10056
rect 15844 10047 15896 10056
rect 15844 10013 15853 10047
rect 15853 10013 15887 10047
rect 15887 10013 15896 10047
rect 15844 10004 15896 10013
rect 17684 10004 17736 10056
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 19432 10047 19484 10056
rect 19432 10013 19441 10047
rect 19441 10013 19475 10047
rect 19475 10013 19484 10047
rect 19432 10004 19484 10013
rect 21916 10047 21968 10056
rect 21916 10013 21925 10047
rect 21925 10013 21959 10047
rect 21959 10013 21968 10047
rect 21916 10004 21968 10013
rect 23204 10004 23256 10056
rect 24032 10004 24084 10056
rect 3700 9868 3752 9920
rect 4252 9868 4304 9920
rect 13728 9936 13780 9988
rect 21456 9936 21508 9988
rect 22560 9936 22612 9988
rect 23664 9936 23716 9988
rect 23940 9936 23992 9988
rect 24308 9936 24360 9988
rect 16580 9868 16632 9920
rect 19248 9868 19300 9920
rect 20628 9868 20680 9920
rect 20720 9868 20772 9920
rect 21088 9868 21140 9920
rect 23388 9868 23440 9920
rect 23848 9868 23900 9920
rect 24032 9868 24084 9920
rect 25412 9911 25464 9920
rect 25412 9877 25421 9911
rect 25421 9877 25455 9911
rect 25455 9877 25464 9911
rect 25412 9868 25464 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2504 9664 2556 9716
rect 4344 9664 4396 9716
rect 4620 9664 4672 9716
rect 6368 9707 6420 9716
rect 6368 9673 6377 9707
rect 6377 9673 6411 9707
rect 6411 9673 6420 9707
rect 6368 9664 6420 9673
rect 8024 9707 8076 9716
rect 8024 9673 8033 9707
rect 8033 9673 8067 9707
rect 8067 9673 8076 9707
rect 8024 9664 8076 9673
rect 8392 9707 8444 9716
rect 8392 9673 8401 9707
rect 8401 9673 8435 9707
rect 8435 9673 8444 9707
rect 8392 9664 8444 9673
rect 10140 9664 10192 9716
rect 11796 9664 11848 9716
rect 13176 9664 13228 9716
rect 14004 9664 14056 9716
rect 1768 9639 1820 9648
rect 1768 9605 1792 9639
rect 1792 9605 1820 9639
rect 1768 9596 1820 9605
rect 2228 9639 2280 9648
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 2228 9605 2237 9639
rect 2237 9605 2271 9639
rect 2271 9605 2280 9639
rect 2228 9596 2280 9605
rect 2964 9639 3016 9648
rect 2964 9605 2973 9639
rect 2973 9605 3007 9639
rect 3007 9605 3016 9639
rect 2964 9596 3016 9605
rect 3148 9596 3200 9648
rect 10784 9639 10836 9648
rect 2136 9528 2188 9580
rect 1308 9460 1360 9512
rect 2228 9460 2280 9512
rect 10784 9605 10793 9639
rect 10793 9605 10827 9639
rect 10827 9605 10836 9639
rect 10784 9596 10836 9605
rect 5264 9571 5316 9580
rect 5264 9537 5273 9571
rect 5273 9537 5307 9571
rect 5307 9537 5316 9571
rect 5264 9528 5316 9537
rect 10232 9528 10284 9580
rect 13360 9571 13412 9580
rect 13360 9537 13369 9571
rect 13369 9537 13403 9571
rect 13403 9537 13412 9571
rect 13360 9528 13412 9537
rect 14280 9528 14332 9580
rect 15752 9664 15804 9716
rect 17500 9664 17552 9716
rect 17316 9596 17368 9648
rect 19340 9664 19392 9716
rect 20260 9707 20312 9716
rect 20260 9673 20269 9707
rect 20269 9673 20303 9707
rect 20303 9673 20312 9707
rect 20260 9664 20312 9673
rect 20996 9664 21048 9716
rect 22008 9664 22060 9716
rect 22744 9707 22796 9716
rect 22744 9673 22753 9707
rect 22753 9673 22787 9707
rect 22787 9673 22796 9707
rect 22744 9664 22796 9673
rect 24860 9664 24912 9716
rect 25320 9664 25372 9716
rect 19248 9571 19300 9580
rect 19248 9537 19257 9571
rect 19257 9537 19291 9571
rect 19291 9537 19300 9571
rect 19248 9528 19300 9537
rect 21824 9571 21876 9580
rect 21824 9537 21833 9571
rect 21833 9537 21867 9571
rect 21867 9537 21876 9571
rect 21824 9528 21876 9537
rect 23020 9528 23072 9580
rect 24032 9528 24084 9580
rect 24216 9571 24268 9580
rect 24216 9537 24225 9571
rect 24225 9537 24259 9571
rect 24259 9537 24268 9571
rect 24216 9528 24268 9537
rect 3608 9503 3660 9512
rect 3608 9469 3617 9503
rect 3617 9469 3651 9503
rect 3651 9469 3660 9503
rect 3608 9460 3660 9469
rect 4804 9503 4856 9512
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5080 9460 5132 9469
rect 6644 9460 6696 9512
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 7656 9460 7708 9512
rect 14832 9460 14884 9512
rect 17408 9460 17460 9512
rect 19064 9460 19116 9512
rect 1952 9392 2004 9444
rect 2872 9392 2924 9444
rect 4620 9435 4672 9444
rect 4620 9401 4629 9435
rect 4629 9401 4663 9435
rect 4663 9401 4672 9435
rect 4620 9392 4672 9401
rect 5264 9392 5316 9444
rect 3148 9324 3200 9376
rect 4344 9367 4396 9376
rect 4344 9333 4353 9367
rect 4353 9333 4387 9367
rect 4387 9333 4396 9367
rect 4344 9324 4396 9333
rect 7012 9367 7064 9376
rect 7012 9333 7021 9367
rect 7021 9333 7055 9367
rect 7055 9333 7064 9367
rect 7012 9324 7064 9333
rect 8760 9435 8812 9444
rect 8760 9401 8769 9435
rect 8769 9401 8803 9435
rect 8803 9401 8812 9435
rect 8760 9392 8812 9401
rect 9588 9392 9640 9444
rect 10232 9435 10284 9444
rect 10232 9401 10241 9435
rect 10241 9401 10275 9435
rect 10275 9401 10284 9435
rect 10232 9392 10284 9401
rect 9220 9324 9272 9376
rect 10140 9324 10192 9376
rect 13176 9435 13228 9444
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 13176 9392 13228 9401
rect 15568 9392 15620 9444
rect 13728 9324 13780 9376
rect 13820 9324 13872 9376
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 15384 9324 15436 9376
rect 15752 9324 15804 9376
rect 16396 9392 16448 9444
rect 17868 9392 17920 9444
rect 19340 9435 19392 9444
rect 19340 9401 19349 9435
rect 19349 9401 19383 9435
rect 19383 9401 19392 9435
rect 19340 9392 19392 9401
rect 20076 9392 20128 9444
rect 16488 9324 16540 9376
rect 17684 9367 17736 9376
rect 17684 9333 17693 9367
rect 17693 9333 17727 9367
rect 17727 9333 17736 9367
rect 17684 9324 17736 9333
rect 18880 9367 18932 9376
rect 18880 9333 18889 9367
rect 18889 9333 18923 9367
rect 18923 9333 18932 9367
rect 18880 9324 18932 9333
rect 20260 9324 20312 9376
rect 25228 9503 25280 9512
rect 25228 9469 25272 9503
rect 25272 9469 25280 9503
rect 25228 9460 25280 9469
rect 21640 9392 21692 9444
rect 22192 9435 22244 9444
rect 22192 9401 22195 9435
rect 22195 9401 22229 9435
rect 22229 9401 22244 9435
rect 22192 9392 22244 9401
rect 23848 9435 23900 9444
rect 23848 9401 23857 9435
rect 23857 9401 23891 9435
rect 23891 9401 23900 9435
rect 23848 9392 23900 9401
rect 21548 9367 21600 9376
rect 21548 9333 21557 9367
rect 21557 9333 21591 9367
rect 21591 9333 21600 9367
rect 21548 9324 21600 9333
rect 25136 9324 25188 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2688 9120 2740 9172
rect 2320 9095 2372 9104
rect 2320 9061 2329 9095
rect 2329 9061 2363 9095
rect 2363 9061 2372 9095
rect 2320 9052 2372 9061
rect 4804 9120 4856 9172
rect 10048 9120 10100 9172
rect 11980 9120 12032 9172
rect 16212 9120 16264 9172
rect 3884 9095 3936 9104
rect 2872 9027 2924 9036
rect 2872 8993 2881 9027
rect 2881 8993 2915 9027
rect 2915 8993 2924 9027
rect 2872 8984 2924 8993
rect 1768 8916 1820 8968
rect 2596 8916 2648 8968
rect 2688 8916 2740 8968
rect 3884 9061 3893 9095
rect 3893 9061 3927 9095
rect 3927 9061 3936 9095
rect 3884 9052 3936 9061
rect 7932 9095 7984 9104
rect 7932 9061 7935 9095
rect 7935 9061 7969 9095
rect 7969 9061 7984 9095
rect 7932 9052 7984 9061
rect 10140 9052 10192 9104
rect 12532 9052 12584 9104
rect 12808 9052 12860 9104
rect 13728 9095 13780 9104
rect 13728 9061 13737 9095
rect 13737 9061 13771 9095
rect 13771 9061 13780 9095
rect 13728 9052 13780 9061
rect 16120 9052 16172 9104
rect 17040 9052 17092 9104
rect 17500 9052 17552 9104
rect 17868 9120 17920 9172
rect 23848 9120 23900 9172
rect 18972 9095 19024 9104
rect 18972 9061 18975 9095
rect 18975 9061 19009 9095
rect 19009 9061 19024 9095
rect 18972 9052 19024 9061
rect 20996 9052 21048 9104
rect 21732 9052 21784 9104
rect 21824 9052 21876 9104
rect 22100 9052 22152 9104
rect 23020 9052 23072 9104
rect 23572 9052 23624 9104
rect 24860 9052 24912 9104
rect 4344 9027 4396 9036
rect 4344 8993 4353 9027
rect 4353 8993 4387 9027
rect 4387 8993 4396 9027
rect 5080 9027 5132 9036
rect 4344 8984 4396 8993
rect 5080 8993 5089 9027
rect 5089 8993 5123 9027
rect 5123 8993 5132 9027
rect 5080 8984 5132 8993
rect 6092 9027 6144 9036
rect 6092 8993 6101 9027
rect 6101 8993 6135 9027
rect 6135 8993 6144 9027
rect 6092 8984 6144 8993
rect 6460 8984 6512 9036
rect 7656 8984 7708 9036
rect 14464 8984 14516 9036
rect 17868 8984 17920 9036
rect 19432 8984 19484 9036
rect 23664 9027 23716 9036
rect 23664 8993 23673 9027
rect 23673 8993 23707 9027
rect 23707 8993 23716 9027
rect 23664 8984 23716 8993
rect 23848 9027 23900 9036
rect 23848 8993 23857 9027
rect 23857 8993 23891 9027
rect 23891 8993 23900 9027
rect 23848 8984 23900 8993
rect 8668 8916 8720 8968
rect 9864 8916 9916 8968
rect 2964 8848 3016 8900
rect 8944 8848 8996 8900
rect 9220 8891 9272 8900
rect 9220 8857 9229 8891
rect 9229 8857 9263 8891
rect 9263 8857 9272 8891
rect 9220 8848 9272 8857
rect 9404 8848 9456 8900
rect 11244 8916 11296 8968
rect 13176 8848 13228 8900
rect 13728 8848 13780 8900
rect 16212 8916 16264 8968
rect 16580 8916 16632 8968
rect 21732 8916 21784 8968
rect 19156 8848 19208 8900
rect 19432 8848 19484 8900
rect 21916 8848 21968 8900
rect 25044 8848 25096 8900
rect 25228 8848 25280 8900
rect 3608 8780 3660 8832
rect 3884 8780 3936 8832
rect 5264 8780 5316 8832
rect 7104 8823 7156 8832
rect 7104 8789 7113 8823
rect 7113 8789 7147 8823
rect 7147 8789 7156 8823
rect 7104 8780 7156 8789
rect 7656 8780 7708 8832
rect 8208 8780 8260 8832
rect 8576 8780 8628 8832
rect 8760 8823 8812 8832
rect 8760 8789 8769 8823
rect 8769 8789 8803 8823
rect 8803 8789 8812 8823
rect 8760 8780 8812 8789
rect 9772 8780 9824 8832
rect 14832 8780 14884 8832
rect 16120 8780 16172 8832
rect 16396 8823 16448 8832
rect 16396 8789 16405 8823
rect 16405 8789 16439 8823
rect 16439 8789 16448 8823
rect 16396 8780 16448 8789
rect 19340 8780 19392 8832
rect 21180 8823 21232 8832
rect 21180 8789 21189 8823
rect 21189 8789 21223 8823
rect 21223 8789 21232 8823
rect 21180 8780 21232 8789
rect 23204 8823 23256 8832
rect 23204 8789 23213 8823
rect 23213 8789 23247 8823
rect 23247 8789 23256 8823
rect 23204 8780 23256 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 4712 8576 4764 8628
rect 6092 8619 6144 8628
rect 1308 8508 1360 8560
rect 3056 8508 3108 8560
rect 2964 8440 3016 8492
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 3148 8415 3200 8424
rect 3148 8381 3157 8415
rect 3157 8381 3191 8415
rect 3191 8381 3200 8415
rect 3148 8372 3200 8381
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 6460 8619 6512 8628
rect 6460 8585 6469 8619
rect 6469 8585 6503 8619
rect 6503 8585 6512 8619
rect 6460 8576 6512 8585
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 8576 8576 8628 8628
rect 8668 8576 8720 8628
rect 8944 8576 8996 8628
rect 9496 8576 9548 8628
rect 11704 8576 11756 8628
rect 13268 8576 13320 8628
rect 14464 8576 14516 8628
rect 15568 8576 15620 8628
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17040 8576 17092 8585
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 19248 8576 19300 8628
rect 20260 8619 20312 8628
rect 20260 8585 20269 8619
rect 20269 8585 20303 8619
rect 20303 8585 20312 8619
rect 20260 8576 20312 8585
rect 20720 8576 20772 8628
rect 22100 8576 22152 8628
rect 22836 8576 22888 8628
rect 23848 8576 23900 8628
rect 24860 8576 24912 8628
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 12164 8508 12216 8560
rect 14372 8508 14424 8560
rect 19800 8551 19852 8560
rect 19800 8517 19809 8551
rect 19809 8517 19843 8551
rect 19843 8517 19852 8551
rect 19800 8508 19852 8517
rect 9588 8440 9640 8492
rect 15200 8440 15252 8492
rect 15844 8440 15896 8492
rect 17960 8440 18012 8492
rect 18972 8483 19024 8492
rect 18972 8449 18981 8483
rect 18981 8449 19015 8483
rect 19015 8449 19024 8483
rect 18972 8440 19024 8449
rect 23664 8508 23716 8560
rect 24768 8508 24820 8560
rect 21180 8440 21232 8492
rect 21824 8483 21876 8492
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 23572 8440 23624 8492
rect 24216 8483 24268 8492
rect 24216 8449 24225 8483
rect 24225 8449 24259 8483
rect 24259 8449 24268 8483
rect 24216 8440 24268 8449
rect 1492 8304 1544 8356
rect 3148 8236 3200 8288
rect 4252 8236 4304 8288
rect 4344 8279 4396 8288
rect 4344 8245 4353 8279
rect 4353 8245 4387 8279
rect 4387 8245 4396 8279
rect 4344 8236 4396 8245
rect 5172 8236 5224 8288
rect 11704 8372 11756 8424
rect 12992 8372 13044 8424
rect 13912 8372 13964 8424
rect 7932 8347 7984 8356
rect 7932 8313 7935 8347
rect 7935 8313 7969 8347
rect 7969 8313 7984 8347
rect 7932 8304 7984 8313
rect 9404 8347 9456 8356
rect 9404 8313 9413 8347
rect 9413 8313 9447 8347
rect 9447 8313 9456 8347
rect 9404 8304 9456 8313
rect 9496 8347 9548 8356
rect 9496 8313 9505 8347
rect 9505 8313 9539 8347
rect 9539 8313 9548 8347
rect 9496 8304 9548 8313
rect 9864 8304 9916 8356
rect 11244 8347 11296 8356
rect 11244 8313 11253 8347
rect 11253 8313 11287 8347
rect 11287 8313 11296 8347
rect 11244 8304 11296 8313
rect 10140 8236 10192 8288
rect 11704 8236 11756 8288
rect 12532 8304 12584 8356
rect 13636 8347 13688 8356
rect 13636 8313 13645 8347
rect 13645 8313 13679 8347
rect 13679 8313 13688 8347
rect 13636 8304 13688 8313
rect 16764 8372 16816 8424
rect 20720 8415 20772 8424
rect 20720 8381 20764 8415
rect 20764 8381 20772 8415
rect 20720 8372 20772 8381
rect 16580 8304 16632 8356
rect 19340 8347 19392 8356
rect 19340 8313 19349 8347
rect 19349 8313 19383 8347
rect 19383 8313 19392 8347
rect 19340 8304 19392 8313
rect 25044 8372 25096 8424
rect 25688 8415 25740 8424
rect 25688 8381 25697 8415
rect 25697 8381 25731 8415
rect 25731 8381 25740 8415
rect 25688 8372 25740 8381
rect 16120 8236 16172 8288
rect 21916 8236 21968 8288
rect 23848 8347 23900 8356
rect 23848 8313 23857 8347
rect 23857 8313 23891 8347
rect 23891 8313 23900 8347
rect 23848 8304 23900 8313
rect 23664 8236 23716 8288
rect 25228 8236 25280 8288
rect 26148 8236 26200 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2688 8032 2740 8084
rect 3700 8032 3752 8084
rect 2320 8007 2372 8016
rect 2320 7973 2329 8007
rect 2329 7973 2363 8007
rect 2363 7973 2372 8007
rect 2320 7964 2372 7973
rect 3516 7964 3568 8016
rect 4712 8032 4764 8084
rect 5172 8075 5224 8084
rect 5172 8041 5181 8075
rect 5181 8041 5215 8075
rect 5215 8041 5224 8075
rect 5172 8032 5224 8041
rect 5816 8075 5868 8084
rect 5816 8041 5825 8075
rect 5825 8041 5859 8075
rect 5859 8041 5868 8075
rect 5816 8032 5868 8041
rect 7748 8032 7800 8084
rect 7932 8032 7984 8084
rect 12348 8075 12400 8084
rect 4252 8007 4304 8016
rect 4252 7973 4261 8007
rect 4261 7973 4295 8007
rect 4295 7973 4304 8007
rect 4252 7964 4304 7973
rect 6276 7964 6328 8016
rect 8760 8007 8812 8016
rect 8760 7973 8769 8007
rect 8769 7973 8803 8007
rect 8803 7973 8812 8007
rect 8760 7964 8812 7973
rect 12348 8041 12357 8075
rect 12357 8041 12391 8075
rect 12391 8041 12400 8075
rect 12348 8032 12400 8041
rect 12992 8075 13044 8084
rect 12992 8041 13001 8075
rect 13001 8041 13035 8075
rect 13035 8041 13044 8075
rect 12992 8032 13044 8041
rect 13268 8032 13320 8084
rect 15108 8075 15160 8084
rect 11704 7964 11756 8016
rect 13728 8007 13780 8016
rect 13728 7973 13737 8007
rect 13737 7973 13771 8007
rect 13771 7973 13780 8007
rect 13728 7964 13780 7973
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 16120 8075 16172 8084
rect 16120 8041 16129 8075
rect 16129 8041 16163 8075
rect 16163 8041 16172 8075
rect 16120 8032 16172 8041
rect 17040 8032 17092 8084
rect 19340 8075 19392 8084
rect 16488 7964 16540 8016
rect 16764 7964 16816 8016
rect 19340 8041 19349 8075
rect 19349 8041 19383 8075
rect 19383 8041 19392 8075
rect 19340 8032 19392 8041
rect 23848 8032 23900 8084
rect 7932 7896 7984 7948
rect 1860 7828 1912 7880
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 2504 7760 2556 7812
rect 5448 7828 5500 7880
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 8300 7896 8352 7948
rect 8668 7896 8720 7948
rect 15568 7939 15620 7948
rect 15568 7905 15612 7939
rect 15612 7905 15620 7939
rect 15568 7896 15620 7905
rect 17408 7896 17460 7948
rect 21916 7964 21968 8016
rect 23664 7964 23716 8016
rect 18328 7939 18380 7948
rect 18328 7905 18337 7939
rect 18337 7905 18371 7939
rect 18371 7905 18380 7939
rect 18328 7896 18380 7905
rect 8760 7828 8812 7880
rect 9772 7828 9824 7880
rect 11244 7828 11296 7880
rect 14004 7871 14056 7880
rect 14004 7837 14013 7871
rect 14013 7837 14047 7871
rect 14047 7837 14056 7871
rect 14004 7828 14056 7837
rect 17316 7828 17368 7880
rect 25780 7896 25832 7948
rect 22008 7828 22060 7880
rect 25044 7828 25096 7880
rect 8024 7760 8076 7812
rect 14740 7760 14792 7812
rect 16672 7760 16724 7812
rect 21732 7760 21784 7812
rect 24216 7803 24268 7812
rect 24216 7769 24225 7803
rect 24225 7769 24259 7803
rect 24259 7769 24268 7803
rect 24216 7760 24268 7769
rect 1768 7692 1820 7744
rect 3608 7735 3660 7744
rect 3608 7701 3617 7735
rect 3617 7701 3651 7735
rect 3651 7701 3660 7735
rect 3608 7692 3660 7701
rect 5448 7735 5500 7744
rect 5448 7701 5457 7735
rect 5457 7701 5491 7735
rect 5491 7701 5500 7735
rect 5448 7692 5500 7701
rect 9404 7735 9456 7744
rect 9404 7701 9413 7735
rect 9413 7701 9447 7735
rect 9447 7701 9456 7735
rect 9404 7692 9456 7701
rect 9680 7692 9732 7744
rect 10140 7692 10192 7744
rect 11704 7692 11756 7744
rect 21824 7692 21876 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1676 7488 1728 7540
rect 2320 7488 2372 7540
rect 3884 7488 3936 7540
rect 4160 7488 4212 7540
rect 6276 7531 6328 7540
rect 6276 7497 6285 7531
rect 6285 7497 6319 7531
rect 6319 7497 6328 7531
rect 6276 7488 6328 7497
rect 8300 7488 8352 7540
rect 8852 7531 8904 7540
rect 8852 7497 8861 7531
rect 8861 7497 8895 7531
rect 8895 7497 8904 7531
rect 8852 7488 8904 7497
rect 11428 7488 11480 7540
rect 13268 7488 13320 7540
rect 15568 7488 15620 7540
rect 17684 7488 17736 7540
rect 18328 7531 18380 7540
rect 18328 7497 18337 7531
rect 18337 7497 18371 7531
rect 18371 7497 18380 7531
rect 22836 7531 22888 7540
rect 18328 7488 18380 7497
rect 10048 7420 10100 7472
rect 13636 7420 13688 7472
rect 4896 7352 4948 7404
rect 5448 7352 5500 7404
rect 6920 7352 6972 7404
rect 7932 7352 7984 7404
rect 9772 7352 9824 7404
rect 17316 7420 17368 7472
rect 19156 7420 19208 7472
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 19524 7352 19576 7404
rect 2504 7284 2556 7336
rect 3608 7284 3660 7336
rect 7104 7327 7156 7336
rect 7104 7293 7113 7327
rect 7113 7293 7147 7327
rect 7147 7293 7156 7327
rect 7104 7284 7156 7293
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 8852 7284 8904 7336
rect 11060 7284 11112 7336
rect 3240 7216 3292 7268
rect 6000 7216 6052 7268
rect 9588 7259 9640 7268
rect 9588 7225 9597 7259
rect 9597 7225 9631 7259
rect 9631 7225 9640 7259
rect 9588 7216 9640 7225
rect 9680 7259 9732 7268
rect 9680 7225 9689 7259
rect 9689 7225 9723 7259
rect 9723 7225 9732 7259
rect 15016 7284 15068 7336
rect 15384 7284 15436 7336
rect 15752 7327 15804 7336
rect 15752 7293 15761 7327
rect 15761 7293 15795 7327
rect 15795 7293 15804 7327
rect 15752 7284 15804 7293
rect 16856 7284 16908 7336
rect 22836 7497 22845 7531
rect 22845 7497 22879 7531
rect 22879 7497 22888 7531
rect 22836 7488 22888 7497
rect 25044 7531 25096 7540
rect 25044 7497 25053 7531
rect 25053 7497 25087 7531
rect 25087 7497 25096 7531
rect 25044 7488 25096 7497
rect 25136 7488 25188 7540
rect 25780 7531 25832 7540
rect 25780 7497 25789 7531
rect 25789 7497 25823 7531
rect 25823 7497 25832 7531
rect 25780 7488 25832 7497
rect 21824 7352 21876 7404
rect 24584 7352 24636 7404
rect 20260 7284 20312 7336
rect 20628 7327 20680 7336
rect 20628 7293 20637 7327
rect 20637 7293 20671 7327
rect 20671 7293 20680 7327
rect 20628 7284 20680 7293
rect 9680 7216 9732 7225
rect 6920 7191 6972 7200
rect 6920 7157 6929 7191
rect 6929 7157 6963 7191
rect 6963 7157 6972 7191
rect 6920 7148 6972 7157
rect 13452 7216 13504 7268
rect 13820 7259 13872 7268
rect 13820 7225 13829 7259
rect 13829 7225 13863 7259
rect 13863 7225 13872 7259
rect 13820 7216 13872 7225
rect 14004 7216 14056 7268
rect 18788 7259 18840 7268
rect 18788 7225 18797 7259
rect 18797 7225 18831 7259
rect 18831 7225 18840 7259
rect 18788 7216 18840 7225
rect 19064 7216 19116 7268
rect 22836 7284 22888 7336
rect 23388 7284 23440 7336
rect 11704 7191 11756 7200
rect 11704 7157 11713 7191
rect 11713 7157 11747 7191
rect 11747 7157 11756 7191
rect 11704 7148 11756 7157
rect 12624 7148 12676 7200
rect 12992 7191 13044 7200
rect 12992 7157 13001 7191
rect 13001 7157 13035 7191
rect 13035 7157 13044 7191
rect 12992 7148 13044 7157
rect 15016 7191 15068 7200
rect 15016 7157 15025 7191
rect 15025 7157 15059 7191
rect 15059 7157 15068 7191
rect 15016 7148 15068 7157
rect 15660 7148 15712 7200
rect 16764 7148 16816 7200
rect 17868 7148 17920 7200
rect 20168 7148 20220 7200
rect 21180 7191 21232 7200
rect 21180 7157 21189 7191
rect 21189 7157 21223 7191
rect 21223 7157 21232 7191
rect 21180 7148 21232 7157
rect 21732 7148 21784 7200
rect 23388 7191 23440 7200
rect 23388 7157 23397 7191
rect 23397 7157 23431 7191
rect 23431 7157 23440 7191
rect 23388 7148 23440 7157
rect 23756 7191 23808 7200
rect 23756 7157 23765 7191
rect 23765 7157 23799 7191
rect 23799 7157 23808 7191
rect 23756 7148 23808 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1216 6944 1268 6996
rect 4252 6944 4304 6996
rect 9772 6987 9824 6996
rect 9772 6953 9781 6987
rect 9781 6953 9815 6987
rect 9815 6953 9824 6987
rect 9772 6944 9824 6953
rect 13820 6944 13872 6996
rect 17408 6987 17460 6996
rect 17408 6953 17417 6987
rect 17417 6953 17451 6987
rect 17451 6953 17460 6987
rect 17408 6944 17460 6953
rect 18788 6987 18840 6996
rect 18788 6953 18797 6987
rect 18797 6953 18831 6987
rect 18831 6953 18840 6987
rect 18788 6944 18840 6953
rect 19524 6944 19576 6996
rect 20260 6987 20312 6996
rect 20260 6953 20269 6987
rect 20269 6953 20303 6987
rect 20303 6953 20312 6987
rect 20260 6944 20312 6953
rect 22744 6944 22796 6996
rect 23296 6944 23348 6996
rect 23664 6944 23716 6996
rect 25136 6987 25188 6996
rect 25136 6953 25145 6987
rect 25145 6953 25179 6987
rect 25179 6953 25188 6987
rect 25136 6944 25188 6953
rect 4896 6919 4948 6928
rect 4896 6885 4905 6919
rect 4905 6885 4939 6919
rect 4939 6885 4948 6919
rect 4896 6876 4948 6885
rect 6092 6919 6144 6928
rect 6092 6885 6095 6919
rect 6095 6885 6129 6919
rect 6129 6885 6144 6919
rect 7656 6919 7708 6928
rect 6092 6876 6144 6885
rect 7656 6885 7665 6919
rect 7665 6885 7699 6919
rect 7699 6885 7708 6919
rect 7656 6876 7708 6885
rect 9036 6876 9088 6928
rect 2872 6808 2924 6860
rect 3976 6808 4028 6860
rect 4528 6808 4580 6860
rect 4712 6851 4764 6860
rect 4712 6817 4721 6851
rect 4721 6817 4755 6851
rect 4755 6817 4764 6851
rect 4712 6808 4764 6817
rect 5540 6808 5592 6860
rect 9680 6851 9732 6860
rect 9680 6817 9689 6851
rect 9689 6817 9723 6851
rect 9723 6817 9732 6851
rect 15752 6876 15804 6928
rect 9680 6808 9732 6817
rect 10784 6808 10836 6860
rect 11612 6808 11664 6860
rect 12072 6808 12124 6860
rect 12440 6808 12492 6860
rect 14648 6808 14700 6860
rect 15292 6851 15344 6860
rect 15292 6817 15336 6851
rect 15336 6817 15344 6851
rect 15292 6808 15344 6817
rect 15476 6808 15528 6860
rect 16488 6851 16540 6860
rect 16488 6817 16497 6851
rect 16497 6817 16531 6851
rect 16531 6817 16540 6851
rect 16488 6808 16540 6817
rect 17868 6876 17920 6928
rect 21824 6876 21876 6928
rect 16764 6851 16816 6860
rect 16764 6817 16773 6851
rect 16773 6817 16807 6851
rect 16807 6817 16816 6851
rect 16764 6808 16816 6817
rect 19432 6808 19484 6860
rect 2688 6740 2740 6792
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 7288 6740 7340 6792
rect 7380 6740 7432 6792
rect 8024 6783 8076 6792
rect 8024 6749 8033 6783
rect 8033 6749 8067 6783
rect 8067 6749 8076 6783
rect 8024 6740 8076 6749
rect 8852 6783 8904 6792
rect 8852 6749 8861 6783
rect 8861 6749 8895 6783
rect 8895 6749 8904 6783
rect 8852 6740 8904 6749
rect 9588 6740 9640 6792
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 13084 6740 13136 6792
rect 18420 6740 18472 6792
rect 22376 6740 22428 6792
rect 1768 6604 1820 6656
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 2964 6604 3016 6656
rect 7656 6672 7708 6724
rect 9680 6672 9732 6724
rect 9956 6672 10008 6724
rect 10876 6672 10928 6724
rect 13176 6715 13228 6724
rect 13176 6681 13185 6715
rect 13185 6681 13219 6715
rect 13219 6681 13228 6715
rect 13176 6672 13228 6681
rect 24216 6808 24268 6860
rect 24676 6851 24728 6860
rect 24676 6817 24685 6851
rect 24685 6817 24719 6851
rect 24719 6817 24728 6851
rect 24676 6808 24728 6817
rect 24860 6851 24912 6860
rect 24860 6817 24869 6851
rect 24869 6817 24903 6851
rect 24903 6817 24912 6851
rect 24860 6808 24912 6817
rect 25320 6808 25372 6860
rect 25872 6808 25924 6860
rect 25596 6740 25648 6792
rect 3884 6604 3936 6656
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 8668 6604 8720 6656
rect 11244 6604 11296 6656
rect 13820 6604 13872 6656
rect 15752 6647 15804 6656
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 15752 6604 15804 6613
rect 16396 6604 16448 6656
rect 18144 6604 18196 6656
rect 21548 6604 21600 6656
rect 22008 6604 22060 6656
rect 23756 6604 23808 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2872 6400 2924 6452
rect 2964 6400 3016 6452
rect 4712 6443 4764 6452
rect 4712 6409 4721 6443
rect 4721 6409 4755 6443
rect 4755 6409 4764 6443
rect 4712 6400 4764 6409
rect 5540 6400 5592 6452
rect 7380 6443 7432 6452
rect 7380 6409 7389 6443
rect 7389 6409 7423 6443
rect 7423 6409 7432 6443
rect 7380 6400 7432 6409
rect 7656 6400 7708 6452
rect 9036 6443 9088 6452
rect 9036 6409 9045 6443
rect 9045 6409 9079 6443
rect 9079 6409 9088 6443
rect 9036 6400 9088 6409
rect 9312 6400 9364 6452
rect 9680 6400 9732 6452
rect 11612 6443 11664 6452
rect 11612 6409 11621 6443
rect 11621 6409 11655 6443
rect 11655 6409 11664 6443
rect 11612 6400 11664 6409
rect 12440 6400 12492 6452
rect 14648 6400 14700 6452
rect 15292 6400 15344 6452
rect 16488 6400 16540 6452
rect 16948 6400 17000 6452
rect 19432 6400 19484 6452
rect 22836 6400 22888 6452
rect 2688 6264 2740 6316
rect 3608 6264 3660 6316
rect 4896 6307 4948 6316
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 7012 6264 7064 6316
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 11244 6307 11296 6316
rect 11244 6273 11253 6307
rect 11253 6273 11287 6307
rect 11287 6273 11296 6307
rect 11244 6264 11296 6273
rect 2504 6196 2556 6248
rect 3976 6196 4028 6248
rect 4528 6196 4580 6248
rect 8208 6196 8260 6248
rect 10508 6239 10560 6248
rect 5172 6128 5224 6180
rect 6000 6060 6052 6112
rect 7932 6060 7984 6112
rect 9772 6060 9824 6112
rect 10140 6060 10192 6112
rect 10508 6205 10517 6239
rect 10517 6205 10551 6239
rect 10551 6205 10560 6239
rect 10508 6196 10560 6205
rect 10784 6196 10836 6248
rect 12808 6239 12860 6248
rect 12808 6205 12810 6239
rect 12810 6205 12860 6239
rect 16028 6332 16080 6384
rect 13820 6307 13872 6316
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 13820 6264 13872 6273
rect 14188 6307 14240 6316
rect 14188 6273 14197 6307
rect 14197 6273 14231 6307
rect 14231 6273 14240 6307
rect 14188 6264 14240 6273
rect 16396 6264 16448 6316
rect 16764 6307 16816 6316
rect 16764 6273 16773 6307
rect 16773 6273 16807 6307
rect 16807 6273 16816 6307
rect 23388 6332 23440 6384
rect 16764 6264 16816 6273
rect 12808 6196 12860 6205
rect 18144 6239 18196 6248
rect 13452 6060 13504 6112
rect 14648 6128 14700 6180
rect 15752 6128 15804 6180
rect 16212 6128 16264 6180
rect 18144 6205 18153 6239
rect 18153 6205 18187 6239
rect 18187 6205 18196 6239
rect 20168 6239 20220 6248
rect 18144 6196 18196 6205
rect 20168 6205 20177 6239
rect 20177 6205 20211 6239
rect 20211 6205 20220 6239
rect 20168 6196 20220 6205
rect 20444 6239 20496 6248
rect 20444 6205 20453 6239
rect 20453 6205 20487 6239
rect 20487 6205 20496 6239
rect 20444 6196 20496 6205
rect 21548 6239 21600 6248
rect 21548 6205 21557 6239
rect 21557 6205 21591 6239
rect 21591 6205 21600 6239
rect 21548 6196 21600 6205
rect 23388 6196 23440 6248
rect 23848 6196 23900 6248
rect 25228 6239 25280 6248
rect 25228 6205 25237 6239
rect 25237 6205 25271 6239
rect 25271 6205 25280 6239
rect 25228 6196 25280 6205
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 17868 6103 17920 6112
rect 17868 6069 17877 6103
rect 17877 6069 17911 6103
rect 17911 6069 17920 6103
rect 17868 6060 17920 6069
rect 19248 6060 19300 6112
rect 20720 6128 20772 6180
rect 20996 6128 21048 6180
rect 21088 6103 21140 6112
rect 21088 6069 21097 6103
rect 21097 6069 21131 6103
rect 21131 6069 21140 6103
rect 21824 6128 21876 6180
rect 21088 6060 21140 6069
rect 22468 6103 22520 6112
rect 22468 6069 22477 6103
rect 22477 6069 22511 6103
rect 22511 6069 22520 6103
rect 22468 6060 22520 6069
rect 23756 6103 23808 6112
rect 23756 6069 23765 6103
rect 23765 6069 23799 6103
rect 23799 6069 23808 6103
rect 23756 6060 23808 6069
rect 24860 6103 24912 6112
rect 24860 6069 24869 6103
rect 24869 6069 24903 6103
rect 24903 6069 24912 6103
rect 24860 6060 24912 6069
rect 26516 6060 26568 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1584 5856 1636 5908
rect 2504 5856 2556 5908
rect 5172 5856 5224 5908
rect 6276 5899 6328 5908
rect 6276 5865 6285 5899
rect 6285 5865 6319 5899
rect 6319 5865 6328 5899
rect 6276 5856 6328 5865
rect 6920 5899 6972 5908
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 7932 5899 7984 5908
rect 7932 5865 7941 5899
rect 7941 5865 7975 5899
rect 7975 5865 7984 5899
rect 7932 5856 7984 5865
rect 10968 5899 11020 5908
rect 10968 5865 10977 5899
rect 10977 5865 11011 5899
rect 11011 5865 11020 5899
rect 10968 5856 11020 5865
rect 13452 5899 13504 5908
rect 13452 5865 13461 5899
rect 13461 5865 13495 5899
rect 13495 5865 13504 5899
rect 13452 5856 13504 5865
rect 3792 5788 3844 5840
rect 4528 5788 4580 5840
rect 6000 5788 6052 5840
rect 1124 5720 1176 5772
rect 2320 5720 2372 5772
rect 2504 5720 2556 5772
rect 7564 5788 7616 5840
rect 13084 5831 13136 5840
rect 13084 5797 13093 5831
rect 13093 5797 13127 5831
rect 13127 5797 13136 5831
rect 13084 5788 13136 5797
rect 18420 5899 18472 5908
rect 18420 5865 18429 5899
rect 18429 5865 18463 5899
rect 18463 5865 18472 5899
rect 18420 5856 18472 5865
rect 20168 5856 20220 5908
rect 20996 5899 21048 5908
rect 20996 5865 21005 5899
rect 21005 5865 21039 5899
rect 21039 5865 21048 5899
rect 20996 5856 21048 5865
rect 23480 5856 23532 5908
rect 23756 5856 23808 5908
rect 24216 5899 24268 5908
rect 24216 5865 24225 5899
rect 24225 5865 24259 5899
rect 24259 5865 24268 5899
rect 24216 5856 24268 5865
rect 25320 5856 25372 5908
rect 13820 5831 13872 5840
rect 13820 5797 13829 5831
rect 13829 5797 13863 5831
rect 13863 5797 13872 5831
rect 13820 5788 13872 5797
rect 15568 5788 15620 5840
rect 17224 5831 17276 5840
rect 17224 5797 17233 5831
rect 17233 5797 17267 5831
rect 17267 5797 17276 5831
rect 17224 5788 17276 5797
rect 18972 5831 19024 5840
rect 18972 5797 18981 5831
rect 18981 5797 19015 5831
rect 19015 5797 19024 5831
rect 18972 5788 19024 5797
rect 19248 5788 19300 5840
rect 20444 5788 20496 5840
rect 22468 5788 22520 5840
rect 23940 5788 23992 5840
rect 24308 5788 24360 5840
rect 7748 5720 7800 5772
rect 12072 5763 12124 5772
rect 12072 5729 12081 5763
rect 12081 5729 12115 5763
rect 12115 5729 12124 5763
rect 12072 5720 12124 5729
rect 12624 5763 12676 5772
rect 12624 5729 12633 5763
rect 12633 5729 12667 5763
rect 12667 5729 12676 5763
rect 12624 5720 12676 5729
rect 14740 5763 14792 5772
rect 14740 5729 14749 5763
rect 14749 5729 14783 5763
rect 14783 5729 14792 5763
rect 14740 5720 14792 5729
rect 20536 5720 20588 5772
rect 20904 5763 20956 5772
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 21364 5763 21416 5772
rect 21364 5729 21373 5763
rect 21373 5729 21407 5763
rect 21407 5729 21416 5763
rect 21364 5720 21416 5729
rect 23848 5720 23900 5772
rect 2688 5652 2740 5704
rect 3976 5652 4028 5704
rect 4068 5652 4120 5704
rect 5908 5695 5960 5704
rect 5908 5661 5917 5695
rect 5917 5661 5951 5695
rect 5951 5661 5960 5695
rect 5908 5652 5960 5661
rect 6920 5652 6972 5704
rect 8208 5652 8260 5704
rect 9772 5652 9824 5704
rect 10508 5652 10560 5704
rect 14832 5652 14884 5704
rect 22652 5695 22704 5704
rect 2872 5584 2924 5636
rect 9680 5584 9732 5636
rect 14188 5584 14240 5636
rect 17040 5584 17092 5636
rect 22652 5661 22661 5695
rect 22661 5661 22695 5695
rect 22695 5661 22704 5695
rect 22652 5652 22704 5661
rect 24216 5720 24268 5772
rect 24676 5652 24728 5704
rect 17316 5584 17368 5636
rect 19156 5584 19208 5636
rect 19524 5627 19576 5636
rect 19524 5593 19533 5627
rect 19533 5593 19567 5627
rect 19567 5593 19576 5627
rect 19524 5584 19576 5593
rect 2228 5559 2280 5568
rect 2228 5525 2237 5559
rect 2237 5525 2271 5559
rect 2271 5525 2280 5559
rect 2228 5516 2280 5525
rect 2688 5559 2740 5568
rect 2688 5525 2697 5559
rect 2697 5525 2731 5559
rect 2731 5525 2740 5559
rect 2688 5516 2740 5525
rect 3332 5516 3384 5568
rect 3792 5516 3844 5568
rect 4160 5516 4212 5568
rect 9864 5516 9916 5568
rect 10416 5516 10468 5568
rect 10784 5516 10836 5568
rect 10876 5516 10928 5568
rect 17868 5516 17920 5568
rect 21916 5559 21968 5568
rect 21916 5525 21925 5559
rect 21925 5525 21959 5559
rect 21959 5525 21968 5559
rect 21916 5516 21968 5525
rect 22376 5559 22428 5568
rect 22376 5525 22385 5559
rect 22385 5525 22419 5559
rect 22419 5525 22428 5559
rect 22376 5516 22428 5525
rect 23388 5516 23440 5568
rect 24216 5516 24268 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2228 5312 2280 5364
rect 2412 5312 2464 5364
rect 4528 5312 4580 5364
rect 6920 5312 6972 5364
rect 8392 5355 8444 5364
rect 8392 5321 8401 5355
rect 8401 5321 8435 5355
rect 8435 5321 8444 5355
rect 8392 5312 8444 5321
rect 9772 5312 9824 5364
rect 10968 5312 11020 5364
rect 11152 5355 11204 5364
rect 11152 5321 11161 5355
rect 11161 5321 11195 5355
rect 11195 5321 11204 5355
rect 11152 5312 11204 5321
rect 12072 5355 12124 5364
rect 12072 5321 12081 5355
rect 12081 5321 12115 5355
rect 12115 5321 12124 5355
rect 12072 5312 12124 5321
rect 12624 5312 12676 5364
rect 14004 5312 14056 5364
rect 14648 5312 14700 5364
rect 17224 5355 17276 5364
rect 17224 5321 17233 5355
rect 17233 5321 17267 5355
rect 17267 5321 17276 5355
rect 17224 5312 17276 5321
rect 19248 5312 19300 5364
rect 2136 5244 2188 5296
rect 2780 5244 2832 5296
rect 2320 5176 2372 5228
rect 2964 5176 3016 5228
rect 10140 5244 10192 5296
rect 10416 5244 10468 5296
rect 19340 5287 19392 5296
rect 19340 5253 19349 5287
rect 19349 5253 19383 5287
rect 19383 5253 19392 5287
rect 19340 5244 19392 5253
rect 4068 5176 4120 5228
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 10508 5176 10560 5228
rect 14740 5176 14792 5228
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 2136 5108 2188 5160
rect 2504 5040 2556 5092
rect 2872 5083 2924 5092
rect 2872 5049 2881 5083
rect 2881 5049 2915 5083
rect 2915 5049 2924 5083
rect 2872 5040 2924 5049
rect 4712 5108 4764 5160
rect 6000 5108 6052 5160
rect 6920 5108 6972 5160
rect 3884 5040 3936 5092
rect 5172 5040 5224 5092
rect 5632 5040 5684 5092
rect 7748 5108 7800 5160
rect 8392 5108 8444 5160
rect 8668 5108 8720 5160
rect 12532 5108 12584 5160
rect 19248 5108 19300 5160
rect 21272 5312 21324 5364
rect 22652 5312 22704 5364
rect 23296 5312 23348 5364
rect 24676 5355 24728 5364
rect 21916 5176 21968 5228
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 24216 5151 24268 5160
rect 24216 5117 24225 5151
rect 24225 5117 24259 5151
rect 24259 5117 24268 5151
rect 24216 5108 24268 5117
rect 25228 5151 25280 5160
rect 25228 5117 25237 5151
rect 25237 5117 25271 5151
rect 25271 5117 25280 5151
rect 25228 5108 25280 5117
rect 7472 5040 7524 5092
rect 8024 5083 8076 5092
rect 8024 5049 8033 5083
rect 8033 5049 8067 5083
rect 8067 5049 8076 5083
rect 8024 5040 8076 5049
rect 8208 5040 8260 5092
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 10048 5040 10100 5092
rect 10876 5040 10928 5092
rect 18328 5083 18380 5092
rect 9680 5015 9732 5024
rect 9680 4981 9689 5015
rect 9689 4981 9723 5015
rect 9723 4981 9732 5015
rect 9680 4972 9732 4981
rect 9956 5015 10008 5024
rect 9956 4981 9965 5015
rect 9965 4981 9999 5015
rect 9999 4981 10008 5015
rect 9956 4972 10008 4981
rect 10784 4972 10836 5024
rect 11428 4972 11480 5024
rect 11704 4972 11756 5024
rect 15660 4972 15712 5024
rect 18328 5049 18337 5083
rect 18337 5049 18371 5083
rect 18371 5049 18380 5083
rect 18328 5040 18380 5049
rect 18420 5083 18472 5092
rect 18420 5049 18438 5083
rect 18438 5049 18472 5083
rect 18420 5040 18472 5049
rect 22376 5083 22428 5092
rect 22376 5049 22385 5083
rect 22385 5049 22419 5083
rect 22419 5049 22428 5083
rect 22376 5040 22428 5049
rect 16580 5015 16632 5024
rect 16580 4981 16589 5015
rect 16589 4981 16623 5015
rect 16623 4981 16632 5015
rect 16580 4972 16632 4981
rect 17500 4972 17552 5024
rect 20260 5015 20312 5024
rect 20260 4981 20269 5015
rect 20269 4981 20303 5015
rect 20303 4981 20312 5015
rect 20260 4972 20312 4981
rect 21088 5015 21140 5024
rect 21088 4981 21097 5015
rect 21097 4981 21131 5015
rect 21131 4981 21140 5015
rect 21088 4972 21140 4981
rect 22100 5015 22152 5024
rect 22100 4981 22109 5015
rect 22109 4981 22143 5015
rect 22143 4981 22152 5015
rect 22100 4972 22152 4981
rect 23480 4972 23532 5024
rect 25504 4972 25556 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1860 4768 1912 4820
rect 2780 4768 2832 4820
rect 2964 4768 3016 4820
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 4160 4768 4212 4820
rect 4712 4811 4764 4820
rect 4712 4777 4721 4811
rect 4721 4777 4755 4811
rect 4755 4777 4764 4811
rect 4712 4768 4764 4777
rect 6920 4811 6972 4820
rect 6920 4777 6929 4811
rect 6929 4777 6963 4811
rect 6963 4777 6972 4811
rect 6920 4768 6972 4777
rect 8576 4811 8628 4820
rect 8576 4777 8585 4811
rect 8585 4777 8619 4811
rect 8619 4777 8628 4811
rect 8576 4768 8628 4777
rect 9036 4811 9088 4820
rect 9036 4777 9045 4811
rect 9045 4777 9079 4811
rect 9079 4777 9088 4811
rect 9036 4768 9088 4777
rect 10784 4811 10836 4820
rect 10784 4777 10793 4811
rect 10793 4777 10827 4811
rect 10827 4777 10836 4811
rect 10784 4768 10836 4777
rect 10968 4768 11020 4820
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 13820 4768 13872 4820
rect 14832 4768 14884 4820
rect 17592 4768 17644 4820
rect 18236 4768 18288 4820
rect 18328 4768 18380 4820
rect 20352 4768 20404 4820
rect 22468 4768 22520 4820
rect 1124 4700 1176 4752
rect 3240 4700 3292 4752
rect 5080 4743 5132 4752
rect 5080 4709 5089 4743
rect 5089 4709 5123 4743
rect 5123 4709 5132 4743
rect 5080 4700 5132 4709
rect 5632 4743 5684 4752
rect 5632 4709 5641 4743
rect 5641 4709 5675 4743
rect 5675 4709 5684 4743
rect 7288 4743 7340 4752
rect 5632 4700 5684 4709
rect 7288 4709 7297 4743
rect 7297 4709 7331 4743
rect 7331 4709 7340 4743
rect 7288 4700 7340 4709
rect 7748 4700 7800 4752
rect 9864 4700 9916 4752
rect 10692 4700 10744 4752
rect 13636 4743 13688 4752
rect 13636 4709 13645 4743
rect 13645 4709 13679 4743
rect 13679 4709 13688 4743
rect 13636 4700 13688 4709
rect 14188 4743 14240 4752
rect 14188 4709 14197 4743
rect 14197 4709 14231 4743
rect 14231 4709 14240 4743
rect 14188 4700 14240 4709
rect 16120 4700 16172 4752
rect 16580 4700 16632 4752
rect 17316 4700 17368 4752
rect 18420 4743 18472 4752
rect 18420 4709 18429 4743
rect 18429 4709 18463 4743
rect 18463 4709 18472 4743
rect 18420 4700 18472 4709
rect 21088 4700 21140 4752
rect 22100 4700 22152 4752
rect 22652 4700 22704 4752
rect 23388 4700 23440 4752
rect 23940 4700 23992 4752
rect 24216 4700 24268 4752
rect 2228 4632 2280 4684
rect 2504 4632 2556 4684
rect 3332 4632 3384 4684
rect 6736 4632 6788 4684
rect 9404 4675 9456 4684
rect 9404 4641 9413 4675
rect 9413 4641 9447 4675
rect 9447 4641 9456 4675
rect 9404 4632 9456 4641
rect 11520 4675 11572 4684
rect 11520 4641 11529 4675
rect 11529 4641 11563 4675
rect 11563 4641 11572 4675
rect 11520 4632 11572 4641
rect 12164 4632 12216 4684
rect 17500 4632 17552 4684
rect 19708 4632 19760 4684
rect 20628 4632 20680 4684
rect 24768 4632 24820 4684
rect 2872 4564 2924 4616
rect 4436 4564 4488 4616
rect 7472 4564 7524 4616
rect 2688 4539 2740 4548
rect 2688 4505 2697 4539
rect 2697 4505 2731 4539
rect 2731 4505 2740 4539
rect 2688 4496 2740 4505
rect 10784 4496 10836 4548
rect 16212 4564 16264 4616
rect 18328 4607 18380 4616
rect 18328 4573 18337 4607
rect 18337 4573 18371 4607
rect 18371 4573 18380 4607
rect 18328 4564 18380 4573
rect 18972 4607 19024 4616
rect 18972 4573 18981 4607
rect 18981 4573 19015 4607
rect 19015 4573 19024 4607
rect 18972 4564 19024 4573
rect 21180 4564 21232 4616
rect 23020 4564 23072 4616
rect 24952 4607 25004 4616
rect 24952 4573 24961 4607
rect 24961 4573 24995 4607
rect 24995 4573 25004 4607
rect 24952 4564 25004 4573
rect 21364 4496 21416 4548
rect 22192 4496 22244 4548
rect 2596 4471 2648 4480
rect 2596 4437 2620 4471
rect 2620 4437 2648 4471
rect 2596 4428 2648 4437
rect 3332 4428 3384 4480
rect 8944 4428 8996 4480
rect 9680 4428 9732 4480
rect 11152 4428 11204 4480
rect 13268 4471 13320 4480
rect 13268 4437 13277 4471
rect 13277 4437 13311 4471
rect 13311 4437 13320 4471
rect 13268 4428 13320 4437
rect 15660 4471 15712 4480
rect 15660 4437 15669 4471
rect 15669 4437 15703 4471
rect 15703 4437 15712 4471
rect 15660 4428 15712 4437
rect 17040 4471 17092 4480
rect 17040 4437 17049 4471
rect 17049 4437 17083 4471
rect 17083 4437 17092 4471
rect 17040 4428 17092 4437
rect 19340 4428 19392 4480
rect 22008 4471 22060 4480
rect 22008 4437 22017 4471
rect 22017 4437 22051 4471
rect 22051 4437 22060 4471
rect 22008 4428 22060 4437
rect 24216 4471 24268 4480
rect 24216 4437 24225 4471
rect 24225 4437 24259 4471
rect 24259 4437 24268 4471
rect 24216 4428 24268 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1952 4267 2004 4276
rect 1952 4233 1961 4267
rect 1961 4233 1995 4267
rect 1995 4233 2004 4267
rect 1952 4224 2004 4233
rect 2872 4267 2924 4276
rect 2872 4233 2881 4267
rect 2881 4233 2915 4267
rect 2915 4233 2924 4267
rect 2872 4224 2924 4233
rect 3332 4267 3384 4276
rect 3332 4233 3341 4267
rect 3341 4233 3375 4267
rect 3375 4233 3384 4267
rect 3332 4224 3384 4233
rect 5356 4224 5408 4276
rect 7748 4224 7800 4276
rect 9680 4267 9732 4276
rect 9680 4233 9689 4267
rect 9689 4233 9723 4267
rect 9723 4233 9732 4267
rect 9680 4224 9732 4233
rect 10048 4267 10100 4276
rect 10048 4233 10057 4267
rect 10057 4233 10091 4267
rect 10091 4233 10100 4267
rect 10048 4224 10100 4233
rect 10784 4267 10836 4276
rect 10784 4233 10793 4267
rect 10793 4233 10827 4267
rect 10827 4233 10836 4267
rect 10784 4224 10836 4233
rect 11520 4224 11572 4276
rect 12164 4267 12216 4276
rect 12164 4233 12173 4267
rect 12173 4233 12207 4267
rect 12207 4233 12216 4267
rect 12164 4224 12216 4233
rect 16120 4267 16172 4276
rect 16120 4233 16129 4267
rect 16129 4233 16163 4267
rect 16163 4233 16172 4267
rect 16120 4224 16172 4233
rect 17500 4267 17552 4276
rect 17500 4233 17509 4267
rect 17509 4233 17543 4267
rect 17543 4233 17552 4267
rect 17500 4224 17552 4233
rect 18420 4224 18472 4276
rect 19708 4267 19760 4276
rect 19708 4233 19717 4267
rect 19717 4233 19751 4267
rect 19751 4233 19760 4267
rect 19708 4224 19760 4233
rect 22008 4224 22060 4276
rect 24768 4267 24820 4276
rect 24768 4233 24777 4267
rect 24777 4233 24811 4267
rect 24811 4233 24820 4267
rect 24768 4224 24820 4233
rect 6736 4156 6788 4208
rect 5080 4088 5132 4140
rect 9404 4156 9456 4208
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 7656 4088 7708 4140
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8944 4131 8996 4140
rect 8300 4088 8352 4097
rect 1492 4020 1544 4072
rect 2688 4020 2740 4072
rect 3148 4020 3200 4072
rect 3700 4020 3752 4072
rect 4252 4020 4304 4072
rect 4712 4020 4764 4072
rect 8944 4097 8953 4131
rect 8953 4097 8987 4131
rect 8987 4097 8996 4131
rect 8944 4088 8996 4097
rect 9036 4088 9088 4140
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 8576 4063 8628 4072
rect 4160 3995 4212 4004
rect 4160 3961 4169 3995
rect 4169 3961 4203 3995
rect 4203 3961 4212 3995
rect 4160 3952 4212 3961
rect 4804 3952 4856 4004
rect 4436 3927 4488 3936
rect 4436 3893 4445 3927
rect 4445 3893 4479 3927
rect 4479 3893 4488 3927
rect 4436 3884 4488 3893
rect 5540 3952 5592 4004
rect 6920 3952 6972 4004
rect 8576 4029 8585 4063
rect 8585 4029 8619 4063
rect 8619 4029 8628 4063
rect 8576 4020 8628 4029
rect 9680 4020 9732 4072
rect 11336 4063 11388 4072
rect 11336 4029 11345 4063
rect 11345 4029 11379 4063
rect 11379 4029 11388 4063
rect 13084 4088 13136 4140
rect 15384 4156 15436 4208
rect 14372 4088 14424 4140
rect 16212 4156 16264 4208
rect 15844 4088 15896 4140
rect 16304 4088 16356 4140
rect 17592 4156 17644 4208
rect 19248 4088 19300 4140
rect 19984 4088 20036 4140
rect 20168 4156 20220 4208
rect 25320 4156 25372 4208
rect 11336 4020 11388 4029
rect 18144 4020 18196 4072
rect 23388 4088 23440 4140
rect 22836 4020 22888 4072
rect 6092 3884 6144 3936
rect 9128 3952 9180 4004
rect 15384 3995 15436 4004
rect 7380 3884 7432 3936
rect 11428 3884 11480 3936
rect 12624 3927 12676 3936
rect 12624 3893 12633 3927
rect 12633 3893 12667 3927
rect 12667 3893 12676 3927
rect 12624 3884 12676 3893
rect 13636 3884 13688 3936
rect 15384 3961 15393 3995
rect 15393 3961 15427 3995
rect 15427 3961 15436 3995
rect 15384 3952 15436 3961
rect 16580 3995 16632 4004
rect 16580 3961 16589 3995
rect 16589 3961 16623 3995
rect 16623 3961 16632 3995
rect 16580 3952 16632 3961
rect 17868 3927 17920 3936
rect 17868 3893 17877 3927
rect 17877 3893 17911 3927
rect 17911 3893 17920 3927
rect 20536 3995 20588 4004
rect 20536 3961 20545 3995
rect 20545 3961 20579 3995
rect 20579 3961 20588 3995
rect 20536 3952 20588 3961
rect 21456 3952 21508 4004
rect 22100 3995 22152 4004
rect 22100 3961 22109 3995
rect 22109 3961 22143 3995
rect 22143 3961 22152 3995
rect 23756 4020 23808 4072
rect 24216 4020 24268 4072
rect 24952 4020 25004 4072
rect 25688 4088 25740 4140
rect 22100 3952 22152 3961
rect 19248 3927 19300 3936
rect 17868 3884 17920 3893
rect 19248 3893 19257 3927
rect 19257 3893 19291 3927
rect 19291 3893 19300 3927
rect 19248 3884 19300 3893
rect 21088 3927 21140 3936
rect 21088 3893 21097 3927
rect 21097 3893 21131 3927
rect 21131 3893 21140 3927
rect 21088 3884 21140 3893
rect 23756 3927 23808 3936
rect 23756 3893 23765 3927
rect 23765 3893 23799 3927
rect 23799 3893 23808 3927
rect 23756 3884 23808 3893
rect 25596 3884 25648 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2228 3723 2280 3732
rect 2228 3689 2237 3723
rect 2237 3689 2271 3723
rect 2271 3689 2280 3723
rect 2228 3680 2280 3689
rect 2688 3680 2740 3732
rect 2780 3680 2832 3732
rect 3700 3680 3752 3732
rect 4252 3723 4304 3732
rect 4252 3689 4261 3723
rect 4261 3689 4295 3723
rect 4295 3689 4304 3723
rect 4252 3680 4304 3689
rect 5080 3680 5132 3732
rect 6368 3723 6420 3732
rect 6368 3689 6377 3723
rect 6377 3689 6411 3723
rect 6411 3689 6420 3723
rect 6368 3680 6420 3689
rect 7288 3680 7340 3732
rect 9404 3723 9456 3732
rect 9404 3689 9413 3723
rect 9413 3689 9447 3723
rect 9447 3689 9456 3723
rect 9404 3680 9456 3689
rect 9680 3680 9732 3732
rect 10140 3680 10192 3732
rect 4804 3655 4856 3664
rect 4804 3621 4807 3655
rect 4807 3621 4841 3655
rect 4841 3621 4856 3655
rect 4804 3612 4856 3621
rect 7380 3655 7432 3664
rect 7380 3621 7389 3655
rect 7389 3621 7423 3655
rect 7423 3621 7432 3655
rect 7380 3612 7432 3621
rect 7748 3612 7800 3664
rect 9220 3612 9272 3664
rect 10048 3612 10100 3664
rect 1492 3587 1544 3596
rect 1492 3553 1510 3587
rect 1510 3553 1544 3587
rect 1492 3544 1544 3553
rect 2872 3587 2924 3596
rect 2872 3553 2881 3587
rect 2881 3553 2915 3587
rect 2915 3553 2924 3587
rect 2872 3544 2924 3553
rect 4160 3544 4212 3596
rect 6184 3587 6236 3596
rect 6184 3553 6193 3587
rect 6193 3553 6227 3587
rect 6227 3553 6236 3587
rect 6184 3544 6236 3553
rect 10784 3587 10836 3596
rect 10784 3553 10790 3587
rect 10790 3553 10836 3587
rect 10784 3544 10836 3553
rect 1952 3476 2004 3528
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 6920 3408 6972 3460
rect 9404 3476 9456 3528
rect 11336 3476 11388 3528
rect 9864 3408 9916 3460
rect 14280 3680 14332 3732
rect 16580 3680 16632 3732
rect 19984 3723 20036 3732
rect 19984 3689 19993 3723
rect 19993 3689 20027 3723
rect 20027 3689 20036 3723
rect 19984 3680 20036 3689
rect 20076 3680 20128 3732
rect 21180 3723 21232 3732
rect 21180 3689 21189 3723
rect 21189 3689 21223 3723
rect 21223 3689 21232 3723
rect 21180 3680 21232 3689
rect 22652 3723 22704 3732
rect 22652 3689 22661 3723
rect 22661 3689 22695 3723
rect 22695 3689 22704 3723
rect 22652 3680 22704 3689
rect 23480 3723 23532 3732
rect 23480 3689 23489 3723
rect 23489 3689 23523 3723
rect 23523 3689 23532 3723
rect 23480 3680 23532 3689
rect 24860 3723 24912 3732
rect 24860 3689 24869 3723
rect 24869 3689 24903 3723
rect 24903 3689 24912 3723
rect 24860 3680 24912 3689
rect 12164 3655 12216 3664
rect 12164 3621 12173 3655
rect 12173 3621 12207 3655
rect 12207 3621 12216 3655
rect 12164 3612 12216 3621
rect 13820 3655 13872 3664
rect 13820 3621 13829 3655
rect 13829 3621 13863 3655
rect 13863 3621 13872 3655
rect 13820 3612 13872 3621
rect 14372 3655 14424 3664
rect 14372 3621 14381 3655
rect 14381 3621 14415 3655
rect 14415 3621 14424 3655
rect 14372 3612 14424 3621
rect 15476 3655 15528 3664
rect 15476 3621 15485 3655
rect 15485 3621 15519 3655
rect 15519 3621 15528 3655
rect 15476 3612 15528 3621
rect 16212 3612 16264 3664
rect 16856 3655 16908 3664
rect 16856 3621 16865 3655
rect 16865 3621 16899 3655
rect 16899 3621 16908 3655
rect 16856 3612 16908 3621
rect 18420 3655 18472 3664
rect 18420 3621 18429 3655
rect 18429 3621 18463 3655
rect 18463 3621 18472 3655
rect 18420 3612 18472 3621
rect 18972 3655 19024 3664
rect 18972 3621 18981 3655
rect 18981 3621 19015 3655
rect 19015 3621 19024 3655
rect 21456 3655 21508 3664
rect 18972 3612 19024 3621
rect 21456 3621 21465 3655
rect 21465 3621 21499 3655
rect 21499 3621 21508 3655
rect 21456 3612 21508 3621
rect 21732 3612 21784 3664
rect 22192 3612 22244 3664
rect 12256 3544 12308 3596
rect 16948 3544 17000 3596
rect 20168 3544 20220 3596
rect 20812 3544 20864 3596
rect 22744 3544 22796 3596
rect 24952 3612 25004 3664
rect 25044 3587 25096 3596
rect 25044 3553 25053 3587
rect 25053 3553 25087 3587
rect 25087 3553 25096 3587
rect 25044 3544 25096 3553
rect 25320 3544 25372 3596
rect 14188 3476 14240 3528
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 18788 3476 18840 3528
rect 21916 3476 21968 3528
rect 23020 3476 23072 3528
rect 1768 3340 1820 3392
rect 1952 3383 2004 3392
rect 1952 3349 1961 3383
rect 1961 3349 1995 3383
rect 1995 3349 2004 3383
rect 1952 3340 2004 3349
rect 7012 3383 7064 3392
rect 7012 3349 7021 3383
rect 7021 3349 7055 3383
rect 7055 3349 7064 3383
rect 7012 3340 7064 3349
rect 9036 3383 9088 3392
rect 9036 3349 9045 3383
rect 9045 3349 9079 3383
rect 9079 3349 9088 3383
rect 9036 3340 9088 3349
rect 10508 3340 10560 3392
rect 10968 3340 11020 3392
rect 11244 3383 11296 3392
rect 11244 3349 11253 3383
rect 11253 3349 11287 3383
rect 11287 3349 11296 3383
rect 11244 3340 11296 3349
rect 12808 3340 12860 3392
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 17316 3340 17368 3349
rect 18144 3383 18196 3392
rect 18144 3349 18153 3383
rect 18153 3349 18187 3383
rect 18187 3349 18196 3383
rect 18144 3340 18196 3349
rect 24216 3383 24268 3392
rect 24216 3349 24225 3383
rect 24225 3349 24259 3383
rect 24259 3349 24268 3383
rect 24216 3340 24268 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1492 3136 1544 3188
rect 2872 3179 2924 3188
rect 2872 3145 2881 3179
rect 2881 3145 2915 3179
rect 2915 3145 2924 3179
rect 6184 3179 6236 3188
rect 2872 3136 2924 3145
rect 6184 3145 6193 3179
rect 6193 3145 6227 3179
rect 6227 3145 6236 3179
rect 6184 3136 6236 3145
rect 5540 3111 5592 3120
rect 5540 3077 5549 3111
rect 5549 3077 5583 3111
rect 5583 3077 5592 3111
rect 5540 3068 5592 3077
rect 2596 3000 2648 3052
rect 3240 3000 3292 3052
rect 4804 3000 4856 3052
rect 6828 3136 6880 3188
rect 7380 3136 7432 3188
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 9956 3136 10008 3188
rect 8576 3043 8628 3052
rect 1952 2975 2004 2984
rect 1952 2941 1961 2975
rect 1961 2941 1995 2975
rect 1995 2941 2004 2975
rect 1952 2932 2004 2941
rect 2320 2932 2372 2984
rect 3424 2975 3476 2984
rect 3424 2941 3433 2975
rect 3433 2941 3467 2975
rect 3467 2941 3476 2975
rect 3424 2932 3476 2941
rect 3792 2975 3844 2984
rect 3792 2941 3801 2975
rect 3801 2941 3835 2975
rect 3835 2941 3844 2975
rect 3792 2932 3844 2941
rect 2504 2907 2556 2916
rect 2504 2873 2513 2907
rect 2513 2873 2547 2907
rect 2547 2873 2556 2907
rect 2504 2864 2556 2873
rect 3976 2864 4028 2916
rect 4988 2907 5040 2916
rect 4988 2873 4997 2907
rect 4997 2873 5031 2907
rect 5031 2873 5040 2907
rect 4988 2864 5040 2873
rect 5080 2907 5132 2916
rect 5080 2873 5089 2907
rect 5089 2873 5123 2907
rect 5123 2873 5132 2907
rect 8576 3009 8585 3043
rect 8585 3009 8619 3043
rect 8619 3009 8628 3043
rect 8576 3000 8628 3009
rect 7012 2932 7064 2984
rect 9312 3000 9364 3052
rect 10784 3136 10836 3188
rect 10968 3136 11020 3188
rect 12164 3179 12216 3188
rect 12164 3145 12173 3179
rect 12173 3145 12207 3179
rect 12207 3145 12216 3179
rect 12164 3136 12216 3145
rect 13820 3136 13872 3188
rect 15476 3179 15528 3188
rect 15476 3145 15485 3179
rect 15485 3145 15519 3179
rect 15519 3145 15528 3179
rect 15476 3136 15528 3145
rect 16948 3136 17000 3188
rect 20168 3136 20220 3188
rect 22376 3136 22428 3188
rect 10508 3111 10560 3120
rect 10508 3077 10517 3111
rect 10517 3077 10551 3111
rect 10551 3077 10560 3111
rect 10508 3068 10560 3077
rect 10692 3111 10744 3120
rect 10692 3077 10701 3111
rect 10701 3077 10735 3111
rect 10735 3077 10744 3111
rect 10692 3068 10744 3077
rect 12440 3000 12492 3052
rect 12808 3043 12860 3052
rect 12808 3009 12817 3043
rect 12817 3009 12851 3043
rect 12851 3009 12860 3043
rect 12808 3000 12860 3009
rect 16856 3000 16908 3052
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 18788 3043 18840 3052
rect 18788 3009 18797 3043
rect 18797 3009 18831 3043
rect 18831 3009 18840 3043
rect 18788 3000 18840 3009
rect 18972 3000 19024 3052
rect 20812 3043 20864 3052
rect 20812 3009 20821 3043
rect 20821 3009 20855 3043
rect 20855 3009 20864 3043
rect 20812 3000 20864 3009
rect 22744 3000 22796 3052
rect 5080 2864 5132 2873
rect 9220 2975 9272 2984
rect 9220 2941 9229 2975
rect 9229 2941 9263 2975
rect 9263 2941 9272 2975
rect 9220 2932 9272 2941
rect 9864 2932 9916 2984
rect 11336 2932 11388 2984
rect 12900 2932 12952 2984
rect 14556 2975 14608 2984
rect 14556 2941 14565 2975
rect 14565 2941 14599 2975
rect 14599 2941 14608 2975
rect 14556 2932 14608 2941
rect 23204 3136 23256 3188
rect 23572 3136 23624 3188
rect 23756 3136 23808 3188
rect 25044 3179 25096 3188
rect 25044 3145 25053 3179
rect 25053 3145 25087 3179
rect 25087 3145 25096 3179
rect 25044 3136 25096 3145
rect 25320 3136 25372 3188
rect 23388 3068 23440 3120
rect 24032 3043 24084 3052
rect 24032 3009 24041 3043
rect 24041 3009 24075 3043
rect 24075 3009 24084 3043
rect 24032 3000 24084 3009
rect 24216 3000 24268 3052
rect 23572 2932 23624 2984
rect 25228 2975 25280 2984
rect 25228 2941 25237 2975
rect 25237 2941 25271 2975
rect 25271 2941 25280 2975
rect 25228 2932 25280 2941
rect 15660 2864 15712 2916
rect 16212 2864 16264 2916
rect 12624 2839 12676 2848
rect 12624 2805 12633 2839
rect 12633 2805 12667 2839
rect 12667 2805 12676 2839
rect 12624 2796 12676 2805
rect 18420 2864 18472 2916
rect 17408 2796 17460 2848
rect 19248 2864 19300 2916
rect 21088 2864 21140 2916
rect 21732 2839 21784 2848
rect 21732 2805 21741 2839
rect 21741 2805 21775 2839
rect 21775 2805 21784 2839
rect 21732 2796 21784 2805
rect 23572 2796 23624 2848
rect 23848 2796 23900 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 4804 2592 4856 2644
rect 4528 2567 4580 2576
rect 1492 2499 1544 2508
rect 1492 2465 1510 2499
rect 1510 2465 1544 2499
rect 4528 2533 4537 2567
rect 4537 2533 4571 2567
rect 4571 2533 4580 2567
rect 4528 2524 4580 2533
rect 6092 2592 6144 2644
rect 7840 2592 7892 2644
rect 8668 2592 8720 2644
rect 9588 2592 9640 2644
rect 7656 2567 7708 2576
rect 7656 2533 7665 2567
rect 7665 2533 7699 2567
rect 7699 2533 7708 2567
rect 7656 2524 7708 2533
rect 8300 2567 8352 2576
rect 8300 2533 8309 2567
rect 8309 2533 8343 2567
rect 8343 2533 8352 2567
rect 8300 2524 8352 2533
rect 1492 2456 1544 2465
rect 3424 2499 3476 2508
rect 3424 2465 3433 2499
rect 3433 2465 3467 2499
rect 3467 2465 3476 2499
rect 3424 2456 3476 2465
rect 5172 2456 5224 2508
rect 11152 2592 11204 2644
rect 12532 2592 12584 2644
rect 13636 2635 13688 2644
rect 13636 2601 13645 2635
rect 13645 2601 13679 2635
rect 13679 2601 13688 2635
rect 13636 2592 13688 2601
rect 14556 2635 14608 2644
rect 14556 2601 14565 2635
rect 14565 2601 14599 2635
rect 14599 2601 14608 2635
rect 14556 2592 14608 2601
rect 15660 2635 15712 2644
rect 15660 2601 15669 2635
rect 15669 2601 15703 2635
rect 15703 2601 15712 2635
rect 15660 2592 15712 2601
rect 16212 2592 16264 2644
rect 17408 2635 17460 2644
rect 12348 2524 12400 2576
rect 12624 2524 12676 2576
rect 17408 2601 17417 2635
rect 17417 2601 17451 2635
rect 17451 2601 17460 2635
rect 17408 2592 17460 2601
rect 18420 2592 18472 2644
rect 20628 2592 20680 2644
rect 21916 2592 21968 2644
rect 17868 2524 17920 2576
rect 21732 2524 21784 2576
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 11152 2499 11204 2508
rect 11152 2465 11161 2499
rect 11161 2465 11195 2499
rect 11195 2465 11204 2499
rect 11152 2456 11204 2465
rect 11428 2499 11480 2508
rect 11428 2465 11437 2499
rect 11437 2465 11471 2499
rect 11471 2465 11480 2499
rect 11428 2456 11480 2465
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 19984 2456 20036 2508
rect 3884 2388 3936 2440
rect 3976 2388 4028 2440
rect 7840 2388 7892 2440
rect 9496 2431 9548 2440
rect 9496 2397 9505 2431
rect 9505 2397 9539 2431
rect 9539 2397 9548 2431
rect 9496 2388 9548 2397
rect 10784 2388 10836 2440
rect 12716 2431 12768 2440
rect 12716 2397 12725 2431
rect 12725 2397 12759 2431
rect 12759 2397 12768 2431
rect 12716 2388 12768 2397
rect 16488 2431 16540 2440
rect 16488 2397 16497 2431
rect 16497 2397 16531 2431
rect 16531 2397 16540 2431
rect 16488 2388 16540 2397
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 21456 2388 21508 2440
rect 23112 2592 23164 2644
rect 23388 2592 23440 2644
rect 24124 2635 24176 2644
rect 24124 2601 24133 2635
rect 24133 2601 24167 2635
rect 24167 2601 24176 2635
rect 24124 2592 24176 2601
rect 25320 2592 25372 2644
rect 23664 2524 23716 2576
rect 26148 2456 26200 2508
rect 22744 2320 22796 2372
rect 2136 2252 2188 2304
rect 5448 2252 5500 2304
rect 8852 2295 8904 2304
rect 8852 2261 8861 2295
rect 8861 2261 8895 2295
rect 8895 2261 8904 2295
rect 8852 2252 8904 2261
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 10048 2252 10100 2304
rect 12624 2252 12676 2304
rect 21640 2252 21692 2304
rect 25136 2252 25188 2304
rect 26148 2295 26200 2304
rect 26148 2261 26157 2295
rect 26157 2261 26191 2295
rect 26191 2261 26200 2295
rect 26148 2252 26200 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 20260 2048 20312 2100
rect 22652 2048 22704 2100
rect 14464 1980 14516 2032
rect 14924 1980 14976 2032
rect 24584 1980 24636 2032
rect 25596 1980 25648 2032
rect 16856 552 16908 604
rect 18052 552 18104 604
<< metal2 >>
rect 662 27520 718 28000
rect 2042 27520 2098 28000
rect 3422 27520 3478 28000
rect 4802 27520 4858 28000
rect 6182 27520 6238 28000
rect 7654 27520 7710 28000
rect 9034 27520 9090 28000
rect 10414 27520 10470 28000
rect 11794 27520 11850 28000
rect 13174 27520 13230 28000
rect 14646 27520 14702 28000
rect 16026 27520 16082 28000
rect 17406 27520 17462 28000
rect 18786 27520 18842 28000
rect 20166 27520 20222 28000
rect 21638 27520 21694 28000
rect 23018 27520 23074 28000
rect 24398 27520 24454 28000
rect 25778 27520 25834 28000
rect 27158 27520 27214 28000
rect 676 23633 704 27520
rect 1398 27296 1454 27305
rect 1398 27231 1454 27240
rect 662 23624 718 23633
rect 662 23559 718 23568
rect 1412 23322 1440 27231
rect 1582 25936 1638 25945
rect 1582 25871 1638 25880
rect 1490 24576 1546 24585
rect 1490 24511 1546 24520
rect 1400 23316 1452 23322
rect 1400 23258 1452 23264
rect 1504 22778 1532 24511
rect 1596 23866 1624 25871
rect 2056 24290 2084 27520
rect 2056 24262 2176 24290
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 2044 23520 2096 23526
rect 2042 23488 2044 23497
rect 2096 23488 2098 23497
rect 2042 23423 2098 23432
rect 1676 23180 1728 23186
rect 1676 23122 1728 23128
rect 1582 23080 1638 23089
rect 1582 23015 1638 23024
rect 1492 22772 1544 22778
rect 1492 22714 1544 22720
rect 1596 21690 1624 23015
rect 1688 22030 1716 23122
rect 2148 22273 2176 24262
rect 2686 22672 2742 22681
rect 2686 22607 2742 22616
rect 2228 22432 2280 22438
rect 2228 22374 2280 22380
rect 2134 22264 2190 22273
rect 2134 22199 2190 22208
rect 1676 22024 1728 22030
rect 1674 21992 1676 22001
rect 1728 21992 1730 22001
rect 1674 21927 1730 21936
rect 1674 21720 1730 21729
rect 1584 21684 1636 21690
rect 1674 21655 1730 21664
rect 1584 21626 1636 21632
rect 1582 20360 1638 20369
rect 1582 20295 1638 20304
rect 1398 19680 1454 19689
rect 1398 19615 1454 19624
rect 1412 17626 1440 19615
rect 1596 19174 1624 20295
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1582 18864 1638 18873
rect 1582 18799 1638 18808
rect 1320 17598 1440 17626
rect 1320 16130 1348 17598
rect 1492 17536 1544 17542
rect 1398 17504 1454 17513
rect 1492 17478 1544 17484
rect 1398 17439 1454 17448
rect 1412 16250 1440 17439
rect 1400 16244 1452 16250
rect 1400 16186 1452 16192
rect 1320 16102 1440 16130
rect 1308 15360 1360 15366
rect 1308 15302 1360 15308
rect 1320 11762 1348 15302
rect 1308 11756 1360 11762
rect 1308 11698 1360 11704
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 1320 9518 1348 9998
rect 1308 9512 1360 9518
rect 1308 9454 1360 9460
rect 1214 9072 1270 9081
rect 1214 9007 1270 9016
rect 1122 7848 1178 7857
rect 1122 7783 1178 7792
rect 1136 5778 1164 7783
rect 1228 7002 1256 9007
rect 1308 8560 1360 8566
rect 1308 8502 1360 8508
rect 1216 6996 1268 7002
rect 1216 6938 1268 6944
rect 1124 5772 1176 5778
rect 1124 5714 1176 5720
rect 1136 4758 1164 5714
rect 1124 4752 1176 4758
rect 1124 4694 1176 4700
rect 478 2408 534 2417
rect 478 2343 534 2352
rect 492 480 520 2343
rect 1320 2145 1348 8502
rect 1306 2136 1362 2145
rect 1306 2071 1362 2080
rect 1412 480 1440 16102
rect 1504 14074 1532 17478
rect 1596 17338 1624 18799
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 1596 16289 1624 17138
rect 1582 16280 1638 16289
rect 1582 16215 1638 16224
rect 1582 16144 1638 16153
rect 1582 16079 1638 16088
rect 1596 14618 1624 16079
rect 1688 15706 1716 21655
rect 2044 21480 2096 21486
rect 2044 21422 2096 21428
rect 1952 20256 2004 20262
rect 1952 20198 2004 20204
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1872 18630 1900 19858
rect 1860 18624 1912 18630
rect 1860 18566 1912 18572
rect 1768 18080 1820 18086
rect 1768 18022 1820 18028
rect 1780 16561 1808 18022
rect 1766 16552 1822 16561
rect 1766 16487 1822 16496
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1676 15428 1728 15434
rect 1676 15370 1728 15376
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1492 14068 1544 14074
rect 1492 14010 1544 14016
rect 1596 13172 1624 14418
rect 1688 13274 1716 15370
rect 1780 13433 1808 16390
rect 1872 14793 1900 18566
rect 1964 16454 1992 20198
rect 2056 17202 2084 21422
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2148 18873 2176 19110
rect 2134 18864 2190 18873
rect 2240 18834 2268 22374
rect 2412 20528 2464 20534
rect 2412 20470 2464 20476
rect 2320 19372 2372 19378
rect 2320 19314 2372 19320
rect 2134 18799 2190 18808
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2228 18692 2280 18698
rect 2228 18634 2280 18640
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2148 16998 2176 17682
rect 2044 16992 2096 16998
rect 2042 16960 2044 16969
rect 2136 16992 2188 16998
rect 2096 16960 2098 16969
rect 2136 16934 2188 16940
rect 2042 16895 2098 16904
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 2056 16266 2084 16390
rect 1964 16238 2084 16266
rect 1964 15162 1992 16238
rect 2042 16144 2098 16153
rect 2042 16079 2044 16088
rect 2096 16079 2098 16088
rect 2044 16050 2096 16056
rect 2042 16008 2098 16017
rect 2042 15943 2098 15952
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 2056 14906 2084 15943
rect 2148 15366 2176 16594
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 1964 14878 2084 14906
rect 1858 14784 1914 14793
rect 1858 14719 1914 14728
rect 1964 14634 1992 14878
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 1872 14606 1992 14634
rect 1766 13424 1822 13433
rect 1766 13359 1822 13368
rect 1688 13246 1808 13274
rect 1676 13184 1728 13190
rect 1596 13144 1676 13172
rect 1676 13126 1728 13132
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1504 11898 1532 12242
rect 1492 11892 1544 11898
rect 1492 11834 1544 11840
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1504 9636 1532 11698
rect 1596 11354 1624 11698
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1582 11248 1638 11257
rect 1582 11183 1584 11192
rect 1636 11183 1638 11192
rect 1584 11154 1636 11160
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1596 10062 1624 11018
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1596 9761 1624 9862
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1504 9608 1624 9636
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 4078 1532 8298
rect 1596 7426 1624 9608
rect 1688 7546 1716 13126
rect 1780 12918 1808 13246
rect 1768 12912 1820 12918
rect 1768 12854 1820 12860
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1780 10810 1808 11154
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1768 10192 1820 10198
rect 1768 10134 1820 10140
rect 1780 9654 1808 10134
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 1780 8974 1808 9590
rect 1872 9489 1900 14606
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1964 10062 1992 12038
rect 2044 11824 2096 11830
rect 2044 11766 2096 11772
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1964 9586 1992 9862
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1858 9480 1914 9489
rect 1858 9415 1914 9424
rect 1952 9444 2004 9450
rect 1952 9386 2004 9392
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1780 7750 1808 8366
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1780 7449 1808 7686
rect 1766 7440 1822 7449
rect 1596 7398 1716 7426
rect 1582 5944 1638 5953
rect 1582 5879 1584 5888
rect 1636 5879 1638 5888
rect 1584 5850 1636 5856
rect 1688 5794 1716 7398
rect 1766 7375 1822 7384
rect 1872 6769 1900 7822
rect 1858 6760 1914 6769
rect 1858 6695 1914 6704
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1780 6361 1808 6598
rect 1766 6352 1822 6361
rect 1766 6287 1822 6296
rect 1596 5766 1716 5794
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1504 3777 1532 4014
rect 1490 3768 1546 3777
rect 1490 3703 1546 3712
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 1504 3505 1532 3538
rect 1490 3496 1546 3505
rect 1490 3431 1546 3440
rect 1504 3194 1532 3431
rect 1596 3233 1624 5766
rect 1872 4826 1900 6695
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1964 4282 1992 9386
rect 2056 5114 2084 11766
rect 2148 10713 2176 14758
rect 2134 10704 2190 10713
rect 2134 10639 2190 10648
rect 2240 9654 2268 18634
rect 2332 16182 2360 19314
rect 2320 16176 2372 16182
rect 2320 16118 2372 16124
rect 2424 15570 2452 20470
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 2502 18728 2558 18737
rect 2502 18663 2558 18672
rect 2516 18426 2544 18663
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2608 18170 2636 19654
rect 2700 18766 2728 22607
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 3068 19514 3096 19858
rect 3160 19825 3188 20198
rect 3146 19816 3202 19825
rect 3146 19751 3202 19760
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 2688 18760 2740 18766
rect 2688 18702 2740 18708
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2516 18142 2636 18170
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 2424 15162 2452 15506
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2332 12481 2360 14894
rect 2516 13326 2544 18142
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 2608 17241 2636 18022
rect 2594 17232 2650 17241
rect 2594 17167 2650 17176
rect 2596 16992 2648 16998
rect 2596 16934 2648 16940
rect 2608 16697 2636 16934
rect 2594 16688 2650 16697
rect 2594 16623 2650 16632
rect 2700 15473 2728 18566
rect 2778 17096 2834 17105
rect 2778 17031 2834 17040
rect 2792 16998 2820 17031
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2686 15464 2742 15473
rect 2686 15399 2742 15408
rect 2792 14226 2820 16594
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2884 15434 2912 15982
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2872 15428 2924 15434
rect 2872 15370 2924 15376
rect 2976 14890 3004 15506
rect 2964 14884 3016 14890
rect 2964 14826 3016 14832
rect 3068 14346 3096 19450
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3252 19009 3280 19110
rect 3238 19000 3294 19009
rect 3238 18935 3294 18944
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3160 18222 3188 18770
rect 3436 18714 3464 27520
rect 4816 24857 4844 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 4802 24848 4858 24857
rect 4802 24783 4858 24792
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5446 23896 5502 23905
rect 5622 23888 5918 23908
rect 5502 23854 5580 23882
rect 5446 23831 5502 23840
rect 5078 23760 5134 23769
rect 5078 23695 5134 23704
rect 5092 23497 5120 23695
rect 5078 23488 5134 23497
rect 5078 23423 5134 23432
rect 5262 23488 5318 23497
rect 5262 23423 5318 23432
rect 5172 22160 5224 22166
rect 5170 22128 5172 22137
rect 5224 22128 5226 22137
rect 5170 22063 5226 22072
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 3792 20392 3844 20398
rect 3792 20334 3844 20340
rect 3516 19712 3568 19718
rect 3804 19689 3832 20334
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3516 19654 3568 19660
rect 3790 19680 3846 19689
rect 3344 18686 3464 18714
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 3160 18086 3188 18158
rect 3148 18080 3200 18086
rect 3148 18022 3200 18028
rect 3160 16454 3188 18022
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3148 14952 3200 14958
rect 3146 14920 3148 14929
rect 3200 14920 3202 14929
rect 3146 14855 3202 14864
rect 3146 14784 3202 14793
rect 3146 14719 3202 14728
rect 3160 14618 3188 14719
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3146 14512 3202 14521
rect 3146 14447 3148 14456
rect 3200 14447 3202 14456
rect 3148 14418 3200 14424
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 2792 14198 3096 14226
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2688 14000 2740 14006
rect 2688 13942 2740 13948
rect 2700 13462 2728 13942
rect 2792 13462 2820 14010
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2780 13456 2832 13462
rect 2780 13398 2832 13404
rect 2870 13424 2926 13433
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2516 12986 2544 13262
rect 2700 12986 2728 13398
rect 2870 13359 2926 13368
rect 2884 13258 2912 13359
rect 2872 13252 2924 13258
rect 2872 13194 2924 13200
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2318 12472 2374 12481
rect 2318 12407 2374 12416
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2332 11558 2360 12242
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2320 11552 2372 11558
rect 2318 11520 2320 11529
rect 2372 11520 2374 11529
rect 2318 11455 2374 11464
rect 2424 11268 2452 12038
rect 2504 11280 2556 11286
rect 2424 11240 2504 11268
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2332 10742 2360 11086
rect 2320 10736 2372 10742
rect 2320 10678 2372 10684
rect 2424 10674 2452 11240
rect 2504 11222 2556 11228
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2608 10810 2636 11154
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2424 10130 2452 10610
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2332 9897 2360 10066
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2318 9888 2374 9897
rect 2318 9823 2374 9832
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2148 5302 2176 9522
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2240 5658 2268 9454
rect 2332 9110 2360 9823
rect 2424 9330 2452 9930
rect 2516 9722 2544 10542
rect 2596 10192 2648 10198
rect 2648 10140 2728 10146
rect 2596 10134 2728 10140
rect 2608 10118 2728 10134
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2424 9302 2544 9330
rect 2410 9208 2466 9217
rect 2410 9143 2466 9152
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 2332 7546 2360 7958
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2332 5778 2360 6598
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2240 5630 2360 5658
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2240 5370 2268 5510
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2136 5296 2188 5302
rect 2136 5238 2188 5244
rect 2332 5234 2360 5630
rect 2424 5370 2452 9143
rect 2516 7818 2544 9302
rect 2608 9058 2636 9998
rect 2700 9178 2728 10118
rect 2792 10033 2820 12582
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 2884 12209 2912 12242
rect 2870 12200 2926 12209
rect 2870 12135 2926 12144
rect 2884 11354 2912 12135
rect 2976 11898 3004 12242
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2870 11248 2926 11257
rect 2870 11183 2926 11192
rect 2884 11150 2912 11183
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2778 10024 2834 10033
rect 2778 9959 2834 9968
rect 2778 9752 2834 9761
rect 2778 9687 2834 9696
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2608 9030 2728 9058
rect 2700 8974 2728 9030
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 2516 7342 2544 7754
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2502 7168 2558 7177
rect 2502 7103 2558 7112
rect 2516 6254 2544 7103
rect 2504 6248 2556 6254
rect 2504 6190 2556 6196
rect 2516 5914 2544 6190
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2136 5160 2188 5166
rect 2056 5108 2136 5114
rect 2056 5102 2188 5108
rect 2056 5086 2176 5102
rect 2516 5098 2544 5714
rect 2504 5092 2556 5098
rect 2504 5034 2556 5040
rect 2410 4856 2466 4865
rect 2410 4791 2466 4800
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 1952 4276 2004 4282
rect 1952 4218 2004 4224
rect 1964 3534 1992 4218
rect 2240 3738 2268 4626
rect 2424 4185 2452 4791
rect 2516 4690 2544 5034
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 2608 4486 2636 8910
rect 2700 8090 2728 8910
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 2700 6322 2728 6734
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2700 5710 2728 6258
rect 2688 5704 2740 5710
rect 2792 5681 2820 9687
rect 2884 9450 2912 10746
rect 2976 9654 3004 11834
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2884 9042 2912 9386
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2884 8786 2912 8978
rect 2976 8906 3004 9590
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 2884 8758 3004 8786
rect 2976 8498 3004 8758
rect 3068 8566 3096 14198
rect 3160 13938 3188 14418
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3146 12472 3202 12481
rect 3146 12407 3202 12416
rect 3160 9654 3188 12407
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2976 7426 3004 8434
rect 3160 8430 3188 9318
rect 3148 8424 3200 8430
rect 3146 8392 3148 8401
rect 3200 8392 3202 8401
rect 3146 8327 3202 8336
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3160 7868 3188 8230
rect 3252 7993 3280 17614
rect 3344 16522 3372 18686
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3332 16516 3384 16522
rect 3332 16458 3384 16464
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 3344 15609 3372 15914
rect 3330 15600 3386 15609
rect 3330 15535 3386 15544
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3344 13870 3372 14554
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3344 13530 3372 13806
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3332 12368 3384 12374
rect 3330 12336 3332 12345
rect 3384 12336 3386 12345
rect 3330 12271 3386 12280
rect 3330 9344 3386 9353
rect 3330 9279 3386 9288
rect 3238 7984 3294 7993
rect 3238 7919 3294 7928
rect 3160 7840 3280 7868
rect 2976 7398 3096 7426
rect 2962 6896 3018 6905
rect 2872 6860 2924 6866
rect 2962 6831 3018 6840
rect 2872 6802 2924 6808
rect 2884 6458 2912 6802
rect 2976 6798 3004 6831
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2976 6458 3004 6598
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2688 5646 2740 5652
rect 2778 5672 2834 5681
rect 2884 5642 2912 6394
rect 2778 5607 2834 5616
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2700 5386 2728 5510
rect 2700 5358 2820 5386
rect 2792 5302 2820 5358
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2686 5128 2742 5137
rect 2686 5063 2742 5072
rect 2700 4554 2728 5063
rect 2792 5001 2820 5238
rect 2884 5216 2912 5578
rect 2976 5409 3004 6394
rect 2962 5400 3018 5409
rect 2962 5335 3018 5344
rect 2964 5228 3016 5234
rect 2884 5188 2964 5216
rect 2964 5170 3016 5176
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2778 4992 2834 5001
rect 2778 4927 2834 4936
rect 2792 4826 2820 4927
rect 2884 4865 2912 5034
rect 2870 4856 2926 4865
rect 2780 4820 2832 4826
rect 2976 4826 3004 5170
rect 2870 4791 2926 4800
rect 2964 4820 3016 4826
rect 2780 4762 2832 4768
rect 2884 4622 2912 4791
rect 2964 4762 3016 4768
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2700 4434 2728 4490
rect 2410 4176 2466 4185
rect 2410 4111 2466 4120
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1582 3224 1638 3233
rect 1492 3188 1544 3194
rect 1582 3159 1638 3168
rect 1492 3130 1544 3136
rect 1504 2961 1532 3130
rect 1780 3097 1808 3334
rect 1766 3088 1822 3097
rect 1766 3023 1822 3032
rect 1964 2990 1992 3334
rect 2608 3058 2636 4422
rect 2700 4406 2820 4434
rect 2688 4072 2740 4078
rect 2686 4040 2688 4049
rect 2740 4040 2742 4049
rect 2686 3975 2742 3984
rect 2792 3738 2820 4406
rect 2884 4282 2912 4558
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 3068 3754 3096 7398
rect 3146 7304 3202 7313
rect 3252 7274 3280 7840
rect 3146 7239 3202 7248
rect 3240 7268 3292 7274
rect 3160 4078 3188 7239
rect 3240 7210 3292 7216
rect 3344 5896 3372 9279
rect 3436 7834 3464 18566
rect 3528 8022 3556 19654
rect 3790 19615 3846 19624
rect 3896 19417 3924 20198
rect 4172 19922 4200 20742
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 3882 19408 3938 19417
rect 3882 19343 3938 19352
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3882 19272 3938 19281
rect 3620 16046 3648 19246
rect 3882 19207 3938 19216
rect 3896 19174 3924 19207
rect 3884 19168 3936 19174
rect 3884 19110 3936 19116
rect 4066 19136 4122 19145
rect 4066 19071 4122 19080
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3700 16652 3752 16658
rect 3700 16594 3752 16600
rect 3608 16040 3660 16046
rect 3712 16017 3740 16594
rect 3608 15982 3660 15988
rect 3698 16008 3754 16017
rect 3620 15745 3648 15982
rect 3698 15943 3700 15952
rect 3752 15943 3754 15952
rect 3700 15914 3752 15920
rect 3606 15736 3662 15745
rect 3606 15671 3662 15680
rect 3620 15502 3648 15671
rect 3608 15496 3660 15502
rect 3608 15438 3660 15444
rect 3700 15428 3752 15434
rect 3700 15370 3752 15376
rect 3608 15360 3660 15366
rect 3608 15302 3660 15308
rect 3620 14482 3648 15302
rect 3712 14958 3740 15370
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3712 14550 3740 14894
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3608 14476 3660 14482
rect 3608 14418 3660 14424
rect 3620 11898 3648 14418
rect 3700 14340 3752 14346
rect 3700 14282 3752 14288
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3712 11150 3740 14282
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3712 9926 3740 10950
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3620 8838 3648 9454
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3712 8090 3740 9862
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3516 8016 3568 8022
rect 3516 7958 3568 7964
rect 3436 7806 3740 7834
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3620 7342 3648 7686
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3620 6322 3648 7278
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3252 5868 3372 5896
rect 3252 4758 3280 5868
rect 3712 5681 3740 7806
rect 3804 5846 3832 17138
rect 3896 12714 3924 18702
rect 4080 18086 4108 19071
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 4172 18222 4200 18906
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 4172 17898 4200 18158
rect 4080 17882 4200 17898
rect 4068 17876 4200 17882
rect 4120 17870 4200 17876
rect 4068 17818 4120 17824
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3988 16697 4016 16934
rect 4066 16824 4122 16833
rect 4066 16759 4068 16768
rect 4120 16759 4122 16768
rect 4068 16730 4120 16736
rect 4252 16720 4304 16726
rect 3974 16688 4030 16697
rect 4252 16662 4304 16668
rect 3974 16623 4030 16632
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 4080 14929 4108 16458
rect 4264 15978 4292 16662
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 4264 15706 4292 15914
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4356 15366 4384 16526
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4356 15026 4384 15302
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4160 14952 4212 14958
rect 4066 14920 4122 14929
rect 4160 14894 4212 14900
rect 4066 14855 4122 14864
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3988 13462 4016 13738
rect 4080 13530 4108 14486
rect 4172 14482 4200 14894
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4172 14074 4200 14418
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 4080 13410 4108 13466
rect 4080 13382 4292 13410
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3988 12714 4016 13126
rect 4080 12986 4108 13262
rect 4068 12980 4120 12986
rect 4120 12940 4200 12968
rect 4068 12922 4120 12928
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 3988 12442 4016 12650
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4080 12322 4108 12786
rect 4172 12442 4200 12940
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 3884 12300 3936 12306
rect 4080 12294 4200 12322
rect 4264 12306 4292 13382
rect 4356 12442 4384 14758
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 3884 12242 3936 12248
rect 3896 11898 3924 12242
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3896 9110 3924 10066
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3896 8537 3924 8774
rect 3882 8528 3938 8537
rect 3882 8463 3938 8472
rect 3896 7546 3924 8463
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3896 6746 3924 7482
rect 3988 6866 4016 11494
rect 4080 11286 4108 11630
rect 4172 11354 4200 12294
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4264 11286 4292 12242
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3896 6718 4016 6746
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3422 5672 3478 5681
rect 3422 5607 3478 5616
rect 3698 5672 3754 5681
rect 3698 5607 3754 5616
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3344 4690 3372 5510
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3344 4486 3372 4626
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3344 4282 3372 4422
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2780 3732 2832 3738
rect 3068 3726 3372 3754
rect 2780 3674 2832 3680
rect 2700 3482 2728 3674
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2700 3454 2820 3482
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 1952 2984 2004 2990
rect 1490 2952 1546 2961
rect 1952 2926 2004 2932
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 1490 2887 1546 2896
rect 1492 2508 1544 2514
rect 1492 2450 1544 2456
rect 1504 2417 1532 2450
rect 1490 2408 1546 2417
rect 1490 2343 1546 2352
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2148 1873 2176 2246
rect 2134 1864 2190 1873
rect 2134 1799 2190 1808
rect 2332 480 2360 2926
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 2516 2825 2544 2858
rect 2502 2816 2558 2825
rect 2502 2751 2558 2760
rect 2792 785 2820 3454
rect 2884 3194 2912 3538
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3252 1465 3280 2994
rect 3238 1456 3294 1465
rect 3238 1391 3294 1400
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 3344 480 3372 3726
rect 3436 2990 3464 5607
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3698 5128 3754 5137
rect 3698 5063 3754 5072
rect 3712 4593 3740 5063
rect 3698 4584 3754 4593
rect 3698 4519 3754 4528
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3712 3738 3740 4014
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3804 3641 3832 5510
rect 3896 5273 3924 6598
rect 3988 6254 4016 6718
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 4080 5794 4108 11086
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4264 9926 4292 10406
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4356 9382 4384 9658
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4356 9042 4384 9318
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4356 8294 4384 8978
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4264 8022 4292 8230
rect 4252 8016 4304 8022
rect 4158 7984 4214 7993
rect 4252 7958 4304 7964
rect 4158 7919 4214 7928
rect 4172 7886 4200 7919
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4172 7546 4200 7822
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4264 7002 4292 7958
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4080 5766 4200 5794
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3882 5264 3938 5273
rect 3882 5199 3938 5208
rect 3882 5128 3938 5137
rect 3882 5063 3884 5072
rect 3936 5063 3938 5072
rect 3884 5034 3936 5040
rect 3896 4826 3924 5034
rect 3988 4842 4016 5646
rect 4080 5234 4108 5646
rect 4172 5574 4200 5766
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3988 4826 4200 4842
rect 3884 4820 3936 4826
rect 3988 4820 4212 4826
rect 3988 4814 4160 4820
rect 3884 4762 3936 4768
rect 4160 4762 4212 4768
rect 4172 4729 4200 4762
rect 4158 4720 4214 4729
rect 4158 4655 4214 4664
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 3790 3632 3846 3641
rect 4172 3602 4200 3946
rect 4264 3738 4292 4014
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4356 3618 4384 8230
rect 4448 4622 4476 21286
rect 5092 21010 5120 21286
rect 5276 21146 5304 23423
rect 5552 22574 5580 23854
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 6196 22216 6224 27520
rect 7668 24721 7696 27520
rect 9048 24834 9076 27520
rect 10428 25786 10456 27520
rect 10428 25758 10824 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 9048 24806 9260 24834
rect 7654 24712 7710 24721
rect 7654 24647 7710 24656
rect 8574 23760 8630 23769
rect 8574 23695 8630 23704
rect 8588 23186 8616 23695
rect 8944 23656 8996 23662
rect 8942 23624 8944 23633
rect 8996 23624 8998 23633
rect 8942 23559 8998 23568
rect 9128 23520 9180 23526
rect 9126 23488 9128 23497
rect 9180 23488 9182 23497
rect 9126 23423 9182 23432
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 8576 23180 8628 23186
rect 8576 23122 8628 23128
rect 6274 22808 6330 22817
rect 6274 22743 6276 22752
rect 6328 22743 6330 22752
rect 6276 22714 6328 22720
rect 6288 22574 6316 22714
rect 7300 22710 7328 23122
rect 7472 23112 7524 23118
rect 7472 23054 7524 23060
rect 7288 22704 7340 22710
rect 7288 22646 7340 22652
rect 7484 22642 7512 23054
rect 7656 22976 7708 22982
rect 7656 22918 7708 22924
rect 8298 22944 8354 22953
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 6276 22568 6328 22574
rect 6276 22510 6328 22516
rect 6736 22500 6788 22506
rect 6736 22442 6788 22448
rect 6196 22188 6408 22216
rect 6184 22092 6236 22098
rect 6184 22034 6236 22040
rect 5540 22024 5592 22030
rect 5538 21992 5540 22001
rect 5592 21992 5594 22001
rect 5538 21927 5594 21936
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6196 21690 6224 22034
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6274 21448 6330 21457
rect 6274 21383 6276 21392
rect 6328 21383 6330 21392
rect 6276 21354 6328 21360
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 5264 21140 5316 21146
rect 5264 21082 5316 21088
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 5080 21004 5132 21010
rect 5080 20946 5132 20952
rect 4724 20262 4752 20946
rect 5276 20398 5304 21082
rect 5632 20936 5684 20942
rect 5552 20884 5632 20890
rect 5552 20878 5684 20884
rect 5552 20862 5672 20878
rect 4896 20392 4948 20398
rect 5264 20392 5316 20398
rect 4896 20334 4948 20340
rect 5078 20360 5134 20369
rect 4712 20256 4764 20262
rect 4712 20198 4764 20204
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 4632 15162 4660 19450
rect 4908 18698 4936 20334
rect 5264 20334 5316 20340
rect 5078 20295 5134 20304
rect 5092 19922 5120 20295
rect 5276 19922 5304 20334
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 5092 19514 5120 19858
rect 5080 19508 5132 19514
rect 5080 19450 5132 19456
rect 5276 19310 5304 19858
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 4896 18692 4948 18698
rect 4896 18634 4948 18640
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4724 17746 4752 18158
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4724 17338 4752 17682
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4710 17232 4766 17241
rect 4710 17167 4712 17176
rect 4764 17167 4766 17176
rect 4712 17138 4764 17144
rect 4724 16726 4752 17138
rect 4816 17066 4844 17478
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4816 16250 4844 17002
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4908 15638 4936 18634
rect 5184 18612 5212 19246
rect 5276 18970 5304 19246
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5264 18624 5316 18630
rect 5184 18584 5264 18612
rect 5264 18566 5316 18572
rect 5276 18290 5304 18566
rect 5354 18320 5410 18329
rect 5264 18284 5316 18290
rect 5354 18255 5410 18264
rect 5264 18226 5316 18232
rect 5368 18222 5396 18255
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5276 17338 5304 17682
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4618 13288 4674 13297
rect 4618 13223 4620 13232
rect 4672 13223 4674 13232
rect 4620 13194 4672 13200
rect 4632 12850 4660 13194
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4724 12170 4752 13806
rect 4896 13456 4948 13462
rect 5000 13433 5028 16934
rect 5092 15094 5120 17274
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5368 16658 5396 17002
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5356 15904 5408 15910
rect 5262 15872 5318 15881
rect 5356 15846 5408 15852
rect 5262 15807 5318 15816
rect 5276 15706 5304 15807
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 5080 15088 5132 15094
rect 5080 15030 5132 15036
rect 5092 14958 5120 15030
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5092 14618 5120 14894
rect 5184 14822 5212 15506
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 5184 13977 5212 14758
rect 5276 14618 5304 15506
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5170 13968 5226 13977
rect 5170 13903 5226 13912
rect 5184 13870 5212 13903
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 4896 13398 4948 13404
rect 4986 13424 5042 13433
rect 4908 12646 4936 13398
rect 4986 13359 5042 13368
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4540 11082 4568 11698
rect 4632 11694 4660 12038
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4632 11218 4660 11630
rect 4724 11257 4752 12106
rect 4710 11248 4766 11257
rect 4620 11212 4672 11218
rect 4710 11183 4766 11192
rect 4620 11154 4672 11160
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4540 10606 4568 11018
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4632 10266 4660 11154
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4632 9722 4660 10066
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4632 9450 4660 9658
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4724 8634 4752 11183
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4816 10810 4844 11086
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4816 10130 4844 10746
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4908 9994 4936 10406
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4908 9518 4936 9930
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4816 9178 4844 9454
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4724 6866 4752 8026
rect 5000 7721 5028 13359
rect 5078 11656 5134 11665
rect 5078 11591 5080 11600
rect 5132 11591 5134 11600
rect 5080 11562 5132 11568
rect 5276 11218 5304 14554
rect 5368 13802 5396 15846
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5460 13682 5488 20198
rect 5552 19990 5580 20862
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5908 20324 5960 20330
rect 5908 20266 5960 20272
rect 5540 19984 5592 19990
rect 5920 19961 5948 20266
rect 5540 19926 5592 19932
rect 5906 19952 5962 19961
rect 5906 19887 5962 19896
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5816 19304 5868 19310
rect 5816 19246 5868 19252
rect 5828 18834 5856 19246
rect 5540 18828 5592 18834
rect 5540 18770 5592 18776
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 5552 17882 5580 18770
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5552 13938 5580 17274
rect 6012 16810 6040 21286
rect 6092 21004 6144 21010
rect 6092 20946 6144 20952
rect 6104 20534 6132 20946
rect 6380 20602 6408 22188
rect 6644 21072 6696 21078
rect 6644 21014 6696 21020
rect 6552 20800 6604 20806
rect 6552 20742 6604 20748
rect 6368 20596 6420 20602
rect 6368 20538 6420 20544
rect 6092 20528 6144 20534
rect 6092 20470 6144 20476
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 6104 18902 6132 20334
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 6196 19378 6224 19790
rect 6184 19372 6236 19378
rect 6380 19360 6408 20538
rect 6380 19332 6500 19360
rect 6184 19314 6236 19320
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 6092 18896 6144 18902
rect 6092 18838 6144 18844
rect 6090 17912 6146 17921
rect 6090 17847 6146 17856
rect 6104 16969 6132 17847
rect 6196 17814 6224 19110
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 6196 16998 6224 17750
rect 6184 16992 6236 16998
rect 6090 16960 6146 16969
rect 6184 16934 6236 16940
rect 6090 16895 6146 16904
rect 6012 16782 6132 16810
rect 6000 16720 6052 16726
rect 5906 16688 5962 16697
rect 6000 16662 6052 16668
rect 5906 16623 5962 16632
rect 5920 16590 5948 16623
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 16250 6040 16662
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5368 13654 5488 13682
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5262 10432 5318 10441
rect 5262 10367 5318 10376
rect 5276 10266 5304 10367
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5092 9518 5120 10066
rect 5262 9888 5318 9897
rect 5262 9823 5318 9832
rect 5276 9586 5304 9823
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5092 9042 5120 9454
rect 5264 9444 5316 9450
rect 5264 9386 5316 9392
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5276 8838 5304 9386
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 8090 5212 8230
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 4986 7712 5042 7721
rect 4986 7647 5042 7656
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4908 6934 4936 7346
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4540 6254 4568 6802
rect 4724 6458 4752 6802
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4528 6248 4580 6254
rect 4526 6216 4528 6225
rect 4580 6216 4582 6225
rect 4526 6151 4582 6160
rect 4528 5840 4580 5846
rect 4528 5782 4580 5788
rect 4540 5370 4568 5782
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4724 5166 4752 6394
rect 4894 6352 4950 6361
rect 4894 6287 4896 6296
rect 4948 6287 4950 6296
rect 4896 6258 4948 6264
rect 5184 6186 5212 6598
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 4802 5944 4858 5953
rect 5184 5914 5212 6122
rect 4802 5879 4858 5888
rect 5172 5908 5224 5914
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4724 4826 4752 5102
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4724 4078 4752 4762
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4816 4010 4844 5879
rect 5172 5850 5224 5856
rect 4894 5672 4950 5681
rect 4894 5607 4950 5616
rect 4908 5234 4936 5607
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 5184 5098 5212 5850
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 5092 4146 5120 4694
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4448 3777 4476 3878
rect 4434 3768 4490 3777
rect 5092 3738 5120 4082
rect 4434 3703 4490 3712
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 3790 3567 3846 3576
rect 4160 3596 4212 3602
rect 3804 2990 3832 3567
rect 4160 3538 4212 3544
rect 4264 3590 4384 3618
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 3436 2514 3464 2926
rect 3804 2650 3832 2926
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3988 2446 4016 2858
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 3896 1601 3924 2382
rect 3882 1592 3938 1601
rect 3882 1527 3938 1536
rect 4264 480 4292 3590
rect 4816 3058 4844 3606
rect 4986 3088 5042 3097
rect 4804 3052 4856 3058
rect 4986 3023 5042 3032
rect 4804 2994 4856 3000
rect 4816 2650 4844 2994
rect 5000 2922 5028 3023
rect 5092 2922 5120 3674
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4528 2576 4580 2582
rect 5000 2553 5028 2858
rect 5170 2680 5226 2689
rect 5170 2615 5226 2624
rect 4528 2518 4580 2524
rect 4986 2544 5042 2553
rect 4540 2417 4568 2518
rect 5184 2514 5212 2615
rect 4986 2479 5042 2488
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 4526 2408 4582 2417
rect 4526 2343 4582 2352
rect 5276 480 5304 8774
rect 5368 4282 5396 13654
rect 5552 11150 5580 13670
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5552 10810 5580 11086
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 6012 10305 6040 12650
rect 6104 12481 6132 16782
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6196 16250 6224 16526
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 6288 16130 6316 18158
rect 6380 18086 6408 18702
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6380 17513 6408 18022
rect 6366 17504 6422 17513
rect 6366 17439 6422 17448
rect 6380 17338 6408 17439
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6196 16102 6316 16130
rect 6196 14414 6224 16102
rect 6380 15978 6408 16934
rect 6368 15972 6420 15978
rect 6368 15914 6420 15920
rect 6380 15638 6408 15914
rect 6368 15632 6420 15638
rect 6368 15574 6420 15580
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6380 15026 6408 15302
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6196 14113 6224 14350
rect 6182 14104 6238 14113
rect 6288 14074 6316 14418
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6182 14039 6184 14048
rect 6236 14039 6238 14048
rect 6276 14068 6328 14074
rect 6184 14010 6236 14016
rect 6276 14010 6328 14016
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6090 12472 6146 12481
rect 6090 12407 6146 12416
rect 6288 12374 6316 13874
rect 6380 13530 6408 14350
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6472 12594 6500 19332
rect 6564 15722 6592 20742
rect 6656 20262 6684 21014
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6656 19990 6684 20198
rect 6644 19984 6696 19990
rect 6644 19926 6696 19932
rect 6656 19174 6684 19926
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6656 17202 6684 18090
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6656 16250 6684 17138
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6564 15694 6684 15722
rect 6550 15600 6606 15609
rect 6550 15535 6552 15544
rect 6604 15535 6606 15544
rect 6552 15506 6604 15512
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6564 13462 6592 14758
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6564 12714 6592 13398
rect 6656 13025 6684 15694
rect 6642 13016 6698 13025
rect 6642 12951 6698 12960
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 6472 12566 6592 12594
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 6104 11830 6132 12242
rect 6288 11898 6316 12310
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6092 11824 6144 11830
rect 6092 11766 6144 11772
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6380 10810 6408 11154
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 5998 10296 6054 10305
rect 5998 10231 6054 10240
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6104 9042 6132 10406
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6380 9722 6408 10066
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6104 8634 6132 8978
rect 6472 8634 6500 8978
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5446 8256 5502 8265
rect 5446 8191 5502 8200
rect 5460 7886 5488 8191
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7410 5488 7686
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5552 6866 5580 8434
rect 5814 8392 5870 8401
rect 5814 8327 5870 8336
rect 5828 8090 5856 8327
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 6012 6916 6040 7210
rect 6104 7041 6132 8570
rect 6366 8528 6422 8537
rect 6472 8514 6500 8570
rect 6564 8537 6592 12566
rect 6656 9518 6684 12854
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6422 8486 6500 8514
rect 6550 8528 6606 8537
rect 6366 8463 6422 8472
rect 6550 8463 6606 8472
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 6288 7546 6316 7958
rect 6552 7880 6604 7886
rect 6550 7848 6552 7857
rect 6604 7848 6606 7857
rect 6550 7783 6606 7792
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6090 7032 6146 7041
rect 6090 6967 6146 6976
rect 6092 6928 6144 6934
rect 6012 6888 6092 6916
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5552 6458 5580 6802
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 6012 6118 6040 6888
rect 6092 6870 6144 6876
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6012 5846 6040 6054
rect 6274 5944 6330 5953
rect 6274 5879 6276 5888
rect 6328 5879 6330 5888
rect 6276 5850 6328 5856
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 5908 5704 5960 5710
rect 5906 5672 5908 5681
rect 5960 5672 5962 5681
rect 5906 5607 5962 5616
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6012 5166 6040 5782
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5644 4758 5672 5034
rect 6366 4992 6422 5001
rect 6366 4927 6422 4936
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6380 4321 6408 4927
rect 6748 4690 6776 22442
rect 7484 22234 7512 22578
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 6920 22160 6972 22166
rect 6920 22102 6972 22108
rect 7470 22128 7526 22137
rect 6828 21344 6880 21350
rect 6932 21298 6960 22102
rect 7470 22063 7526 22072
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 7300 21418 7328 21626
rect 7288 21412 7340 21418
rect 7288 21354 7340 21360
rect 7380 21412 7432 21418
rect 7380 21354 7432 21360
rect 6880 21292 6960 21298
rect 6828 21286 6960 21292
rect 6840 21270 6960 21286
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 6840 17921 6868 20470
rect 6932 20058 6960 21270
rect 7392 21146 7420 21354
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7012 20800 7064 20806
rect 7012 20742 7064 20748
rect 7024 20398 7052 20742
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 7024 18426 7052 18770
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 7024 18329 7052 18362
rect 7104 18352 7156 18358
rect 7010 18320 7066 18329
rect 6920 18284 6972 18290
rect 7104 18294 7156 18300
rect 7010 18255 7066 18264
rect 6920 18226 6972 18232
rect 6826 17912 6882 17921
rect 6826 17847 6882 17856
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6840 16794 6868 17614
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6932 16674 6960 18226
rect 6840 16646 6960 16674
rect 6840 16590 6868 16646
rect 6828 16584 6880 16590
rect 7116 16538 7144 18294
rect 7484 18272 7512 22063
rect 7576 22030 7604 22578
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 7576 21554 7604 21966
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7562 19816 7618 19825
rect 7562 19751 7618 19760
rect 6828 16526 6880 16532
rect 6932 16510 7144 16538
rect 7392 18244 7512 18272
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6840 14890 6868 15574
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6840 12238 6868 12718
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6840 10033 6868 11630
rect 6932 11540 6960 16510
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 7024 15162 7052 15506
rect 7194 15464 7250 15473
rect 7194 15399 7250 15408
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 7024 12306 7052 14894
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7116 12102 7144 12650
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7012 11552 7064 11558
rect 6932 11520 7012 11540
rect 7064 11520 7066 11529
rect 6932 11512 7010 11520
rect 7010 11455 7066 11464
rect 6918 10296 6974 10305
rect 6918 10231 6974 10240
rect 6932 10062 6960 10231
rect 7024 10130 7052 11455
rect 7116 11286 7144 12038
rect 7208 11762 7236 15399
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 13802 7328 14214
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7300 13530 7328 13738
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7208 11354 7236 11698
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7208 10810 7236 11086
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7300 10674 7328 12718
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6920 10056 6972 10062
rect 6826 10024 6882 10033
rect 6920 9998 6972 10004
rect 6826 9959 6882 9968
rect 7286 9616 7342 9625
rect 7286 9551 7342 9560
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7024 8634 7052 9318
rect 7116 8838 7144 9454
rect 7300 9217 7328 9551
rect 7286 9208 7342 9217
rect 7286 9143 7342 9152
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6932 7313 6960 7346
rect 7116 7342 7144 8774
rect 7104 7336 7156 7342
rect 6918 7304 6974 7313
rect 6918 7239 6974 7248
rect 7102 7304 7104 7313
rect 7288 7336 7340 7342
rect 7156 7304 7158 7313
rect 7288 7278 7340 7284
rect 7102 7239 7158 7248
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 7194 7168 7250 7177
rect 6932 5914 6960 7142
rect 7194 7103 7250 7112
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6920 5908 6972 5914
rect 6840 5868 6920 5896
rect 6840 5234 6868 5868
rect 6920 5850 6972 5856
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6932 5370 6960 5646
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6932 4826 6960 5102
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6366 4312 6422 4321
rect 5356 4276 5408 4282
rect 6366 4247 6422 4256
rect 5356 4218 5408 4224
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5552 3126 5580 3946
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5998 2952 6054 2961
rect 5998 2887 6054 2896
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5460 2009 5488 2246
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5446 2000 5502 2009
rect 5446 1935 5502 1944
rect 6012 1737 6040 2887
rect 6104 2650 6132 3878
rect 6380 3738 6408 4247
rect 6748 4214 6776 4626
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6932 4128 6960 4762
rect 6840 4100 6960 4128
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6196 3194 6224 3538
rect 6840 3194 6868 4100
rect 7024 4026 7052 6258
rect 6932 4010 7052 4026
rect 6920 4004 7052 4010
rect 6972 3998 7052 4004
rect 6920 3946 6972 3952
rect 6932 3466 6960 3946
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 5998 1728 6054 1737
rect 5998 1663 6054 1672
rect 6196 480 6224 3130
rect 7024 2990 7052 3334
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7208 480 7236 7103
rect 7300 6905 7328 7278
rect 7286 6896 7342 6905
rect 7286 6831 7342 6840
rect 7300 6798 7328 6831
rect 7392 6798 7420 18244
rect 7472 18148 7524 18154
rect 7472 18090 7524 18096
rect 7484 17882 7512 18090
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7470 16824 7526 16833
rect 7470 16759 7526 16768
rect 7484 16114 7512 16759
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7484 13530 7512 13942
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7576 11558 7604 19751
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7668 11370 7696 22918
rect 8298 22879 8354 22888
rect 7840 22704 7892 22710
rect 7840 22646 7892 22652
rect 7748 22432 7800 22438
rect 7748 22374 7800 22380
rect 7760 20602 7788 22374
rect 7852 22137 7880 22646
rect 7838 22128 7894 22137
rect 7838 22063 7894 22072
rect 8024 21956 8076 21962
rect 8024 21898 8076 21904
rect 8036 21146 8064 21898
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 8036 21049 8064 21082
rect 8022 21040 8078 21049
rect 8022 20975 8078 20984
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 7760 19310 7788 19654
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7760 19145 7788 19246
rect 7746 19136 7802 19145
rect 7746 19071 7802 19080
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7760 18601 7788 18770
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 7746 18592 7802 18601
rect 7746 18527 7802 18536
rect 7760 18358 7788 18527
rect 7748 18352 7800 18358
rect 7748 18294 7800 18300
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 7944 17338 7972 17750
rect 8036 17338 8064 18702
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 8128 18086 8156 18566
rect 8208 18284 8260 18290
rect 8312 18272 8340 22879
rect 8588 22778 8616 23122
rect 8760 22976 8812 22982
rect 8760 22918 8812 22924
rect 8576 22772 8628 22778
rect 8576 22714 8628 22720
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 8680 21350 8708 22374
rect 8772 22234 8800 22918
rect 8850 22536 8906 22545
rect 8850 22471 8906 22480
rect 8864 22273 8892 22471
rect 8850 22264 8906 22273
rect 8760 22228 8812 22234
rect 8850 22199 8906 22208
rect 8760 22170 8812 22176
rect 8772 21622 8800 22170
rect 8760 21616 8812 21622
rect 8760 21558 8812 21564
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8390 19408 8446 19417
rect 8390 19343 8446 19352
rect 8404 18737 8432 19343
rect 8680 19310 8708 21286
rect 8864 21010 8892 22199
rect 9128 22092 9180 22098
rect 9128 22034 9180 22040
rect 9140 21554 9168 22034
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 8852 21004 8904 21010
rect 8852 20946 8904 20952
rect 8864 20602 8892 20946
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 9048 20466 9076 20742
rect 9140 20466 9168 21490
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 8772 19854 8800 20266
rect 9048 20058 9076 20402
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 9232 19417 9260 24806
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10690 24304 10746 24313
rect 10690 24239 10692 24248
rect 10744 24239 10746 24248
rect 10692 24210 10744 24216
rect 10048 24064 10100 24070
rect 10048 24006 10100 24012
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 9864 23248 9916 23254
rect 9864 23190 9916 23196
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9784 22778 9812 23054
rect 9588 22772 9640 22778
rect 9588 22714 9640 22720
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9312 22500 9364 22506
rect 9312 22442 9364 22448
rect 9324 21894 9352 22442
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9508 21078 9536 21966
rect 9600 21570 9628 22714
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9692 21962 9720 22578
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9692 21690 9720 21898
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9600 21542 9720 21570
rect 9496 21072 9548 21078
rect 9496 21014 9548 21020
rect 9692 21026 9720 21542
rect 9784 21146 9812 22714
rect 9876 22438 9904 23190
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 9876 21690 9904 22374
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9692 20998 9812 21026
rect 9678 19952 9734 19961
rect 9404 19916 9456 19922
rect 9678 19887 9680 19896
rect 9404 19858 9456 19864
rect 9732 19887 9734 19896
rect 9680 19858 9732 19864
rect 9218 19408 9274 19417
rect 9416 19378 9444 19858
rect 9692 19446 9720 19858
rect 9680 19440 9732 19446
rect 9680 19382 9732 19388
rect 9218 19343 9274 19352
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 8666 19000 8722 19009
rect 8666 18935 8722 18944
rect 8680 18834 8708 18935
rect 9324 18902 9352 19110
rect 8944 18896 8996 18902
rect 8944 18838 8996 18844
rect 9312 18896 9364 18902
rect 9416 18873 9444 19314
rect 9496 19304 9548 19310
rect 9494 19272 9496 19281
rect 9548 19272 9550 19281
rect 9494 19207 9550 19216
rect 9508 18970 9536 19207
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9312 18838 9364 18844
rect 9402 18864 9458 18873
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8390 18728 8446 18737
rect 8390 18663 8446 18672
rect 8260 18244 8340 18272
rect 8208 18226 8260 18232
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 8128 17649 8156 18022
rect 8312 17814 8340 18244
rect 8680 18222 8708 18770
rect 8668 18216 8720 18222
rect 8666 18184 8668 18193
rect 8720 18184 8722 18193
rect 8666 18119 8722 18128
rect 8482 17912 8538 17921
rect 8482 17847 8538 17856
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8114 17640 8170 17649
rect 8114 17575 8170 17584
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7944 16794 7972 17274
rect 8128 17218 8156 17575
rect 8036 17190 8156 17218
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7840 16720 7892 16726
rect 7840 16662 7892 16668
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7760 15366 7788 16526
rect 7852 16250 7880 16662
rect 8036 16590 8064 17190
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7852 15978 7880 16186
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 7852 15706 7880 15914
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7760 14550 7788 14758
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 8036 14414 8064 16526
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 8128 15706 8156 16050
rect 8116 15700 8168 15706
rect 8116 15642 8168 15648
rect 8208 15360 8260 15366
rect 8260 15320 8340 15348
rect 8208 15302 8260 15308
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 7944 13190 7972 14350
rect 8128 14074 8156 14486
rect 8312 14074 8340 15320
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8404 13870 8432 16390
rect 8496 15570 8524 17847
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8680 16794 8708 17614
rect 8956 17066 8984 18838
rect 9402 18799 9458 18808
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 9048 18426 9076 18634
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9048 18222 9076 18362
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 8944 17060 8996 17066
rect 8944 17002 8996 17008
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8680 16590 8708 16730
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8680 16114 8708 16526
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8496 14822 8524 15506
rect 8680 15026 8708 16050
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8484 14816 8536 14822
rect 8680 14793 8708 14826
rect 8484 14758 8536 14764
rect 8666 14784 8722 14793
rect 8496 14249 8524 14758
rect 8666 14719 8722 14728
rect 8680 14618 8708 14719
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8772 14550 8800 14826
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 8482 14240 8538 14249
rect 8482 14175 8538 14184
rect 8758 14104 8814 14113
rect 8758 14039 8814 14048
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8220 13682 8248 13806
rect 8220 13654 8340 13682
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 7932 13184 7984 13190
rect 7930 13152 7932 13161
rect 7984 13152 7986 13161
rect 7930 13087 7986 13096
rect 8128 12986 8156 13262
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8220 12850 8248 13398
rect 8312 13326 8340 13654
rect 8300 13320 8352 13326
rect 8298 13288 8300 13297
rect 8352 13288 8354 13297
rect 8298 13223 8354 13232
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11626 8064 12038
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7484 11342 7696 11370
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7300 6361 7328 6598
rect 7392 6458 7420 6734
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7286 6352 7342 6361
rect 7286 6287 7342 6296
rect 7484 5216 7512 11342
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7668 10810 7696 11222
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7760 10554 7788 11494
rect 8036 11354 8064 11562
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 7838 10704 7894 10713
rect 7838 10639 7840 10648
rect 7892 10639 7894 10648
rect 7840 10610 7892 10616
rect 7760 10526 7880 10554
rect 8036 10538 8064 11290
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7668 9042 7696 9454
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7668 8838 7696 8978
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7668 6730 7696 6870
rect 7656 6724 7708 6730
rect 7656 6666 7708 6672
rect 7668 6458 7696 6666
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7576 5846 7604 6258
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 7760 5778 7788 8026
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7392 5188 7512 5216
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7300 4146 7328 4694
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7392 4026 7420 5188
rect 7760 5166 7788 5714
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7472 5092 7524 5098
rect 7472 5034 7524 5040
rect 7484 4622 7512 5034
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 4758 7788 4966
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7300 3998 7420 4026
rect 7300 3738 7328 3998
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7300 3534 7328 3674
rect 7392 3670 7420 3878
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7392 3194 7420 3606
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7484 2689 7512 4558
rect 7760 4282 7788 4694
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7470 2680 7526 2689
rect 7470 2615 7526 2624
rect 7668 2582 7696 4082
rect 7748 3664 7800 3670
rect 7746 3632 7748 3641
rect 7800 3632 7802 3641
rect 7746 3567 7802 3576
rect 7852 2650 7880 10526
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 8036 10266 8064 10474
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8404 10130 8432 11154
rect 8496 10713 8524 12922
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8588 11898 8616 12242
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8680 11762 8708 13942
rect 8772 12986 8800 14039
rect 9140 13802 9168 16118
rect 9232 13954 9260 18158
rect 9312 15904 9364 15910
rect 9310 15872 9312 15881
rect 9364 15872 9366 15881
rect 9310 15807 9366 15816
rect 9232 13926 9352 13954
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9140 13530 9168 13738
rect 9232 13734 9260 13806
rect 9324 13734 9352 13926
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9232 13297 9260 13670
rect 9218 13288 9274 13297
rect 9416 13258 9444 18799
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 16250 9536 16934
rect 9600 16726 9628 18566
rect 9784 18306 9812 20998
rect 9692 18278 9812 18306
rect 9588 16720 9640 16726
rect 9588 16662 9640 16668
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9600 15706 9628 16662
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9586 15600 9642 15609
rect 9586 15535 9588 15544
rect 9640 15535 9642 15544
rect 9588 15506 9640 15512
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9600 13530 9628 14350
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9218 13223 9274 13232
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8850 12064 8906 12073
rect 8850 11999 8906 12008
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8482 10704 8538 10713
rect 8482 10639 8538 10648
rect 8496 10606 8524 10639
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8036 9722 8064 10066
rect 8404 9722 8432 10066
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7944 8362 7972 9046
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8208 8832 8260 8838
rect 8576 8832 8628 8838
rect 8260 8780 8340 8786
rect 8208 8774 8340 8780
rect 8576 8774 8628 8780
rect 8220 8758 8340 8774
rect 7932 8356 7984 8362
rect 7932 8298 7984 8304
rect 7944 8090 7972 8298
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 8312 7954 8340 8758
rect 8588 8634 8616 8774
rect 8680 8634 8708 8910
rect 8772 8838 8800 9386
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8760 8016 8812 8022
rect 8758 7984 8760 7993
rect 8812 7984 8814 7993
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8668 7948 8720 7954
rect 8758 7919 8814 7928
rect 8668 7890 8720 7896
rect 7944 7410 7972 7890
rect 8298 7848 8354 7857
rect 8024 7812 8076 7818
rect 8298 7783 8354 7792
rect 8024 7754 8076 7760
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 8036 6798 8064 7754
rect 8312 7546 8340 7783
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8298 7440 8354 7449
rect 8298 7375 8354 7384
rect 8206 7168 8262 7177
rect 8206 7103 8262 7112
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8036 6322 8064 6734
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7944 5914 7972 6054
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8036 5098 8064 6258
rect 8220 6254 8248 7103
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8220 5098 8248 5646
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 8312 4146 8340 7375
rect 8390 7032 8446 7041
rect 8390 6967 8446 6976
rect 8404 5409 8432 6967
rect 8574 6896 8630 6905
rect 8574 6831 8630 6840
rect 8390 5400 8446 5409
rect 8390 5335 8392 5344
rect 8444 5335 8446 5344
rect 8392 5306 8444 5312
rect 8404 5166 8432 5306
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8588 5148 8616 6831
rect 8680 6662 8708 7890
rect 8760 7880 8812 7886
rect 8758 7848 8760 7857
rect 8812 7848 8814 7857
rect 8758 7783 8814 7792
rect 8864 7546 8892 11999
rect 8956 11830 8984 12174
rect 8944 11824 8996 11830
rect 8942 11792 8944 11801
rect 8996 11792 8998 11801
rect 8942 11727 8998 11736
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8956 8634 8984 8842
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8864 7342 8892 7482
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 9048 6934 9076 12378
rect 9600 12306 9628 13466
rect 9692 13190 9720 18278
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9784 17882 9812 18158
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9784 17134 9812 17818
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9876 17082 9904 21490
rect 9968 20602 9996 23462
rect 10060 21554 10088 24006
rect 10704 23866 10732 24210
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 10152 22642 10180 23054
rect 10140 22636 10192 22642
rect 10140 22578 10192 22584
rect 10796 22574 10824 25758
rect 11518 24712 11574 24721
rect 11518 24647 11574 24656
rect 11150 24440 11206 24449
rect 11150 24375 11206 24384
rect 11164 23662 11192 24375
rect 11152 23656 11204 23662
rect 11152 23598 11204 23604
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10784 22568 10836 22574
rect 10784 22510 10836 22516
rect 10692 22432 10744 22438
rect 10692 22374 10744 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10140 22160 10192 22166
rect 10140 22102 10192 22108
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 10152 21434 10180 22102
rect 10704 22030 10732 22374
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10060 21406 10180 21434
rect 10060 21350 10088 21406
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 10060 20806 10088 21286
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10704 21078 10732 21626
rect 10692 21072 10744 21078
rect 10506 21040 10562 21049
rect 10744 21020 10824 21026
rect 10692 21014 10824 21020
rect 10704 20998 10824 21014
rect 10506 20975 10562 20984
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 10060 20330 10088 20742
rect 10520 20466 10548 20975
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10048 20324 10100 20330
rect 10048 20266 10100 20272
rect 9956 19984 10008 19990
rect 9956 19926 10008 19932
rect 9968 19242 9996 19926
rect 10060 19514 10088 20266
rect 10704 20262 10732 20878
rect 10796 20602 10824 20998
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10704 20058 10732 20198
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10796 19922 10824 20538
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9968 18902 9996 19178
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 10152 18850 10180 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10888 18902 10916 20402
rect 10324 18896 10376 18902
rect 10152 18844 10324 18850
rect 10152 18838 10376 18844
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10152 18822 10364 18838
rect 10046 18592 10102 18601
rect 10046 18527 10102 18536
rect 10060 18086 10088 18527
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10152 17882 10180 18822
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10140 17264 10192 17270
rect 10140 17206 10192 17212
rect 9876 17054 10088 17082
rect 9772 16992 9824 16998
rect 9956 16992 10008 16998
rect 9824 16952 9904 16980
rect 9772 16934 9824 16940
rect 9876 16726 9904 16952
rect 9956 16934 10008 16940
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9770 15736 9826 15745
rect 9770 15671 9826 15680
rect 9784 15570 9812 15671
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9784 15162 9812 15506
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9784 14482 9812 15098
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9784 14074 9812 14418
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9876 13462 9904 15846
rect 9968 15570 9996 16934
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9968 15094 9996 15506
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 9968 14793 9996 15030
rect 9954 14784 10010 14793
rect 9954 14719 10010 14728
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9784 12764 9812 13262
rect 9692 12736 9812 12764
rect 9692 12374 9720 12736
rect 9876 12714 9904 13398
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9784 12374 9812 12582
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9876 11626 9904 12650
rect 9968 12442 9996 14554
rect 10060 12646 10088 17054
rect 10152 16590 10180 17206
rect 10796 17066 10824 17750
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10690 16416 10746 16425
rect 10690 16351 10746 16360
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10612 15201 10640 15438
rect 10598 15192 10654 15201
rect 10598 15127 10654 15136
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10152 13802 10180 14214
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10152 13530 10180 13738
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10152 12714 10180 13466
rect 10322 13016 10378 13025
rect 10322 12951 10378 12960
rect 10336 12850 10364 12951
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10046 12472 10102 12481
rect 9956 12436 10008 12442
rect 10152 12442 10180 12650
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10046 12407 10102 12416
rect 10140 12436 10192 12442
rect 9956 12378 10008 12384
rect 9968 11762 9996 12378
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9416 11286 9444 11494
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9324 10198 9352 10542
rect 9416 10538 9444 11222
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9692 10674 9720 11154
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9692 10441 9720 10610
rect 9678 10432 9734 10441
rect 9678 10367 9734 10376
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 8945 9260 9318
rect 9218 8936 9274 8945
rect 9218 8871 9220 8880
rect 9272 8871 9274 8880
rect 9404 8900 9456 8906
rect 9220 8842 9272 8848
rect 9404 8842 9456 8848
rect 9416 8362 9444 8842
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9508 8362 9536 8570
rect 9600 8498 9628 9386
rect 9770 9344 9826 9353
rect 9770 9279 9826 9288
rect 9784 8838 9812 9279
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9416 7750 9444 8298
rect 9600 8265 9628 8434
rect 9876 8362 9904 8910
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9586 8256 9642 8265
rect 9586 8191 9642 8200
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9416 7449 9444 7686
rect 9402 7440 9458 7449
rect 9402 7375 9458 7384
rect 9692 7274 9720 7686
rect 9784 7410 9812 7822
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9036 6928 9088 6934
rect 9036 6870 9088 6876
rect 8852 6792 8904 6798
rect 8850 6760 8852 6769
rect 8904 6760 8906 6769
rect 8850 6695 8906 6704
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8680 5681 8708 6598
rect 9048 6458 9076 6870
rect 9600 6798 9628 7210
rect 9784 7002 9812 7346
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9692 6730 9720 6802
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9692 6458 9720 6666
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 8666 5672 8722 5681
rect 8666 5607 8722 5616
rect 9034 5264 9090 5273
rect 9034 5199 9090 5208
rect 8668 5160 8720 5166
rect 8588 5120 8668 5148
rect 8588 4826 8616 5120
rect 8668 5102 8720 5108
rect 9048 4826 9076 5199
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 8942 4584 8998 4593
rect 8942 4519 8998 4528
rect 8956 4486 8984 4519
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 4146 8984 4422
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 8576 4072 8628 4078
rect 8114 4040 8170 4049
rect 8114 3975 8170 3984
rect 8574 4040 8576 4049
rect 8628 4040 8630 4049
rect 8574 3975 8630 3984
rect 8128 3233 8156 3975
rect 9048 3398 9076 4082
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 8114 3224 8170 3233
rect 8114 3159 8170 3168
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7852 2446 7880 2586
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 8128 480 8156 3159
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8300 2576 8352 2582
rect 8298 2544 8300 2553
rect 8588 2553 8616 2994
rect 8666 2816 8722 2825
rect 8666 2751 8722 2760
rect 8680 2650 8708 2751
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8352 2544 8354 2553
rect 8298 2479 8354 2488
rect 8574 2544 8630 2553
rect 8574 2479 8630 2488
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 8864 1465 8892 2246
rect 8850 1456 8906 1465
rect 8850 1391 8906 1400
rect 9140 480 9168 3946
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9232 2990 9260 3606
rect 9324 3058 9352 6394
rect 9772 6112 9824 6118
rect 9876 6089 9904 8298
rect 9968 6730 9996 11018
rect 10060 10062 10088 12407
rect 10140 12378 10192 12384
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10612 11898 10640 12310
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10152 10198 10180 10406
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10060 9178 10088 9998
rect 10152 9722 10180 10134
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10152 9382 10180 9658
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10244 9489 10272 9522
rect 10230 9480 10286 9489
rect 10230 9415 10232 9424
rect 10284 9415 10286 9424
rect 10232 9386 10284 9392
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 10046 8936 10102 8945
rect 10046 8871 10102 8880
rect 10060 7478 10088 8871
rect 10152 8294 10180 9046
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10152 7750 10180 8230
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 10506 6352 10562 6361
rect 10506 6287 10562 6296
rect 10520 6254 10548 6287
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10140 6112 10192 6118
rect 9772 6054 9824 6060
rect 9862 6080 9918 6089
rect 9784 5710 9812 6054
rect 10140 6054 10192 6060
rect 9862 6015 9918 6024
rect 10152 5817 10180 6054
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10138 5808 10194 5817
rect 10138 5743 10194 5752
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9692 5030 9720 5578
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9402 4720 9458 4729
rect 9402 4655 9404 4664
rect 9456 4655 9458 4664
rect 9404 4626 9456 4632
rect 9416 4214 9444 4626
rect 9692 4486 9720 4966
rect 9680 4480 9732 4486
rect 9784 4457 9812 5306
rect 9876 4758 9904 5510
rect 10428 5302 10456 5510
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 10048 5092 10100 5098
rect 10048 5034 10100 5040
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9968 4865 9996 4966
rect 9954 4856 10010 4865
rect 9954 4791 10010 4800
rect 9864 4752 9916 4758
rect 9864 4694 9916 4700
rect 9680 4422 9732 4428
rect 9770 4448 9826 4457
rect 9692 4321 9720 4422
rect 9770 4383 9826 4392
rect 9678 4312 9734 4321
rect 9678 4247 9680 4256
rect 9732 4247 9734 4256
rect 9680 4218 9732 4224
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9416 3738 9444 4150
rect 9692 4078 9720 4218
rect 9680 4072 9732 4078
rect 9586 4040 9642 4049
rect 9680 4014 9732 4020
rect 9586 3975 9642 3984
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9416 3534 9444 3674
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9600 2650 9628 3975
rect 9692 3738 9720 4014
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9784 3194 9812 4383
rect 9876 3466 9904 4694
rect 9864 3460 9916 3466
rect 9864 3402 9916 3408
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9876 2990 9904 3402
rect 9968 3194 9996 4791
rect 10060 4282 10088 5034
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10060 3670 10088 4218
rect 10152 4146 10180 5238
rect 10520 5234 10548 5646
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10704 4758 10732 16351
rect 10796 16250 10824 17002
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10888 13977 10916 18090
rect 10980 17678 11008 23462
rect 11164 23322 11192 23598
rect 11152 23316 11204 23322
rect 11152 23258 11204 23264
rect 11336 23180 11388 23186
rect 11336 23122 11388 23128
rect 11152 22976 11204 22982
rect 11152 22918 11204 22924
rect 11164 22234 11192 22918
rect 11348 22438 11376 23122
rect 11336 22432 11388 22438
rect 11334 22400 11336 22409
rect 11388 22400 11390 22409
rect 11334 22335 11390 22344
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 11164 21554 11192 22170
rect 11334 22128 11390 22137
rect 11532 22098 11560 24647
rect 11808 24313 11836 27520
rect 13188 24449 13216 27520
rect 13174 24440 13230 24449
rect 13174 24375 13230 24384
rect 11794 24304 11850 24313
rect 11612 24268 11664 24274
rect 11794 24239 11850 24248
rect 12438 24304 12494 24313
rect 12438 24239 12494 24248
rect 11612 24210 11664 24216
rect 11624 23526 11652 24210
rect 11888 24064 11940 24070
rect 11888 24006 11940 24012
rect 11612 23520 11664 23526
rect 11612 23462 11664 23468
rect 11624 22114 11652 23462
rect 11334 22063 11390 22072
rect 11520 22092 11572 22098
rect 11152 21548 11204 21554
rect 11152 21490 11204 21496
rect 11150 21040 11206 21049
rect 11150 20975 11152 20984
rect 11204 20975 11206 20984
rect 11152 20946 11204 20952
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11242 19136 11298 19145
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 11058 17640 11114 17649
rect 10980 16726 11008 17614
rect 11058 17575 11060 17584
rect 11112 17575 11114 17584
rect 11060 17546 11112 17552
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11072 16794 11100 17138
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 11058 16688 11114 16697
rect 11058 16623 11114 16632
rect 11072 14657 11100 16623
rect 11058 14648 11114 14657
rect 11058 14583 11114 14592
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11072 14074 11100 14418
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10874 13968 10930 13977
rect 10874 13903 10930 13912
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 11058 13832 11114 13841
rect 10874 13560 10930 13569
rect 10874 13495 10930 13504
rect 10784 13320 10836 13326
rect 10888 13297 10916 13495
rect 10784 13262 10836 13268
rect 10874 13288 10930 13297
rect 10796 12986 10824 13262
rect 10874 13223 10930 13232
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10796 10713 10824 12106
rect 10888 11558 10916 12310
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 11286 10916 11494
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10888 10810 10916 11222
rect 10980 11132 11008 13806
rect 11058 13767 11114 13776
rect 11072 13530 11100 13767
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 11058 13288 11114 13297
rect 11058 13223 11060 13232
rect 11112 13223 11114 13232
rect 11060 13194 11112 13200
rect 11058 13152 11114 13161
rect 11058 13087 11114 13096
rect 11072 12850 11100 13087
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 11072 12170 11100 12650
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 11060 11688 11112 11694
rect 11058 11656 11060 11665
rect 11112 11656 11114 11665
rect 11058 11591 11114 11600
rect 11060 11144 11112 11150
rect 10980 11104 11060 11132
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10782 10704 10838 10713
rect 10782 10639 10838 10648
rect 10796 9654 10824 10639
rect 10980 10198 11008 11104
rect 11060 11086 11112 11092
rect 10968 10192 11020 10198
rect 10968 10134 11020 10140
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10874 8256 10930 8265
rect 10874 8191 10930 8200
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10796 6254 10824 6802
rect 10888 6730 10916 8191
rect 11060 7336 11112 7342
rect 10980 7296 11060 7324
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10980 5914 11008 7296
rect 11060 7278 11112 7284
rect 11058 7168 11114 7177
rect 11058 7103 11114 7112
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10796 5030 10824 5510
rect 10888 5098 10916 5510
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 10876 5092 10928 5098
rect 10876 5034 10928 5040
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10796 4826 10824 4966
rect 10980 4826 11008 5306
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10796 4282 10824 4490
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10152 3738 10180 4082
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 10796 3602 10824 4218
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10520 3126 10548 3334
rect 10796 3194 10824 3538
rect 10980 3398 11008 4762
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10980 3194 11008 3334
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10508 3120 10560 3126
rect 10692 3120 10744 3126
rect 10508 3062 10560 3068
rect 10690 3088 10692 3097
rect 10744 3088 10746 3097
rect 10690 3023 10746 3032
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9496 2440 9548 2446
rect 9494 2408 9496 2417
rect 9548 2408 9550 2417
rect 9494 2343 9550 2352
rect 9784 2009 9812 2450
rect 10796 2446 10824 3130
rect 10980 2961 11008 3130
rect 10966 2952 11022 2961
rect 10966 2887 11022 2896
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 9968 2009 9996 2246
rect 9770 2000 9826 2009
rect 9770 1935 9826 1944
rect 9954 2000 10010 2009
rect 9954 1935 10010 1944
rect 10060 480 10088 2246
rect 10796 1465 10824 2382
rect 10782 1456 10838 1465
rect 10782 1391 10838 1400
rect 11072 480 11100 7103
rect 11164 5370 11192 19110
rect 11242 19071 11298 19080
rect 11256 18970 11284 19071
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11348 16810 11376 22063
rect 11624 22086 11698 22114
rect 11520 22034 11572 22040
rect 11532 22001 11560 22034
rect 11670 22012 11698 22086
rect 11518 21992 11574 22001
rect 11518 21927 11574 21936
rect 11624 21984 11698 22012
rect 11532 21690 11560 21927
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11440 18290 11468 19110
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11440 16998 11468 17682
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11256 16782 11376 16810
rect 11256 12782 11284 16782
rect 11336 16720 11388 16726
rect 11336 16662 11388 16668
rect 11348 16250 11376 16662
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11348 15042 11376 15506
rect 11440 15162 11468 16934
rect 11532 16697 11560 18362
rect 11518 16688 11574 16697
rect 11518 16623 11574 16632
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11532 15910 11560 16526
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11532 15609 11560 15846
rect 11518 15600 11574 15609
rect 11518 15535 11574 15544
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11348 15014 11468 15042
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11348 14618 11376 14894
rect 11440 14890 11468 15014
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11334 14104 11390 14113
rect 11334 14039 11390 14048
rect 11348 13841 11376 14039
rect 11334 13832 11390 13841
rect 11334 13767 11390 13776
rect 11336 13728 11388 13734
rect 11440 13682 11468 14826
rect 11388 13676 11468 13682
rect 11336 13670 11468 13676
rect 11348 13654 11468 13670
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11242 12200 11298 12209
rect 11242 12135 11298 12144
rect 11256 11150 11284 12135
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11256 10266 11284 10950
rect 11348 10810 11376 13654
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11440 12986 11468 13330
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11426 11792 11482 11801
rect 11426 11727 11482 11736
rect 11440 11257 11468 11727
rect 11518 11656 11574 11665
rect 11518 11591 11574 11600
rect 11532 11558 11560 11591
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11426 11248 11482 11257
rect 11426 11183 11482 11192
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11256 8362 11284 8910
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11256 7970 11284 8298
rect 11256 7942 11376 7970
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11256 6662 11284 7822
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11256 6322 11284 6598
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11348 4826 11376 7942
rect 11440 7546 11468 11086
rect 11624 8809 11652 21984
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11808 18426 11836 18770
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 11704 18080 11756 18086
rect 11756 18040 11836 18068
rect 11704 18022 11756 18028
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 11716 16590 11744 17546
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11716 14074 11744 14418
rect 11808 14414 11836 18040
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11702 13424 11758 13433
rect 11702 13359 11758 13368
rect 11610 8800 11666 8809
rect 11610 8735 11666 8744
rect 11716 8634 11744 13359
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11808 10130 11836 13126
rect 11900 11014 11928 24006
rect 12452 23662 12480 24239
rect 14554 24168 14610 24177
rect 14554 24103 14610 24112
rect 14568 23866 14596 24103
rect 14556 23860 14608 23866
rect 14556 23802 14608 23808
rect 14278 23760 14334 23769
rect 14278 23695 14334 23704
rect 12440 23656 12492 23662
rect 13820 23656 13872 23662
rect 12440 23598 12492 23604
rect 12714 23624 12770 23633
rect 13820 23598 13872 23604
rect 12714 23559 12770 23568
rect 12256 23180 12308 23186
rect 12256 23122 12308 23128
rect 12162 22808 12218 22817
rect 12162 22743 12218 22752
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 12084 20602 12112 20946
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 12084 20369 12112 20538
rect 12070 20360 12126 20369
rect 12070 20295 12126 20304
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11992 19174 12020 19858
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11992 17649 12020 19110
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 11978 17640 12034 17649
rect 11978 17575 12034 17584
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 11992 15162 12020 15506
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11992 14958 12020 15098
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 12084 14414 12112 18566
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 12084 13462 12112 13670
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11992 10248 12020 12922
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 12084 11393 12112 12718
rect 12070 11384 12126 11393
rect 12070 11319 12126 11328
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12084 10470 12112 11154
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 11900 10220 12020 10248
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11808 9722 11836 10066
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11900 9625 11928 10220
rect 12084 10169 12112 10406
rect 12070 10160 12126 10169
rect 12070 10095 12126 10104
rect 11886 9616 11942 9625
rect 11886 9551 11942 9560
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11716 8430 11744 8570
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11716 8022 11744 8230
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11716 7750 11744 7958
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11716 7206 11744 7686
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11624 6458 11652 6802
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11518 5128 11574 5137
rect 11518 5063 11574 5072
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 2650 11192 4422
rect 11336 4072 11388 4078
rect 11334 4040 11336 4049
rect 11388 4040 11390 4049
rect 11334 3975 11390 3984
rect 11440 3942 11468 4966
rect 11532 4690 11560 5063
rect 11716 5030 11744 7142
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11532 4282 11560 4626
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11256 2825 11284 3334
rect 11348 2990 11376 3470
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11242 2816 11298 2825
rect 11242 2751 11298 2760
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11150 2544 11206 2553
rect 11150 2479 11152 2488
rect 11204 2479 11206 2488
rect 11428 2508 11480 2514
rect 11152 2450 11204 2456
rect 11428 2450 11480 2456
rect 11440 2417 11468 2450
rect 11426 2408 11482 2417
rect 11426 2343 11482 2352
rect 11992 480 12020 9114
rect 12176 8786 12204 22743
rect 12268 22642 12296 23122
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12360 22234 12388 22918
rect 12438 22672 12494 22681
rect 12438 22607 12494 22616
rect 12452 22574 12480 22607
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12348 22228 12400 22234
rect 12348 22170 12400 22176
rect 12728 21457 12756 23559
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 12808 22500 12860 22506
rect 12808 22442 12860 22448
rect 12820 21554 12848 22442
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12808 21548 12860 21554
rect 12808 21490 12860 21496
rect 12714 21448 12770 21457
rect 12912 21418 12940 21830
rect 12714 21383 12770 21392
rect 12900 21412 12952 21418
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12636 20602 12664 20946
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12452 19378 12480 19790
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12268 18086 12296 18294
rect 12348 18284 12400 18290
rect 12452 18272 12480 19314
rect 12544 19310 12572 19654
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12400 18244 12480 18272
rect 12348 18226 12400 18232
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 12268 15706 12296 18022
rect 12544 17678 12572 19246
rect 12636 18970 12664 20538
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12636 18154 12664 18906
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12636 17746 12664 18090
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12636 17270 12664 17682
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12346 17096 12402 17105
rect 12346 17031 12402 17040
rect 12360 16726 12388 17031
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12440 16788 12492 16794
rect 12440 16730 12492 16736
rect 12348 16720 12400 16726
rect 12348 16662 12400 16668
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12360 15570 12388 16662
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12268 14550 12296 15438
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 12360 15026 12388 15302
rect 12452 15162 12480 16730
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 12438 13968 12494 13977
rect 12438 13903 12440 13912
rect 12492 13903 12494 13912
rect 12440 13874 12492 13880
rect 12452 13530 12480 13874
rect 12544 13841 12572 16934
rect 12622 15192 12678 15201
rect 12728 15162 12756 21383
rect 12900 21354 12952 21360
rect 13096 19281 13124 22374
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13280 20466 13308 20878
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13082 19272 13138 19281
rect 13082 19207 13138 19216
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13188 18154 13216 18702
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 13188 17882 13216 18090
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12912 17513 12940 17682
rect 12898 17504 12954 17513
rect 12898 17439 12954 17448
rect 12912 16998 12940 17439
rect 13268 17128 13320 17134
rect 13266 17096 13268 17105
rect 13320 17096 13322 17105
rect 13266 17031 13322 17040
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12622 15127 12678 15136
rect 12716 15156 12768 15162
rect 12530 13832 12586 13841
rect 12530 13767 12586 13776
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12452 12730 12480 12786
rect 12084 8758 12204 8786
rect 12268 12702 12480 12730
rect 12084 6905 12112 8758
rect 12268 8650 12296 12702
rect 12346 12608 12402 12617
rect 12346 12543 12402 12552
rect 12360 10266 12388 12543
rect 12438 12336 12494 12345
rect 12438 12271 12494 12280
rect 12452 12238 12480 12271
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12544 11694 12572 13767
rect 12636 13394 12664 15127
rect 12716 15098 12768 15104
rect 12728 14958 12756 15098
rect 12716 14952 12768 14958
rect 12768 14912 12848 14940
rect 12716 14894 12768 14900
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12728 13818 12756 14758
rect 12820 13954 12848 14912
rect 12912 14822 12940 16934
rect 13280 16726 13308 17031
rect 13268 16720 13320 16726
rect 13268 16662 13320 16668
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 13096 15638 13124 15982
rect 13188 15706 13216 16526
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13280 15638 13308 15846
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13280 14822 13308 15574
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12912 14074 12940 14350
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13004 14006 13032 14486
rect 12992 14000 13044 14006
rect 12820 13926 12940 13954
rect 12992 13942 13044 13948
rect 12728 13790 12848 13818
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12636 12442 12664 13330
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12728 12073 12756 12718
rect 12714 12064 12770 12073
rect 12714 11999 12770 12008
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12544 11354 12572 11630
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12820 11286 12848 13790
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12532 11144 12584 11150
rect 12820 11121 12848 11222
rect 12532 11086 12584 11092
rect 12806 11112 12862 11121
rect 12544 10674 12572 11086
rect 12806 11047 12862 11056
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12176 8622 12296 8650
rect 12176 8566 12204 8622
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12452 8276 12480 10202
rect 12544 9489 12572 10610
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12636 10266 12664 10474
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12714 10160 12770 10169
rect 12714 10095 12716 10104
rect 12768 10095 12770 10104
rect 12716 10066 12768 10072
rect 12530 9480 12586 9489
rect 12530 9415 12586 9424
rect 12820 9110 12848 10746
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12544 8362 12572 9046
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12360 8248 12480 8276
rect 12360 8090 12388 8248
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12162 7168 12218 7177
rect 12162 7103 12218 7112
rect 12070 6896 12126 6905
rect 12070 6831 12072 6840
rect 12124 6831 12126 6840
rect 12072 6802 12124 6808
rect 12084 6771 12112 6802
rect 12072 5772 12124 5778
rect 12176 5760 12204 7103
rect 12452 6866 12480 8248
rect 12806 7712 12862 7721
rect 12806 7647 12862 7656
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12452 6458 12480 6802
rect 12636 6798 12664 7142
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12820 6254 12848 7647
rect 12912 7313 12940 13926
rect 12992 13456 13044 13462
rect 13096 13444 13124 14758
rect 13044 13416 13124 13444
rect 12992 13398 13044 13404
rect 13004 12918 13032 13398
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 13004 12374 13032 12854
rect 12992 12368 13044 12374
rect 12992 12310 13044 12316
rect 13084 12232 13136 12238
rect 12990 12200 13046 12209
rect 13084 12174 13136 12180
rect 12990 12135 13046 12144
rect 13004 11694 13032 12135
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 13096 11354 13124 12174
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 13280 11218 13308 11562
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13280 10266 13308 11154
rect 13372 10674 13400 23462
rect 13832 23338 13860 23598
rect 13740 23322 13860 23338
rect 13728 23316 13860 23322
rect 13780 23310 13860 23316
rect 13728 23258 13780 23264
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13556 22953 13584 23122
rect 13542 22944 13598 22953
rect 13542 22879 13598 22888
rect 13556 22778 13584 22879
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 13452 22024 13504 22030
rect 13452 21966 13504 21972
rect 13464 21554 13492 21966
rect 13648 21690 13676 22102
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13544 21412 13596 21418
rect 13544 21354 13596 21360
rect 13556 21049 13584 21354
rect 13542 21040 13598 21049
rect 13542 20975 13598 20984
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13464 19990 13492 20198
rect 13452 19984 13504 19990
rect 13452 19926 13504 19932
rect 13464 19174 13492 19926
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13464 18902 13492 19110
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13464 18086 13492 18838
rect 13556 18834 13584 20975
rect 13648 19310 13676 21626
rect 13728 20936 13780 20942
rect 13832 20890 13860 22646
rect 14002 22536 14058 22545
rect 14002 22471 14004 22480
rect 14056 22471 14058 22480
rect 14004 22442 14056 22448
rect 13912 21616 13964 21622
rect 13912 21558 13964 21564
rect 13924 21078 13952 21558
rect 14188 21344 14240 21350
rect 14188 21286 14240 21292
rect 13912 21072 13964 21078
rect 13912 21014 13964 21020
rect 13780 20884 13860 20890
rect 13728 20878 13860 20884
rect 13740 20862 13860 20878
rect 13832 20058 13860 20862
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13924 19922 13952 21014
rect 14200 20602 14228 21286
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 14188 18216 14240 18222
rect 14292 18193 14320 23695
rect 14660 23497 14688 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14738 24848 14794 24857
rect 14738 24783 14794 24792
rect 14646 23488 14702 23497
rect 14646 23423 14702 23432
rect 14752 23338 14780 24783
rect 16040 24177 16068 27520
rect 17130 24440 17186 24449
rect 17130 24375 17132 24384
rect 17184 24375 17186 24384
rect 17132 24346 17184 24352
rect 17316 24268 17368 24274
rect 17316 24210 17368 24216
rect 16026 24168 16082 24177
rect 16026 24103 16082 24112
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 16210 23896 16266 23905
rect 16210 23831 16212 23840
rect 16264 23831 16266 23840
rect 16212 23802 16264 23808
rect 16028 23656 16080 23662
rect 16026 23624 16028 23633
rect 16080 23624 16082 23633
rect 16026 23559 16082 23568
rect 17328 23526 17356 24210
rect 17420 23905 17448 27520
rect 18328 26648 18380 26654
rect 18328 26590 18380 26596
rect 18234 24712 18290 24721
rect 18234 24647 18290 24656
rect 18248 24410 18276 24647
rect 18236 24404 18288 24410
rect 18236 24346 18288 24352
rect 18234 24304 18290 24313
rect 18234 24239 18290 24248
rect 17406 23896 17462 23905
rect 18248 23866 18276 24239
rect 17406 23831 17462 23840
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 18144 23656 18196 23662
rect 18144 23598 18196 23604
rect 17316 23520 17368 23526
rect 16762 23488 16818 23497
rect 17316 23462 17368 23468
rect 16762 23423 16818 23432
rect 14660 23310 14780 23338
rect 14464 22568 14516 22574
rect 14464 22510 14516 22516
rect 14476 22001 14504 22510
rect 14462 21992 14518 22001
rect 14518 21950 14596 21978
rect 14462 21927 14518 21936
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14384 21078 14412 21490
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14476 19922 14504 20198
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14188 18158 14240 18164
rect 14278 18184 14334 18193
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13910 18048 13966 18057
rect 13464 17066 13492 18022
rect 13542 17912 13598 17921
rect 13542 17847 13598 17856
rect 13556 17746 13584 17847
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13832 17270 13860 18022
rect 13910 17983 13966 17992
rect 13820 17264 13872 17270
rect 13542 17232 13598 17241
rect 13820 17206 13872 17212
rect 13542 17167 13598 17176
rect 13452 17060 13504 17066
rect 13452 17002 13504 17008
rect 13464 16726 13492 17002
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13464 15978 13492 16662
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13556 15858 13584 17167
rect 13464 15830 13584 15858
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13188 9722 13216 10134
rect 13372 10062 13400 10474
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13188 9602 13216 9658
rect 13188 9574 13308 9602
rect 13372 9586 13400 9998
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13188 8906 13216 9386
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13280 8634 13308 9574
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13372 8945 13400 9522
rect 13358 8936 13414 8945
rect 13358 8871 13414 8880
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 13004 8090 13032 8366
rect 13280 8090 13308 8570
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13004 7993 13032 8026
rect 12990 7984 13046 7993
rect 12990 7919 13046 7928
rect 13280 7546 13308 8026
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13174 7440 13230 7449
rect 13174 7375 13230 7384
rect 12898 7304 12954 7313
rect 12898 7239 12954 7248
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12124 5732 12204 5760
rect 12624 5772 12676 5778
rect 12072 5714 12124 5720
rect 12624 5714 12676 5720
rect 12084 5409 12112 5714
rect 12162 5672 12218 5681
rect 12162 5607 12218 5616
rect 12070 5400 12126 5409
rect 12070 5335 12072 5344
rect 12124 5335 12126 5344
rect 12072 5306 12124 5312
rect 12176 4690 12204 5607
rect 12636 5370 12664 5714
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12176 4282 12204 4626
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12164 3664 12216 3670
rect 12162 3632 12164 3641
rect 12216 3632 12218 3641
rect 12162 3567 12218 3576
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12162 3224 12218 3233
rect 12268 3210 12296 3538
rect 12218 3182 12296 3210
rect 12162 3159 12164 3168
rect 12216 3159 12218 3168
rect 12164 3130 12216 3136
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12452 2938 12480 2994
rect 12360 2910 12480 2938
rect 12360 2582 12388 2910
rect 12544 2689 12572 5102
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12636 3641 12664 3878
rect 12622 3632 12678 3641
rect 12622 3567 12678 3576
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12820 3058 12848 3334
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12530 2680 12586 2689
rect 12530 2615 12532 2624
rect 12584 2615 12586 2624
rect 12532 2586 12584 2592
rect 12348 2576 12400 2582
rect 12544 2555 12572 2586
rect 12636 2582 12664 2790
rect 12624 2576 12676 2582
rect 12348 2518 12400 2524
rect 12624 2518 12676 2524
rect 12636 2310 12664 2518
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12728 1601 12756 2382
rect 12912 1601 12940 2926
rect 12714 1592 12770 1601
rect 12714 1527 12770 1536
rect 12898 1592 12954 1601
rect 12898 1527 12954 1536
rect 13004 480 13032 7142
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13096 5846 13124 6734
rect 13188 6730 13216 7375
rect 13464 7274 13492 15830
rect 13924 15026 13952 17983
rect 14200 17814 14228 18158
rect 14278 18119 14334 18128
rect 14188 17808 14240 17814
rect 14188 17750 14240 17756
rect 14200 16794 14228 17750
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14292 15722 14320 18119
rect 14016 15694 14320 15722
rect 13912 15020 13964 15026
rect 13832 14980 13912 15008
rect 13832 14618 13860 14980
rect 13912 14962 13964 14968
rect 13912 14884 13964 14890
rect 13912 14826 13964 14832
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13820 14408 13872 14414
rect 13740 14368 13820 14396
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 13556 12986 13584 14282
rect 13636 14000 13688 14006
rect 13634 13968 13636 13977
rect 13688 13968 13690 13977
rect 13634 13903 13690 13912
rect 13740 13954 13768 14368
rect 13924 14396 13952 14826
rect 13872 14368 13952 14396
rect 13820 14350 13872 14356
rect 13820 14000 13872 14006
rect 13740 13948 13820 13954
rect 13740 13942 13872 13948
rect 13740 13926 13860 13942
rect 13740 13530 13768 13926
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13832 12850 13860 13126
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13740 12442 13768 12650
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 11286 13768 11494
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13740 10810 13768 11222
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13464 5914 13492 6054
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 13082 5264 13138 5273
rect 13082 5199 13138 5208
rect 13096 4146 13124 5199
rect 13556 5001 13584 10610
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13740 9602 13768 9930
rect 14016 9722 14044 15694
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14108 14550 14136 14962
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 14108 12850 14136 14486
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14108 12238 14136 12786
rect 14384 12458 14412 19314
rect 14568 18737 14596 21950
rect 14554 18728 14610 18737
rect 14554 18663 14610 18672
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14568 17202 14596 17478
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14660 17082 14688 23310
rect 15566 23216 15622 23225
rect 16776 23186 16804 23423
rect 15566 23151 15568 23160
rect 15620 23151 15622 23160
rect 16764 23180 16816 23186
rect 15568 23122 15620 23128
rect 16764 23122 16816 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15580 22778 15608 23122
rect 15936 22976 15988 22982
rect 15936 22918 15988 22924
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15660 22432 15712 22438
rect 15660 22374 15712 22380
rect 15568 22160 15620 22166
rect 15568 22102 15620 22108
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15016 21412 15068 21418
rect 15016 21354 15068 21360
rect 15028 20913 15056 21354
rect 15580 21350 15608 22102
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15580 21049 15608 21286
rect 15672 21078 15700 22374
rect 15752 21956 15804 21962
rect 15752 21898 15804 21904
rect 15660 21072 15712 21078
rect 15566 21040 15622 21049
rect 15660 21014 15712 21020
rect 15566 20975 15622 20984
rect 15014 20904 15070 20913
rect 15014 20839 15070 20848
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15672 20602 15700 21014
rect 15764 20806 15792 21898
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15856 21146 15884 21626
rect 15948 21554 15976 22918
rect 16776 22778 16804 23122
rect 16764 22772 16816 22778
rect 16764 22714 16816 22720
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 15844 21140 15896 21146
rect 15844 21082 15896 21088
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15566 20496 15622 20505
rect 15566 20431 15568 20440
rect 15620 20431 15622 20440
rect 15568 20402 15620 20408
rect 14740 20392 14792 20398
rect 14740 20334 14792 20340
rect 14752 19446 14780 20334
rect 15764 20330 15792 20742
rect 15752 20324 15804 20330
rect 15752 20266 15804 20272
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14752 18630 14780 19246
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14752 18290 14780 18566
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14200 12430 14412 12458
rect 14476 17054 14688 17082
rect 14752 17066 14780 18022
rect 14740 17060 14792 17066
rect 14200 12288 14228 12430
rect 14200 12260 14320 12288
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14186 12200 14242 12209
rect 14186 12135 14242 12144
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14108 11694 14136 12038
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 14108 10713 14136 11630
rect 14094 10704 14150 10713
rect 14094 10639 14150 10648
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 13740 9574 13860 9602
rect 13832 9382 13860 9574
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 13740 9110 13768 9318
rect 13728 9104 13780 9110
rect 13726 9072 13728 9081
rect 13780 9072 13782 9081
rect 13726 9007 13782 9016
rect 14108 8945 14136 9318
rect 14094 8936 14150 8945
rect 13728 8900 13780 8906
rect 14094 8871 14150 8880
rect 13728 8842 13780 8848
rect 13634 8392 13690 8401
rect 13634 8327 13636 8336
rect 13688 8327 13690 8336
rect 13636 8298 13688 8304
rect 13648 7478 13676 8298
rect 13740 8276 13768 8842
rect 13910 8800 13966 8809
rect 13910 8735 13966 8744
rect 13924 8430 13952 8735
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13740 8248 13860 8276
rect 13728 8016 13780 8022
rect 13726 7984 13728 7993
rect 13780 7984 13782 7993
rect 13726 7919 13782 7928
rect 13636 7472 13688 7478
rect 13636 7414 13688 7420
rect 13832 7274 13860 8248
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13832 7002 13860 7210
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13832 6322 13860 6598
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13542 4992 13598 5001
rect 13542 4927 13598 4936
rect 13832 4826 13860 5782
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13636 4752 13688 4758
rect 13636 4694 13688 4700
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13280 1873 13308 4422
rect 13648 3942 13676 4694
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13648 2650 13676 3878
rect 13832 3670 13860 4762
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13832 3194 13860 3606
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13266 1864 13322 1873
rect 13266 1799 13322 1808
rect 13924 480 13952 8366
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14016 7449 14044 7822
rect 14002 7440 14058 7449
rect 14002 7375 14004 7384
rect 14056 7375 14058 7384
rect 14004 7346 14056 7352
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 14016 5370 14044 7210
rect 14200 6440 14228 12135
rect 14292 10146 14320 12260
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14384 10266 14412 10542
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14292 10118 14412 10146
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14292 8548 14320 9522
rect 14384 9217 14412 10118
rect 14370 9208 14426 9217
rect 14370 9143 14426 9152
rect 14476 9042 14504 17054
rect 14740 17002 14792 17008
rect 14646 16552 14702 16561
rect 14646 16487 14702 16496
rect 14740 16516 14792 16522
rect 14660 16114 14688 16487
rect 14740 16458 14792 16464
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14752 15910 14780 16458
rect 14844 16130 14872 20198
rect 15856 20058 15884 21082
rect 16132 20942 16160 21558
rect 16120 20936 16172 20942
rect 16684 20913 16712 22510
rect 17328 22409 17356 23462
rect 18052 23180 18104 23186
rect 18052 23122 18104 23128
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17314 22400 17370 22409
rect 17314 22335 17370 22344
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 16960 21418 16988 21966
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16948 21412 17000 21418
rect 16948 21354 17000 21360
rect 16776 21146 16804 21354
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16120 20878 16172 20884
rect 16670 20904 16726 20913
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15658 19272 15714 19281
rect 15658 19207 15714 19216
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15304 17814 15332 18702
rect 15580 18086 15608 18838
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15304 16726 15332 16934
rect 15292 16720 15344 16726
rect 15292 16662 15344 16668
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15488 16182 15516 16526
rect 15476 16176 15528 16182
rect 14844 16114 15240 16130
rect 15476 16118 15528 16124
rect 14844 16108 15252 16114
rect 14844 16102 15200 16108
rect 15200 16050 15252 16056
rect 14740 15904 14792 15910
rect 14792 15864 14872 15892
rect 14740 15846 14792 15852
rect 14844 15706 14872 15864
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14740 15632 14792 15638
rect 14740 15574 14792 15580
rect 14752 15366 14780 15574
rect 15488 15502 15516 16118
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14752 15162 14780 15302
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14646 14240 14702 14249
rect 14646 14175 14702 14184
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14568 12646 14596 13262
rect 14556 12640 14608 12646
rect 14554 12608 14556 12617
rect 14608 12608 14610 12617
rect 14554 12543 14610 12552
rect 14660 11098 14688 14175
rect 14844 13530 14872 14350
rect 15304 14346 15332 15370
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15396 13977 15424 14826
rect 15672 14532 15700 19207
rect 15856 18426 15884 19994
rect 16132 19854 16160 20878
rect 16670 20839 16726 20848
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16592 20346 16620 20742
rect 16684 20466 16712 20839
rect 16776 20602 16804 21082
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16500 20330 16620 20346
rect 16488 20324 16620 20330
rect 16540 20318 16620 20324
rect 16488 20266 16540 20272
rect 16212 19984 16264 19990
rect 16212 19926 16264 19932
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16132 19378 16160 19790
rect 16224 19514 16252 19926
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16500 18970 16528 20266
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16028 18896 16080 18902
rect 16028 18838 16080 18844
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15856 18154 15884 18362
rect 16040 18290 16068 18838
rect 16592 18358 16620 20198
rect 16684 19786 16712 20402
rect 16868 19990 16896 21286
rect 16856 19984 16908 19990
rect 16856 19926 16908 19932
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17040 18828 17092 18834
rect 17040 18770 17092 18776
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 17052 18086 17080 18770
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 17052 17921 17080 18022
rect 17038 17912 17094 17921
rect 16120 17876 16172 17882
rect 17038 17847 17094 17856
rect 16120 17818 16172 17824
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15764 16998 15792 17682
rect 16132 17202 16160 17818
rect 16948 17808 17000 17814
rect 16948 17750 17000 17756
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15764 16096 15792 16934
rect 16500 16833 16528 17478
rect 16486 16824 16542 16833
rect 16684 16794 16712 17682
rect 16960 17066 16988 17750
rect 17144 17746 17172 18906
rect 17236 18873 17264 19110
rect 17222 18864 17278 18873
rect 17222 18799 17278 18808
rect 17328 17785 17356 22335
rect 17314 17776 17370 17785
rect 17132 17740 17184 17746
rect 17314 17711 17370 17720
rect 17132 17682 17184 17688
rect 17130 17640 17186 17649
rect 17130 17575 17186 17584
rect 16948 17060 17000 17066
rect 16948 17002 17000 17008
rect 16486 16759 16542 16768
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15856 16250 15884 16662
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 16408 16204 16620 16232
rect 15764 16068 15884 16096
rect 15474 14512 15530 14521
rect 15672 14504 15792 14532
rect 15474 14447 15530 14456
rect 15488 14414 15516 14447
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15382 13968 15438 13977
rect 15200 13932 15252 13938
rect 15382 13903 15438 13912
rect 15200 13874 15252 13880
rect 15212 13841 15240 13874
rect 15198 13832 15254 13841
rect 15198 13767 15254 13776
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 15396 13462 15424 13903
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15396 12986 15424 13398
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15474 12608 15530 12617
rect 15474 12543 15530 12552
rect 15384 12368 15436 12374
rect 15304 12316 15384 12322
rect 15304 12310 15436 12316
rect 15304 12294 15424 12310
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14752 11218 14780 12174
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11558 15332 12294
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15304 11354 15332 11494
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14660 11070 14780 11098
rect 14646 10432 14702 10441
rect 14646 10367 14702 10376
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14476 8634 14504 8978
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14372 8560 14424 8566
rect 14292 8520 14372 8548
rect 14292 7324 14320 8520
rect 14372 8502 14424 8508
rect 14476 7449 14504 8570
rect 14462 7440 14518 7449
rect 14462 7375 14518 7384
rect 14292 7296 14504 7324
rect 14200 6412 14320 6440
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 14200 5642 14228 6258
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 14200 4758 14228 5578
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14292 3738 14320 6412
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14188 3528 14240 3534
rect 14292 3516 14320 3674
rect 14384 3670 14412 4082
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 14240 3488 14320 3516
rect 14188 3470 14240 3476
rect 14476 2038 14504 7296
rect 14660 6866 14688 10367
rect 14752 7818 14780 11070
rect 14844 10266 14872 11222
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15396 10810 15424 11698
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15212 10266 15240 10406
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 15382 9480 15438 9489
rect 14844 8838 14872 9454
rect 15382 9415 15438 9424
rect 15396 9382 15424 9415
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15108 8084 15160 8090
rect 15212 8072 15240 8434
rect 15160 8044 15240 8072
rect 15108 8026 15160 8032
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 15382 7712 15438 7721
rect 14956 7644 15252 7664
rect 15382 7647 15438 7656
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15396 7342 15424 7647
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15028 7206 15056 7278
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15028 7041 15056 7142
rect 15014 7032 15070 7041
rect 15014 6967 15070 6976
rect 15488 6866 15516 12543
rect 15580 11286 15608 12786
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15672 10266 15700 11222
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15764 10130 15792 14504
rect 15856 12356 15884 16068
rect 16304 16040 16356 16046
rect 16408 16028 16436 16204
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16356 16000 16436 16028
rect 16304 15982 16356 15988
rect 16500 15706 16528 16050
rect 16592 15978 16620 16204
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16118 15464 16174 15473
rect 16118 15399 16174 15408
rect 15936 15088 15988 15094
rect 15936 15030 15988 15036
rect 15948 13938 15976 15030
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 16040 13462 16068 14350
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15948 12714 15976 12854
rect 16040 12850 16068 13398
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 16132 12730 16160 15399
rect 16592 15094 16620 15914
rect 16764 15632 16816 15638
rect 16764 15574 16816 15580
rect 16776 15162 16804 15574
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16580 15088 16632 15094
rect 16394 15056 16450 15065
rect 16580 15030 16632 15036
rect 17144 15026 17172 17575
rect 17222 15600 17278 15609
rect 17222 15535 17278 15544
rect 17236 15502 17264 15535
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 16394 14991 16396 15000
rect 16448 14991 16450 15000
rect 17132 15020 17184 15026
rect 16396 14962 16448 14968
rect 17132 14962 17184 14968
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 16040 12702 16160 12730
rect 16040 12374 16068 12702
rect 16028 12368 16080 12374
rect 15856 12328 15976 12356
rect 15842 11112 15898 11121
rect 15842 11047 15898 11056
rect 15856 10810 15884 11047
rect 15948 10996 15976 12328
rect 16028 12310 16080 12316
rect 16212 12368 16264 12374
rect 16212 12310 16264 12316
rect 16040 11762 16068 12310
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16040 11150 16068 11698
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15948 10968 16068 10996
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15856 10606 15884 10746
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15672 9602 15700 9998
rect 15764 9722 15792 10066
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15672 9574 15792 9602
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 15580 8634 15608 9386
rect 15764 9382 15792 9574
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15764 8378 15792 9318
rect 15856 8498 15884 9998
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15764 8350 15884 8378
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15580 7546 15608 7890
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15580 7313 15608 7482
rect 15752 7336 15804 7342
rect 15566 7304 15622 7313
rect 15752 7278 15804 7284
rect 15566 7239 15622 7248
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 14660 6458 14688 6802
rect 15304 6769 15332 6802
rect 15290 6760 15346 6769
rect 15290 6695 15346 6704
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15304 6458 15332 6695
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14660 5370 14688 6122
rect 15568 5840 15620 5846
rect 14738 5808 14794 5817
rect 15568 5782 15620 5788
rect 14738 5743 14740 5752
rect 14792 5743 14794 5752
rect 14740 5714 14792 5720
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14752 5234 14780 5714
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14844 4826 14872 5646
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15580 5012 15608 5782
rect 15672 5234 15700 7142
rect 15764 6934 15792 7278
rect 15752 6928 15804 6934
rect 15752 6870 15804 6876
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 6186 15792 6598
rect 15856 6497 15884 8350
rect 16040 7585 16068 10968
rect 16224 9178 16252 12310
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 16132 8838 16160 9046
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16120 8832 16172 8838
rect 16224 8809 16252 8910
rect 16120 8774 16172 8780
rect 16210 8800 16266 8809
rect 16132 8294 16160 8774
rect 16210 8735 16266 8744
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16132 8090 16160 8230
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16026 7576 16082 7585
rect 16026 7511 16082 7520
rect 15842 6488 15898 6497
rect 15842 6423 15898 6432
rect 16040 6390 16068 7511
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15660 5024 15712 5030
rect 15580 4984 15660 5012
rect 15660 4966 15712 4972
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 15672 4486 15700 4966
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15396 4049 15424 4150
rect 15382 4040 15438 4049
rect 15382 3975 15384 3984
rect 15436 3975 15438 3984
rect 15384 3946 15436 3952
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14554 3088 14610 3097
rect 14554 3023 14610 3032
rect 14568 2990 14596 3023
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 14568 2650 14596 2926
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14464 2032 14516 2038
rect 14464 1974 14516 1980
rect 14924 2032 14976 2038
rect 14924 1974 14976 1980
rect 14936 480 14964 1974
rect 15396 1873 15424 3470
rect 15488 3194 15516 3606
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15672 2922 15700 4422
rect 16132 4282 16160 4694
rect 16224 4622 16252 6122
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16224 4214 16252 4558
rect 16212 4208 16264 4214
rect 16212 4150 16264 4156
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 15474 2816 15530 2825
rect 15474 2751 15530 2760
rect 15488 2514 15516 2751
rect 15658 2680 15714 2689
rect 15658 2615 15660 2624
rect 15712 2615 15714 2624
rect 15660 2586 15712 2592
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15382 1864 15438 1873
rect 15382 1799 15438 1808
rect 15856 480 15884 4082
rect 16224 3670 16252 4150
rect 16316 4146 16344 14894
rect 16946 14784 17002 14793
rect 16946 14719 17002 14728
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16394 12744 16450 12753
rect 16394 12679 16450 12688
rect 16408 12646 16436 12679
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16408 12442 16436 12582
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16868 12374 16896 13806
rect 16856 12368 16908 12374
rect 16856 12310 16908 12316
rect 16580 9920 16632 9926
rect 16500 9868 16580 9874
rect 16500 9862 16632 9868
rect 16500 9846 16620 9862
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16408 8838 16436 9386
rect 16500 9382 16528 9846
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16592 8362 16620 8910
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16580 8356 16632 8362
rect 16500 8316 16580 8344
rect 16500 8022 16528 8316
rect 16580 8298 16632 8304
rect 16776 8022 16804 8366
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16764 8016 16816 8022
rect 16764 7958 16816 7964
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16396 6656 16448 6662
rect 16500 6633 16528 6802
rect 16396 6598 16448 6604
rect 16486 6624 16542 6633
rect 16408 6322 16436 6598
rect 16486 6559 16542 6568
rect 16500 6458 16528 6559
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 16408 3233 16436 6258
rect 16500 6225 16528 6394
rect 16486 6216 16542 6225
rect 16486 6151 16542 6160
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16592 4758 16620 4966
rect 16580 4752 16632 4758
rect 16684 4729 16712 7754
rect 16776 7206 16804 7958
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16868 6905 16896 7278
rect 16854 6896 16910 6905
rect 16764 6860 16816 6866
rect 16854 6831 16910 6840
rect 16764 6802 16816 6808
rect 16776 6322 16804 6802
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16580 4694 16632 4700
rect 16670 4720 16726 4729
rect 16670 4655 16726 4664
rect 16868 4264 16896 6831
rect 16960 6458 16988 14719
rect 17236 14618 17264 15438
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17328 14498 17356 17711
rect 17420 14550 17448 22918
rect 18064 22710 18092 23122
rect 18052 22704 18104 22710
rect 18052 22646 18104 22652
rect 18156 21486 18184 23598
rect 18340 23322 18368 26590
rect 18800 24449 18828 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 20180 24721 20208 27520
rect 20166 24712 20222 24721
rect 20166 24647 20222 24656
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 18786 24440 18842 24449
rect 19622 24432 19918 24452
rect 18786 24375 18842 24384
rect 18696 24268 18748 24274
rect 18696 24210 18748 24216
rect 18708 23526 18736 24210
rect 21454 24032 21510 24041
rect 21454 23967 21510 23976
rect 20350 23896 20406 23905
rect 21468 23866 21496 23967
rect 21652 23905 21680 27520
rect 22558 24168 22614 24177
rect 22558 24103 22614 24112
rect 21638 23896 21694 23905
rect 20350 23831 20352 23840
rect 20404 23831 20406 23840
rect 21456 23860 21508 23866
rect 20352 23802 20404 23808
rect 22572 23866 22600 24103
rect 23032 24041 23060 27520
rect 24412 27418 24440 27520
rect 24228 27390 24440 27418
rect 23478 27296 23534 27305
rect 23478 27231 23534 27240
rect 23492 26654 23520 27231
rect 23480 26648 23532 26654
rect 23480 26590 23532 26596
rect 24228 24177 24256 27390
rect 24766 25936 24822 25945
rect 24766 25871 24822 25880
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24674 24576 24730 24585
rect 24674 24511 24730 24520
rect 24214 24168 24270 24177
rect 24214 24103 24270 24112
rect 23018 24032 23074 24041
rect 23018 23967 23074 23976
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 21638 23831 21694 23840
rect 22560 23860 22612 23866
rect 21456 23802 21508 23808
rect 22560 23802 22612 23808
rect 21270 23760 21326 23769
rect 21270 23695 21326 23704
rect 21284 23662 21312 23695
rect 21272 23656 21324 23662
rect 21272 23598 21324 23604
rect 22192 23656 22244 23662
rect 22192 23598 22244 23604
rect 24584 23656 24636 23662
rect 24584 23598 24636 23604
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 18328 23316 18380 23322
rect 18328 23258 18380 23264
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 17868 21412 17920 21418
rect 17868 21354 17920 21360
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17880 21298 17908 21354
rect 17512 21078 17540 21286
rect 17880 21270 18000 21298
rect 17500 21072 17552 21078
rect 17500 21014 17552 21020
rect 17512 20602 17540 21014
rect 17972 20602 18000 21270
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 18708 20398 18736 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18696 20392 18748 20398
rect 18696 20334 18748 20340
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 17868 19984 17920 19990
rect 17868 19926 17920 19932
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17590 19408 17646 19417
rect 17590 19343 17646 19352
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17512 16726 17540 17478
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17512 16250 17540 16662
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17236 14470 17356 14498
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 17236 13870 17264 14470
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17316 13796 17368 13802
rect 17316 13738 17368 13744
rect 17130 13560 17186 13569
rect 17130 13495 17186 13504
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 17052 12714 17080 13398
rect 17144 12889 17172 13495
rect 17328 13326 17356 13738
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17130 12880 17186 12889
rect 17130 12815 17186 12824
rect 17040 12708 17092 12714
rect 17040 12650 17092 12656
rect 17236 12646 17264 13262
rect 17224 12640 17276 12646
rect 17222 12608 17224 12617
rect 17276 12608 17278 12617
rect 17222 12543 17278 12552
rect 17328 11898 17356 13262
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17420 11762 17448 12310
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17038 11656 17094 11665
rect 17038 11591 17094 11600
rect 17052 10810 17080 11591
rect 17420 11286 17448 11698
rect 17408 11280 17460 11286
rect 17314 11248 17370 11257
rect 17408 11222 17460 11228
rect 17314 11183 17316 11192
rect 17368 11183 17370 11192
rect 17316 11154 17368 11160
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17328 10266 17356 11154
rect 17420 10742 17448 11222
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17512 9722 17540 10134
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 17052 8634 17080 9046
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17052 8090 17080 8570
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17328 7886 17356 9590
rect 17408 9512 17460 9518
rect 17406 9480 17408 9489
rect 17460 9480 17462 9489
rect 17406 9415 17462 9424
rect 17512 9110 17540 9658
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17328 7478 17356 7822
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 17420 7002 17448 7890
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17604 6769 17632 19343
rect 17696 19242 17724 19790
rect 17788 19310 17816 19790
rect 17880 19514 17908 19926
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 17776 19304 17828 19310
rect 17972 19258 18000 19654
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 17776 19246 17828 19252
rect 17684 19236 17736 19242
rect 17684 19178 17736 19184
rect 17880 19230 18000 19258
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17696 18970 17724 19178
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17880 18902 17908 19230
rect 17960 19168 18012 19174
rect 17958 19136 17960 19145
rect 18012 19136 18014 19145
rect 17958 19071 18014 19080
rect 17868 18896 17920 18902
rect 17868 18838 17920 18844
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17788 18086 17816 18770
rect 18064 18766 18092 19246
rect 18052 18760 18104 18766
rect 17880 18708 18052 18714
rect 17880 18702 18104 18708
rect 17880 18686 18092 18702
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 17788 17814 17816 18022
rect 17776 17808 17828 17814
rect 17776 17750 17828 17756
rect 17788 17134 17816 17750
rect 17776 17128 17828 17134
rect 17774 17096 17776 17105
rect 17828 17096 17830 17105
rect 17774 17031 17830 17040
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17696 15638 17724 16526
rect 17684 15632 17736 15638
rect 17684 15574 17736 15580
rect 17880 15484 17908 18686
rect 18064 18637 18092 18686
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 17270 18276 17478
rect 18236 17264 18288 17270
rect 18236 17206 18288 17212
rect 18248 17066 18276 17206
rect 18144 17060 18196 17066
rect 18144 17002 18196 17008
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 18156 16794 18184 17002
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18234 16688 18290 16697
rect 18234 16623 18290 16632
rect 18248 15706 18276 16623
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 17696 15456 17908 15484
rect 17696 13308 17724 15456
rect 18248 15026 18276 15642
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17880 13530 17908 14554
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17696 13280 17816 13308
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17696 11558 17724 12174
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17696 11121 17724 11494
rect 17682 11112 17738 11121
rect 17682 11047 17738 11056
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17696 9382 17724 9998
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 7546 17724 9318
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17590 6760 17646 6769
rect 17590 6695 17646 6704
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17040 5636 17092 5642
rect 17040 5578 17092 5584
rect 17052 4486 17080 5578
rect 17236 5370 17264 5782
rect 17420 5681 17448 6054
rect 17406 5672 17462 5681
rect 17316 5636 17368 5642
rect 17406 5607 17462 5616
rect 17316 5578 17368 5584
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 17328 4758 17356 5578
rect 17590 5128 17646 5137
rect 17590 5063 17646 5072
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17316 4752 17368 4758
rect 17316 4694 17368 4700
rect 17512 4690 17540 4966
rect 17604 4826 17632 5063
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16868 4236 16988 4264
rect 16854 4176 16910 4185
rect 16854 4111 16910 4120
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16592 3738 16620 3946
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16868 3670 16896 4111
rect 16856 3664 16908 3670
rect 16856 3606 16908 3612
rect 16394 3224 16450 3233
rect 16394 3159 16450 3168
rect 16868 3058 16896 3606
rect 16960 3602 16988 4236
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16960 3194 16988 3538
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 17052 3058 17080 4422
rect 17512 4282 17540 4626
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17604 4214 17632 4762
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 16224 2650 16252 2858
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16500 2281 16528 2382
rect 16486 2272 16542 2281
rect 16486 2207 16542 2216
rect 17130 2136 17186 2145
rect 17130 2071 17186 2080
rect 17144 1737 17172 2071
rect 17328 1737 17356 3334
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17420 2650 17448 2790
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17130 1728 17186 1737
rect 17130 1663 17186 1672
rect 17314 1728 17370 1737
rect 17314 1663 17370 1672
rect 16856 604 16908 610
rect 16856 546 16908 552
rect 16868 480 16896 546
rect 17788 480 17816 13280
rect 17972 12850 18000 14826
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 18064 14006 18092 14486
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 18064 13818 18092 13942
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18064 13802 18184 13818
rect 18064 13796 18196 13802
rect 18064 13790 18144 13796
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 18064 12442 18092 13790
rect 18144 13738 18196 13744
rect 18248 13530 18276 13874
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18156 12306 18184 12786
rect 18340 12617 18368 19314
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18432 17202 18460 18158
rect 18524 17241 18552 20198
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18510 17232 18566 17241
rect 18420 17196 18472 17202
rect 18510 17167 18566 17176
rect 18420 17138 18472 17144
rect 18432 16590 18460 17138
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18616 16114 18644 18566
rect 18708 18086 18736 18770
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18708 16998 18736 17682
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18616 15706 18644 16050
rect 18604 15700 18656 15706
rect 18604 15642 18656 15648
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18616 14793 18644 15438
rect 18602 14784 18658 14793
rect 18602 14719 18658 14728
rect 18604 13456 18656 13462
rect 18604 13398 18656 13404
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 18326 12608 18382 12617
rect 18326 12543 18382 12552
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18432 11354 18460 12650
rect 18524 12646 18552 13262
rect 18616 12714 18644 13398
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18602 12608 18658 12617
rect 18524 12442 18552 12582
rect 18602 12543 18658 12552
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17866 9480 17922 9489
rect 17866 9415 17868 9424
rect 17920 9415 17922 9424
rect 17868 9386 17920 9392
rect 17880 9178 17908 9386
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17880 8634 17908 8978
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17972 8498 18000 10678
rect 18064 10606 18092 10746
rect 18142 10704 18198 10713
rect 18142 10639 18198 10648
rect 18328 10668 18380 10674
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 18156 10470 18184 10639
rect 18328 10610 18380 10616
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18340 10266 18368 10610
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 18064 8809 18092 9998
rect 18050 8800 18106 8809
rect 18050 8735 18106 8744
rect 18616 8650 18644 12543
rect 18708 10810 18736 16934
rect 18800 16289 18828 21286
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 19076 19417 19104 20334
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 19062 19408 19118 19417
rect 19260 19378 19288 19858
rect 19062 19343 19118 19352
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19064 19304 19116 19310
rect 19062 19272 19064 19281
rect 19892 19304 19944 19310
rect 19116 19272 19118 19281
rect 19890 19272 19892 19281
rect 19944 19272 19946 19281
rect 19062 19207 19118 19216
rect 19340 19236 19392 19242
rect 19890 19207 19946 19216
rect 19340 19178 19392 19184
rect 19248 19168 19300 19174
rect 19246 19136 19248 19145
rect 19300 19136 19302 19145
rect 19246 19071 19302 19080
rect 19246 18320 19302 18329
rect 19246 18255 19248 18264
rect 19300 18255 19302 18264
rect 19248 18226 19300 18232
rect 19248 18080 19300 18086
rect 19352 18057 19380 19178
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19614 18728 19670 18737
rect 19614 18663 19670 18672
rect 19628 18222 19656 18663
rect 19628 18216 19703 18222
rect 19628 18176 19651 18216
rect 19651 18158 19703 18164
rect 19248 18022 19300 18028
rect 19338 18048 19394 18057
rect 19260 17513 19288 18022
rect 19338 17983 19394 17992
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19246 17504 19302 17513
rect 19246 17439 19302 17448
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18786 16280 18842 16289
rect 18786 16215 18842 16224
rect 18892 16153 18920 17070
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 18970 16824 19026 16833
rect 18970 16759 19026 16768
rect 18984 16658 19012 16759
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 18878 16144 18934 16153
rect 18878 16079 18934 16088
rect 18788 15972 18840 15978
rect 18788 15914 18840 15920
rect 18800 15638 18828 15914
rect 19076 15910 19104 16526
rect 19432 16176 19484 16182
rect 19432 16118 19484 16124
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 18788 15632 18840 15638
rect 18788 15574 18840 15580
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 18800 15026 18828 15574
rect 18892 15162 18920 15574
rect 19062 15328 19118 15337
rect 19062 15263 19118 15272
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18972 14544 19024 14550
rect 18972 14486 19024 14492
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18800 14006 18828 14350
rect 18984 14074 19012 14486
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18788 14000 18840 14006
rect 18788 13942 18840 13948
rect 18800 13326 18828 13942
rect 18880 13796 18932 13802
rect 18880 13738 18932 13744
rect 18788 13320 18840 13326
rect 18892 13297 18920 13738
rect 18788 13262 18840 13268
rect 18878 13288 18934 13297
rect 18878 13223 18934 13232
rect 18892 12918 18920 13223
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18984 12696 19012 14010
rect 19076 12866 19104 15263
rect 19260 14890 19288 15846
rect 19444 15638 19472 16118
rect 19536 16114 19564 16934
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19892 16720 19944 16726
rect 19892 16662 19944 16668
rect 19904 16114 19932 16662
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19536 15706 19564 16050
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19340 14816 19392 14822
rect 19338 14784 19340 14793
rect 19524 14816 19576 14822
rect 19392 14784 19394 14793
rect 19524 14758 19576 14764
rect 19338 14719 19394 14728
rect 19536 14550 19564 14758
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19524 14544 19576 14550
rect 19524 14486 19576 14492
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19260 13462 19288 14350
rect 19996 14226 20024 20198
rect 20076 18828 20128 18834
rect 20076 18770 20128 18776
rect 20088 18426 20116 18770
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20168 14544 20220 14550
rect 20168 14486 20220 14492
rect 19904 14198 20024 14226
rect 19904 13784 19932 14198
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19904 13756 20024 13784
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19248 13456 19300 13462
rect 19248 13398 19300 13404
rect 19798 13016 19854 13025
rect 19798 12951 19854 12960
rect 19076 12838 19196 12866
rect 18892 12668 19012 12696
rect 18892 12374 18920 12668
rect 19168 12628 19196 12838
rect 19812 12782 19840 12951
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 18984 12600 19196 12628
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18892 11898 18920 12310
rect 18984 12209 19012 12600
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19616 12368 19668 12374
rect 19522 12336 19578 12345
rect 19616 12310 19668 12316
rect 19522 12271 19578 12280
rect 19340 12232 19392 12238
rect 18970 12200 19026 12209
rect 18970 12135 19026 12144
rect 19338 12200 19340 12209
rect 19392 12200 19394 12209
rect 19338 12135 19394 12144
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 18880 11892 18932 11898
rect 18932 11852 19012 11880
rect 18880 11834 18932 11840
rect 18880 11688 18932 11694
rect 18878 11656 18880 11665
rect 18932 11656 18934 11665
rect 18984 11626 19012 11852
rect 18878 11591 18934 11600
rect 18972 11620 19024 11626
rect 18892 11354 18920 11591
rect 18972 11562 19024 11568
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18892 9761 18920 10066
rect 18878 9752 18934 9761
rect 18878 9687 18934 9696
rect 18892 9382 18920 9687
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18694 8664 18750 8673
rect 18616 8622 18694 8650
rect 18694 8599 18750 8608
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 18326 8256 18382 8265
rect 18326 8191 18382 8200
rect 18340 7954 18368 8191
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 18340 7546 18368 7890
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17880 6934 17908 7142
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17880 6118 17908 6870
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18156 6254 18184 6598
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17880 5574 17908 6054
rect 18432 5914 18460 6734
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17880 3942 17908 5510
rect 18050 5400 18106 5409
rect 18050 5335 18106 5344
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17880 2582 17908 3878
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 18064 610 18092 5335
rect 18328 5092 18380 5098
rect 18328 5034 18380 5040
rect 18420 5092 18472 5098
rect 18420 5034 18472 5040
rect 18340 5001 18368 5034
rect 18326 4992 18382 5001
rect 18248 4950 18326 4978
rect 18248 4826 18276 4950
rect 18326 4927 18382 4936
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18340 4622 18368 4762
rect 18432 4758 18460 5034
rect 18420 4752 18472 4758
rect 18420 4694 18472 4700
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 18432 4282 18460 4694
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18156 3398 18184 4014
rect 18420 3664 18472 3670
rect 18420 3606 18472 3612
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18144 3392 18196 3398
rect 18340 3369 18368 3470
rect 18144 3334 18196 3340
rect 18326 3360 18382 3369
rect 18156 2553 18184 3334
rect 18326 3295 18382 3304
rect 18432 2922 18460 3606
rect 18708 2938 18736 8599
rect 18892 7857 18920 9318
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 18984 8498 19012 9046
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18878 7848 18934 7857
rect 18878 7783 18934 7792
rect 19076 7274 19104 9454
rect 19168 8906 19196 12038
rect 19352 11286 19380 12135
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19352 10470 19380 11086
rect 19444 10538 19472 11154
rect 19432 10532 19484 10538
rect 19432 10474 19484 10480
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9586 19288 9862
rect 19352 9722 19380 10406
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19156 8900 19208 8906
rect 19156 8842 19208 8848
rect 19260 8634 19288 9522
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19352 8838 19380 9386
rect 19444 9042 19472 9998
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19352 8362 19380 8774
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19352 8090 19380 8298
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19444 7698 19472 8842
rect 19352 7670 19472 7698
rect 19156 7472 19208 7478
rect 19156 7414 19208 7420
rect 18788 7268 18840 7274
rect 18788 7210 18840 7216
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 18800 7002 18828 7210
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18970 6216 19026 6225
rect 18970 6151 19026 6160
rect 18984 5846 19012 6151
rect 18972 5840 19024 5846
rect 18972 5782 19024 5788
rect 19168 5642 19196 7414
rect 19352 6338 19380 7670
rect 19536 7562 19564 12271
rect 19628 11830 19656 12310
rect 19616 11824 19668 11830
rect 19616 11766 19668 11772
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19798 8800 19854 8809
rect 19798 8735 19854 8744
rect 19812 8566 19840 8735
rect 19800 8560 19852 8566
rect 19800 8502 19852 8508
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19444 7534 19564 7562
rect 19444 6866 19472 7534
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19536 7002 19564 7346
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19444 6458 19472 6802
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19352 6310 19472 6338
rect 19338 6216 19394 6225
rect 19338 6151 19394 6160
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19260 5846 19288 6054
rect 19248 5840 19300 5846
rect 19248 5782 19300 5788
rect 19156 5636 19208 5642
rect 19156 5578 19208 5584
rect 19260 5370 19288 5782
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 19352 5302 19380 6151
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19248 5160 19300 5166
rect 19248 5102 19300 5108
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 18984 3670 19012 4558
rect 19260 4146 19288 5102
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19352 4185 19380 4422
rect 19338 4176 19394 4185
rect 19248 4140 19300 4146
rect 19338 4111 19394 4120
rect 19248 4082 19300 4088
rect 19444 4049 19472 6310
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5636 19576 5642
rect 19524 5578 19576 5584
rect 19430 4040 19486 4049
rect 19430 3975 19486 3984
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18800 3058 18828 3470
rect 18984 3058 19012 3606
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18420 2916 18472 2922
rect 18708 2910 18828 2938
rect 19260 2922 19288 3878
rect 19536 3074 19564 5578
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19708 4684 19760 4690
rect 19708 4626 19760 4632
rect 19720 4457 19748 4626
rect 19706 4448 19762 4457
rect 19706 4383 19762 4392
rect 19720 4282 19748 4383
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 19996 4162 20024 13756
rect 20088 13530 20116 13874
rect 20180 13802 20208 14486
rect 20168 13796 20220 13802
rect 20168 13738 20220 13744
rect 20166 13560 20222 13569
rect 20076 13524 20128 13530
rect 20166 13495 20222 13504
rect 20076 13466 20128 13472
rect 20180 13462 20208 13495
rect 20168 13456 20220 13462
rect 20168 13398 20220 13404
rect 20272 12102 20300 18022
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20166 11112 20222 11121
rect 20166 11047 20222 11056
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 20088 9353 20116 9386
rect 20074 9344 20130 9353
rect 20074 9279 20130 9288
rect 20074 8120 20130 8129
rect 20074 8055 20130 8064
rect 20088 7721 20116 8055
rect 20074 7712 20130 7721
rect 20074 7647 20130 7656
rect 20180 7206 20208 11047
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20272 9722 20300 10066
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20272 8634 20300 9318
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20258 7712 20314 7721
rect 20258 7647 20314 7656
rect 20272 7342 20300 7647
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20272 7002 20300 7278
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20258 6760 20314 6769
rect 20258 6695 20314 6704
rect 20272 6497 20300 6695
rect 20074 6488 20130 6497
rect 20074 6423 20130 6432
rect 20258 6488 20314 6497
rect 20258 6423 20314 6432
rect 20088 6089 20116 6423
rect 20166 6352 20222 6361
rect 20166 6287 20222 6296
rect 20180 6254 20208 6287
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 20074 6080 20130 6089
rect 20074 6015 20130 6024
rect 20180 5914 20208 6190
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20168 4208 20220 4214
rect 19996 4146 20116 4162
rect 20168 4150 20220 4156
rect 19984 4140 20116 4146
rect 20036 4134 20116 4140
rect 19984 4082 20036 4088
rect 19982 4040 20038 4049
rect 19982 3975 20038 3984
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19996 3738 20024 3975
rect 20088 3738 20116 4134
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 20180 3641 20208 4150
rect 20166 3632 20222 3641
rect 20166 3567 20168 3576
rect 20220 3567 20222 3576
rect 20168 3538 20220 3544
rect 20180 3194 20208 3538
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 19536 3046 20024 3074
rect 18420 2858 18472 2864
rect 18432 2650 18460 2858
rect 18420 2644 18472 2650
rect 18420 2586 18472 2592
rect 18142 2544 18198 2553
rect 18142 2479 18198 2488
rect 18328 2440 18380 2446
rect 18326 2408 18328 2417
rect 18380 2408 18382 2417
rect 18326 2343 18382 2352
rect 18052 604 18104 610
rect 18052 546 18104 552
rect 18800 480 18828 2910
rect 19248 2916 19300 2922
rect 19248 2858 19300 2864
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19996 2514 20024 3046
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 20272 2106 20300 4966
rect 20364 4826 20392 18566
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20640 16425 20668 18022
rect 20810 17776 20866 17785
rect 20810 17711 20812 17720
rect 20864 17711 20866 17720
rect 20812 17682 20864 17688
rect 20824 17338 20852 17682
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20718 17232 20774 17241
rect 20718 17167 20774 17176
rect 20732 17134 20760 17167
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20810 16960 20866 16969
rect 20732 16697 20760 16934
rect 20810 16895 20866 16904
rect 20718 16688 20774 16697
rect 20718 16623 20774 16632
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20626 16416 20682 16425
rect 20626 16351 20682 16360
rect 20732 16250 20760 16458
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20548 14618 20576 14894
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20732 13954 20760 15914
rect 20640 13938 20760 13954
rect 20628 13932 20760 13938
rect 20680 13926 20760 13932
rect 20628 13874 20680 13880
rect 20720 13252 20772 13258
rect 20720 13194 20772 13200
rect 20442 13152 20498 13161
rect 20732 13138 20760 13194
rect 20442 13087 20498 13096
rect 20548 13110 20760 13138
rect 20456 11014 20484 13087
rect 20548 12374 20576 13110
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20536 12368 20588 12374
rect 20536 12310 20588 12316
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20548 11626 20576 12106
rect 20536 11620 20588 11626
rect 20536 11562 20588 11568
rect 20640 11286 20668 12786
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20732 11762 20760 12038
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20824 11642 20852 16895
rect 20732 11614 20852 11642
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20444 11008 20496 11014
rect 20444 10950 20496 10956
rect 20444 10464 20496 10470
rect 20548 10452 20576 11154
rect 20628 10532 20680 10538
rect 20628 10474 20680 10480
rect 20496 10424 20576 10452
rect 20444 10406 20496 10412
rect 20456 8129 20484 10406
rect 20640 9926 20668 10474
rect 20732 9926 20760 11614
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20534 9480 20590 9489
rect 20534 9415 20590 9424
rect 20548 8673 20576 9415
rect 20534 8664 20590 8673
rect 20534 8599 20590 8608
rect 20640 8514 20668 9862
rect 20718 9616 20774 9625
rect 20718 9551 20774 9560
rect 20732 8634 20760 9551
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20548 8486 20668 8514
rect 20442 8120 20498 8129
rect 20442 8055 20498 8064
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20456 5846 20484 6190
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 20548 5778 20576 8486
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20626 7848 20682 7857
rect 20626 7783 20682 7792
rect 20640 7342 20668 7783
rect 20732 7449 20760 8366
rect 20718 7440 20774 7449
rect 20718 7375 20774 7384
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20720 6180 20772 6186
rect 20720 6122 20772 6128
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20628 4684 20680 4690
rect 20732 4672 20760 6122
rect 20680 4644 20760 4672
rect 20628 4626 20680 4632
rect 20536 4004 20588 4010
rect 20536 3946 20588 3952
rect 20548 3913 20576 3946
rect 20534 3904 20590 3913
rect 20534 3839 20590 3848
rect 20824 3602 20852 11494
rect 20916 6225 20944 18702
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21088 16652 21140 16658
rect 21088 16594 21140 16600
rect 21100 16114 21128 16594
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 21192 15638 21220 18022
rect 21284 16794 21312 23462
rect 21638 18728 21694 18737
rect 21638 18663 21694 18672
rect 21364 17536 21416 17542
rect 21364 17478 21416 17484
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 21180 15632 21232 15638
rect 21180 15574 21232 15580
rect 21192 15162 21220 15574
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 21376 14940 21404 17478
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21456 15632 21508 15638
rect 21456 15574 21508 15580
rect 21468 14958 21496 15574
rect 21284 14912 21404 14940
rect 21456 14952 21508 14958
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21008 14414 21036 14758
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 21008 13530 21036 14350
rect 21100 14074 21128 14486
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21100 12850 21128 13126
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21180 12708 21232 12714
rect 21180 12650 21232 12656
rect 21192 12374 21220 12650
rect 21180 12368 21232 12374
rect 21180 12310 21232 12316
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 21008 11762 21036 12174
rect 21192 12170 21220 12310
rect 21180 12164 21232 12170
rect 21180 12106 21232 12112
rect 21284 12050 21312 14912
rect 21456 14894 21508 14900
rect 21560 14770 21588 16934
rect 21652 14958 21680 18663
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 21732 16108 21784 16114
rect 21732 16050 21784 16056
rect 21744 15434 21772 16050
rect 21824 15904 21876 15910
rect 21824 15846 21876 15852
rect 21732 15428 21784 15434
rect 21732 15370 21784 15376
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 21192 12022 21312 12050
rect 21376 14742 21588 14770
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 21008 11354 21036 11698
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 21008 10606 21036 10950
rect 21192 10674 21220 12022
rect 21270 11928 21326 11937
rect 21270 11863 21326 11872
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 20996 10600 21048 10606
rect 20996 10542 21048 10548
rect 21008 9722 21036 10542
rect 21180 10532 21232 10538
rect 21180 10474 21232 10480
rect 21086 10432 21142 10441
rect 21086 10367 21142 10376
rect 21100 10266 21128 10367
rect 21192 10266 21220 10474
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 21180 10260 21232 10266
rect 21180 10202 21232 10208
rect 21088 9920 21140 9926
rect 21088 9862 21140 9868
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 20902 6216 20958 6225
rect 21008 6186 21036 9046
rect 21100 6202 21128 9862
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21192 8498 21220 8774
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 21180 7200 21232 7206
rect 21178 7168 21180 7177
rect 21232 7168 21234 7177
rect 21178 7103 21234 7112
rect 20902 6151 20958 6160
rect 20996 6180 21048 6186
rect 21100 6174 21220 6202
rect 20996 6122 21048 6128
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 21008 5817 21036 5850
rect 20994 5808 21050 5817
rect 20904 5772 20956 5778
rect 20994 5743 21050 5752
rect 20904 5714 20956 5720
rect 20916 5273 20944 5714
rect 20902 5264 20958 5273
rect 20902 5199 20958 5208
rect 21100 5030 21128 6054
rect 21192 5137 21220 6174
rect 21284 5370 21312 11863
rect 21376 11558 21404 14742
rect 21652 14634 21680 14894
rect 21560 14606 21680 14634
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21468 13326 21496 14350
rect 21560 13682 21588 14606
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21652 13802 21680 14214
rect 21744 13938 21772 15370
rect 21732 13932 21784 13938
rect 21732 13874 21784 13880
rect 21640 13796 21692 13802
rect 21640 13738 21692 13744
rect 21560 13654 21680 13682
rect 21548 13456 21600 13462
rect 21548 13398 21600 13404
rect 21456 13320 21508 13326
rect 21454 13288 21456 13297
rect 21508 13288 21510 13297
rect 21454 13223 21510 13232
rect 21560 12986 21588 13398
rect 21652 13138 21680 13654
rect 21744 13258 21772 13874
rect 21732 13252 21784 13258
rect 21732 13194 21784 13200
rect 21652 13110 21772 13138
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21376 5930 21404 10610
rect 21468 10130 21496 12786
rect 21560 11898 21588 12922
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21560 10810 21588 11018
rect 21744 10962 21772 13110
rect 21652 10934 21772 10962
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21652 10248 21680 10934
rect 21836 10826 21864 15846
rect 21928 11082 21956 18226
rect 22204 17649 22232 23598
rect 24596 23225 24624 23598
rect 24688 23322 24716 24511
rect 24780 23866 24808 25871
rect 25792 24313 25820 27520
rect 25778 24304 25834 24313
rect 25778 24239 25834 24248
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 27172 23497 27200 27520
rect 24766 23488 24822 23497
rect 24766 23423 24822 23432
rect 27158 23488 27214 23497
rect 27158 23423 27214 23432
rect 24676 23316 24728 23322
rect 24676 23258 24728 23264
rect 23386 23216 23442 23225
rect 24582 23216 24638 23225
rect 23386 23151 23442 23160
rect 24124 23180 24176 23186
rect 23400 17898 23428 23151
rect 24780 23202 24808 23423
rect 24582 23151 24638 23160
rect 24688 23174 24808 23202
rect 24124 23122 24176 23128
rect 23754 22536 23810 22545
rect 23754 22471 23810 22480
rect 23662 21584 23718 21593
rect 23662 21519 23718 21528
rect 23216 17870 23428 17898
rect 22836 17740 22888 17746
rect 22836 17682 22888 17688
rect 22190 17640 22246 17649
rect 22190 17575 22246 17584
rect 22006 17504 22062 17513
rect 22006 17439 22062 17448
rect 22020 12850 22048 17439
rect 22204 17134 22232 17575
rect 22376 17536 22428 17542
rect 22376 17478 22428 17484
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22284 16584 22336 16590
rect 22284 16526 22336 16532
rect 22098 16280 22154 16289
rect 22098 16215 22154 16224
rect 22112 15978 22140 16215
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22204 15609 22232 15846
rect 22190 15600 22246 15609
rect 22190 15535 22246 15544
rect 22296 15502 22324 16526
rect 22100 15496 22152 15502
rect 22098 15464 22100 15473
rect 22284 15496 22336 15502
rect 22152 15464 22154 15473
rect 22284 15438 22336 15444
rect 22098 15399 22154 15408
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22296 14006 22324 14214
rect 22284 14000 22336 14006
rect 22284 13942 22336 13948
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22100 13252 22152 13258
rect 22100 13194 22152 13200
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22008 12708 22060 12714
rect 22008 12650 22060 12656
rect 22020 12442 22048 12650
rect 22008 12436 22060 12442
rect 22008 12378 22060 12384
rect 22112 12306 22140 13194
rect 22204 12714 22232 13738
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22296 12646 22324 12854
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22100 12096 22152 12102
rect 22204 12073 22232 12378
rect 22296 12374 22324 12582
rect 22284 12368 22336 12374
rect 22284 12310 22336 12316
rect 22282 12200 22338 12209
rect 22282 12135 22338 12144
rect 22100 12038 22152 12044
rect 22190 12064 22246 12073
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 21836 10798 21956 10826
rect 21824 10260 21876 10266
rect 21652 10220 21772 10248
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21456 9988 21508 9994
rect 21456 9930 21508 9936
rect 21468 7449 21496 9930
rect 21652 9450 21680 10066
rect 21640 9444 21692 9450
rect 21640 9386 21692 9392
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21560 8537 21588 9318
rect 21546 8528 21602 8537
rect 21546 8463 21602 8472
rect 21454 7440 21510 7449
rect 21454 7375 21510 7384
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21560 6254 21588 6598
rect 21548 6248 21600 6254
rect 21546 6216 21548 6225
rect 21600 6216 21602 6225
rect 21546 6151 21602 6160
rect 21376 5902 21496 5930
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 21178 5128 21234 5137
rect 21178 5063 21234 5072
rect 21088 5024 21140 5030
rect 21088 4966 21140 4972
rect 21100 4758 21128 4966
rect 21088 4752 21140 4758
rect 21088 4694 21140 4700
rect 21100 3942 21128 4694
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20810 3496 20866 3505
rect 20810 3431 20866 3440
rect 20824 3058 20852 3431
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 21100 2922 21128 3878
rect 21192 3777 21220 4558
rect 21376 4554 21404 5714
rect 21364 4548 21416 4554
rect 21364 4490 21416 4496
rect 21468 4162 21496 5902
rect 21376 4134 21496 4162
rect 21178 3768 21234 3777
rect 21178 3703 21180 3712
rect 21232 3703 21234 3712
rect 21180 3674 21232 3680
rect 21376 3369 21404 4134
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 21468 3670 21496 3946
rect 21456 3664 21508 3670
rect 21456 3606 21508 3612
rect 21362 3360 21418 3369
rect 21362 3295 21418 3304
rect 21088 2916 21140 2922
rect 21088 2858 21140 2864
rect 20626 2680 20682 2689
rect 20626 2615 20628 2624
rect 20680 2615 20682 2624
rect 20628 2586 20680 2592
rect 21468 2446 21496 3606
rect 21456 2440 21508 2446
rect 21652 2394 21680 9386
rect 21744 9110 21772 10220
rect 21824 10202 21876 10208
rect 21836 9586 21864 10202
rect 21928 10169 21956 10798
rect 22020 10198 22048 11494
rect 22112 10470 22140 12038
rect 22190 11999 22246 12008
rect 22204 11393 22232 11999
rect 22296 11898 22324 12135
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22190 11384 22246 11393
rect 22190 11319 22246 11328
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22296 10606 22324 10950
rect 22284 10600 22336 10606
rect 22284 10542 22336 10548
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22008 10192 22060 10198
rect 21914 10160 21970 10169
rect 22008 10134 22060 10140
rect 22100 10192 22152 10198
rect 22100 10134 22152 10140
rect 21914 10095 21970 10104
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21744 7818 21772 8910
rect 21836 8786 21864 9046
rect 21928 8906 21956 9998
rect 22008 9716 22060 9722
rect 22008 9658 22060 9664
rect 21916 8900 21968 8906
rect 21916 8842 21968 8848
rect 21836 8758 21956 8786
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21836 8265 21864 8434
rect 21928 8294 21956 8758
rect 22020 8650 22048 9658
rect 22112 9432 22140 10134
rect 22192 9444 22244 9450
rect 22112 9404 22192 9432
rect 22112 9110 22140 9404
rect 22192 9386 22244 9392
rect 22100 9104 22152 9110
rect 22100 9046 22152 9052
rect 22020 8634 22140 8650
rect 22020 8628 22152 8634
rect 22020 8622 22100 8628
rect 22100 8570 22152 8576
rect 21916 8288 21968 8294
rect 21822 8256 21878 8265
rect 21916 8230 21968 8236
rect 21822 8191 21878 8200
rect 21928 8022 21956 8230
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21732 7812 21784 7818
rect 21732 7754 21784 7760
rect 21744 7206 21772 7754
rect 21824 7744 21876 7750
rect 21928 7732 21956 7958
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 21876 7704 21956 7732
rect 21824 7686 21876 7692
rect 21836 7410 21864 7686
rect 21914 7440 21970 7449
rect 21824 7404 21876 7410
rect 21914 7375 21970 7384
rect 21824 7346 21876 7352
rect 21732 7200 21784 7206
rect 21732 7142 21784 7148
rect 21836 6934 21864 7346
rect 21824 6928 21876 6934
rect 21824 6870 21876 6876
rect 21836 6186 21864 6870
rect 21824 6180 21876 6186
rect 21824 6122 21876 6128
rect 21928 6066 21956 7375
rect 22020 6662 22048 7822
rect 22296 7177 22324 10542
rect 22282 7168 22338 7177
rect 22282 7103 22338 7112
rect 22388 6916 22416 17478
rect 22480 16969 22508 17478
rect 22848 16998 22876 17682
rect 22836 16992 22888 16998
rect 22466 16960 22522 16969
rect 22836 16934 22888 16940
rect 22466 16895 22522 16904
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22560 15972 22612 15978
rect 22560 15914 22612 15920
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22480 14521 22508 15302
rect 22466 14512 22522 14521
rect 22466 14447 22522 14456
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22480 12986 22508 13262
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22480 12442 22508 12786
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22466 12336 22522 12345
rect 22466 12271 22522 12280
rect 22480 11694 22508 12271
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 22466 11384 22522 11393
rect 22466 11319 22522 11328
rect 22204 6888 22416 6916
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 21836 6038 21956 6066
rect 21836 5409 21864 6038
rect 21916 5568 21968 5574
rect 21916 5510 21968 5516
rect 21822 5400 21878 5409
rect 21822 5335 21878 5344
rect 21928 5273 21956 5510
rect 21914 5264 21970 5273
rect 21914 5199 21916 5208
rect 21968 5199 21970 5208
rect 21916 5170 21968 5176
rect 21928 5139 21956 5170
rect 22204 5114 22232 6888
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 22388 5574 22416 6734
rect 22480 6361 22508 11319
rect 22572 9994 22600 15914
rect 22560 9988 22612 9994
rect 22560 9930 22612 9936
rect 22466 6352 22522 6361
rect 22466 6287 22522 6296
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 22480 5846 22508 6054
rect 22468 5840 22520 5846
rect 22468 5782 22520 5788
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22020 5086 22232 5114
rect 22374 5128 22430 5137
rect 22020 4570 22048 5086
rect 22374 5063 22376 5072
rect 22428 5063 22430 5072
rect 22376 5034 22428 5040
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 22112 4758 22140 4966
rect 22480 4826 22508 5782
rect 22664 5710 22692 16526
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 22756 13870 22784 14418
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22756 12850 22784 13806
rect 22848 13682 22876 16934
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 23112 16652 23164 16658
rect 23112 16594 23164 16600
rect 22940 16046 22968 16594
rect 22928 16040 22980 16046
rect 22926 16008 22928 16017
rect 22980 16008 22982 16017
rect 22926 15943 22982 15952
rect 22940 15570 22968 15943
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 22940 15162 22968 15506
rect 22928 15156 22980 15162
rect 22928 15098 22980 15104
rect 22928 14476 22980 14482
rect 22928 14418 22980 14424
rect 22940 13802 22968 14418
rect 23020 14000 23072 14006
rect 23020 13942 23072 13948
rect 22928 13796 22980 13802
rect 22928 13738 22980 13744
rect 22848 13654 22968 13682
rect 22834 13424 22890 13433
rect 22834 13359 22890 13368
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22756 12238 22784 12582
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22756 11354 22784 12174
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 22848 10577 22876 13359
rect 22834 10568 22890 10577
rect 22834 10503 22890 10512
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22756 9722 22784 10406
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 22836 8628 22888 8634
rect 22836 8570 22888 8576
rect 22848 7546 22876 8570
rect 22836 7540 22888 7546
rect 22836 7482 22888 7488
rect 22848 7342 22876 7482
rect 22836 7336 22888 7342
rect 22836 7278 22888 7284
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22664 5370 22692 5646
rect 22652 5364 22704 5370
rect 22652 5306 22704 5312
rect 22468 4820 22520 4826
rect 22468 4762 22520 4768
rect 22100 4752 22152 4758
rect 22100 4694 22152 4700
rect 22652 4752 22704 4758
rect 22652 4694 22704 4700
rect 21928 4542 22048 4570
rect 22192 4548 22244 4554
rect 21732 3664 21784 3670
rect 21732 3606 21784 3612
rect 21744 2854 21772 3606
rect 21928 3534 21956 4542
rect 22192 4490 22244 4496
rect 22008 4480 22060 4486
rect 22008 4422 22060 4428
rect 22020 4282 22048 4422
rect 22008 4276 22060 4282
rect 22008 4218 22060 4224
rect 22020 4026 22048 4218
rect 22020 4010 22140 4026
rect 22020 4004 22152 4010
rect 22020 3998 22100 4004
rect 22100 3946 22152 3952
rect 22204 3670 22232 4490
rect 22664 3738 22692 4694
rect 22652 3732 22704 3738
rect 22652 3674 22704 3680
rect 22192 3664 22244 3670
rect 22192 3606 22244 3612
rect 22756 3602 22784 6938
rect 22848 6458 22876 7278
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 22836 4072 22888 4078
rect 22834 4040 22836 4049
rect 22888 4040 22890 4049
rect 22834 3975 22890 3984
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 21744 2582 21772 2790
rect 21928 2650 21956 3470
rect 22374 3224 22430 3233
rect 22374 3159 22376 3168
rect 22428 3159 22430 3168
rect 22376 3130 22428 3136
rect 22756 3058 22784 3538
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 21732 2576 21784 2582
rect 21732 2518 21784 2524
rect 21456 2382 21508 2388
rect 21560 2366 21680 2394
rect 22756 2378 22784 2994
rect 22744 2372 22796 2378
rect 21560 2145 21588 2366
rect 22744 2314 22796 2320
rect 21640 2304 21692 2310
rect 21640 2246 21692 2252
rect 21546 2136 21602 2145
rect 20260 2100 20312 2106
rect 21546 2071 21602 2080
rect 20260 2042 20312 2048
rect 19706 2000 19762 2009
rect 19706 1935 19762 1944
rect 19720 480 19748 1935
rect 20718 1728 20774 1737
rect 20718 1663 20774 1672
rect 20732 480 20760 1663
rect 21652 480 21680 2246
rect 22652 2100 22704 2106
rect 22652 2042 22704 2048
rect 22664 480 22692 2042
rect 22940 785 22968 13654
rect 23032 12238 23060 13942
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23032 9761 23060 12038
rect 23018 9752 23074 9761
rect 23018 9687 23074 9696
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 23032 9353 23060 9522
rect 23018 9344 23074 9353
rect 23018 9279 23074 9288
rect 23032 9110 23060 9279
rect 23020 9104 23072 9110
rect 23020 9046 23072 9052
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 23032 3913 23060 4558
rect 23018 3904 23074 3913
rect 23018 3839 23074 3848
rect 23032 3534 23060 3839
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23124 2650 23152 16594
rect 23216 13433 23244 17870
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 23400 16998 23428 17682
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23400 14929 23428 16934
rect 23480 15360 23532 15366
rect 23478 15328 23480 15337
rect 23532 15328 23534 15337
rect 23478 15263 23534 15272
rect 23386 14920 23442 14929
rect 23386 14855 23442 14864
rect 23572 14884 23624 14890
rect 23572 14826 23624 14832
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23492 13841 23520 14758
rect 23478 13832 23534 13841
rect 23478 13767 23534 13776
rect 23480 13728 23532 13734
rect 23480 13670 23532 13676
rect 23492 13569 23520 13670
rect 23478 13560 23534 13569
rect 23478 13495 23534 13504
rect 23388 13456 23440 13462
rect 23202 13424 23258 13433
rect 23388 13398 23440 13404
rect 23202 13359 23258 13368
rect 23400 12986 23428 13398
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23296 12640 23348 12646
rect 23296 12582 23348 12588
rect 23204 12368 23256 12374
rect 23204 12310 23256 12316
rect 23216 11830 23244 12310
rect 23204 11824 23256 11830
rect 23204 11766 23256 11772
rect 23308 11744 23336 12582
rect 23308 11716 23428 11744
rect 23296 11620 23348 11626
rect 23296 11562 23348 11568
rect 23204 11552 23256 11558
rect 23204 11494 23256 11500
rect 23216 11354 23244 11494
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23216 10538 23244 11290
rect 23204 10532 23256 10538
rect 23204 10474 23256 10480
rect 23308 10146 23336 11562
rect 23400 11286 23428 11716
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23400 10266 23428 11222
rect 23492 10470 23520 11222
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23388 10260 23440 10266
rect 23388 10202 23440 10208
rect 23308 10118 23520 10146
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23216 8838 23244 9998
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 23294 9752 23350 9761
rect 23294 9687 23350 9696
rect 23204 8832 23256 8838
rect 23202 8800 23204 8809
rect 23256 8800 23258 8809
rect 23202 8735 23258 8744
rect 23308 7002 23336 9687
rect 23400 7342 23428 9862
rect 23492 7721 23520 10118
rect 23584 9110 23612 14826
rect 23676 12617 23704 21519
rect 23768 15570 23796 22471
rect 24136 22438 24164 23122
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24124 22432 24176 22438
rect 24124 22374 24176 22380
rect 24136 20505 24164 22374
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24122 20496 24178 20505
rect 24122 20431 24178 20440
rect 24136 19417 24164 20431
rect 24122 19408 24178 19417
rect 24122 19343 24178 19352
rect 24122 17504 24178 17513
rect 24122 17439 24178 17448
rect 24136 17134 24164 17439
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 24228 15570 24256 21286
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24584 19304 24636 19310
rect 24584 19246 24636 19252
rect 24596 18737 24624 19246
rect 24688 18970 24716 23174
rect 24766 23080 24822 23089
rect 24766 23015 24822 23024
rect 24780 21690 24808 23015
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24766 20360 24822 20369
rect 24766 20295 24822 20304
rect 24780 19514 24808 20295
rect 24768 19508 24820 19514
rect 24768 19450 24820 19456
rect 25778 19408 25834 19417
rect 25778 19343 25834 19352
rect 24676 18964 24728 18970
rect 24676 18906 24728 18912
rect 24766 18864 24822 18873
rect 24676 18828 24728 18834
rect 24766 18799 24822 18808
rect 24676 18770 24728 18776
rect 24582 18728 24638 18737
rect 24582 18663 24638 18672
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24584 18352 24636 18358
rect 24582 18320 24584 18329
rect 24636 18320 24638 18329
rect 24688 18306 24716 18770
rect 24638 18278 24716 18306
rect 24582 18255 24638 18264
rect 24674 17504 24730 17513
rect 24289 17436 24585 17456
rect 24674 17439 24730 17448
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 16810 24716 17439
rect 24780 17338 24808 18799
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 25044 17060 25096 17066
rect 25044 17002 25096 17008
rect 24688 16782 24808 16810
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 24216 15564 24268 15570
rect 24216 15506 24268 15512
rect 23952 14822 23980 15506
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24032 14952 24084 14958
rect 24032 14894 24084 14900
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23768 13870 23796 14214
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23662 12608 23718 12617
rect 23662 12543 23718 12552
rect 23768 12238 23796 13806
rect 23848 13796 23900 13802
rect 23848 13738 23900 13744
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 23664 12096 23716 12102
rect 23664 12038 23716 12044
rect 23676 11694 23704 12038
rect 23860 11694 23888 13738
rect 23952 12084 23980 14758
rect 24044 13705 24072 14894
rect 24688 14482 24716 16662
rect 24780 16250 24808 16782
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24766 16144 24822 16153
rect 24766 16079 24822 16088
rect 24780 14618 24808 16079
rect 24858 15056 24914 15065
rect 24858 14991 24914 15000
rect 24768 14612 24820 14618
rect 24768 14554 24820 14560
rect 24766 14512 24822 14521
rect 24676 14476 24728 14482
rect 24766 14447 24822 14456
rect 24676 14418 24728 14424
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 14074 24716 14418
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24030 13696 24086 13705
rect 24030 13631 24086 13640
rect 24030 13560 24086 13569
rect 24030 13495 24086 13504
rect 24044 13161 24072 13495
rect 24214 13424 24270 13433
rect 24214 13359 24216 13368
rect 24268 13359 24270 13368
rect 24216 13330 24268 13336
rect 24030 13152 24086 13161
rect 24030 13087 24086 13096
rect 24228 12918 24256 13330
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24780 12986 24808 14447
rect 24872 14074 24900 14991
rect 24950 14920 25006 14929
rect 24950 14855 25006 14864
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24964 13870 24992 14855
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24216 12912 24268 12918
rect 24216 12854 24268 12860
rect 24766 12880 24822 12889
rect 24766 12815 24822 12824
rect 24860 12844 24912 12850
rect 24030 12608 24086 12617
rect 24030 12543 24086 12552
rect 24044 12209 24072 12543
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24030 12200 24086 12209
rect 24030 12135 24086 12144
rect 23952 12056 24072 12084
rect 23664 11688 23716 11694
rect 23848 11688 23900 11694
rect 23664 11630 23716 11636
rect 23754 11656 23810 11665
rect 23676 11234 23704 11630
rect 23848 11630 23900 11636
rect 23754 11591 23810 11600
rect 23768 11558 23796 11591
rect 23756 11552 23808 11558
rect 23756 11494 23808 11500
rect 23860 11354 23888 11630
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23676 11206 23796 11234
rect 23768 11200 23796 11206
rect 23768 11172 23980 11200
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23676 9994 23704 11086
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23756 11008 23808 11014
rect 23756 10950 23808 10956
rect 23768 10538 23796 10950
rect 23756 10532 23808 10538
rect 23756 10474 23808 10480
rect 23768 10441 23796 10474
rect 23754 10432 23810 10441
rect 23754 10367 23810 10376
rect 23860 10282 23888 11018
rect 23768 10254 23888 10282
rect 23664 9988 23716 9994
rect 23664 9930 23716 9936
rect 23572 9104 23624 9110
rect 23572 9046 23624 9052
rect 23584 8498 23612 9046
rect 23664 9036 23716 9042
rect 23664 8978 23716 8984
rect 23676 8566 23704 8978
rect 23664 8560 23716 8566
rect 23664 8502 23716 8508
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23768 8378 23796 10254
rect 23952 10180 23980 11172
rect 23860 10152 23980 10180
rect 23860 9926 23888 10152
rect 24044 10062 24072 12056
rect 24032 10056 24084 10062
rect 24136 10033 24164 12378
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24596 12186 24624 12242
rect 24596 12158 24716 12186
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11626 24716 12158
rect 24676 11620 24728 11626
rect 24676 11562 24728 11568
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24308 10464 24360 10470
rect 24308 10406 24360 10412
rect 24216 10192 24268 10198
rect 24216 10134 24268 10140
rect 24032 9998 24084 10004
rect 24122 10024 24178 10033
rect 23940 9988 23992 9994
rect 24122 9959 24178 9968
rect 23940 9930 23992 9936
rect 23848 9920 23900 9926
rect 23848 9862 23900 9868
rect 23848 9444 23900 9450
rect 23848 9386 23900 9392
rect 23860 9178 23888 9386
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23860 8634 23888 8978
rect 23848 8628 23900 8634
rect 23848 8570 23900 8576
rect 23584 8350 23796 8378
rect 23848 8356 23900 8362
rect 23478 7712 23534 7721
rect 23478 7647 23534 7656
rect 23388 7336 23440 7342
rect 23388 7278 23440 7284
rect 23400 7206 23428 7278
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 23478 7168 23534 7177
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 23400 6633 23428 7142
rect 23478 7103 23534 7112
rect 23386 6624 23442 6633
rect 23308 6582 23386 6610
rect 23202 5672 23258 5681
rect 23202 5607 23258 5616
rect 23216 3194 23244 5607
rect 23308 5370 23336 6582
rect 23386 6559 23442 6568
rect 23388 6384 23440 6390
rect 23386 6352 23388 6361
rect 23440 6352 23442 6361
rect 23386 6287 23442 6296
rect 23400 6254 23428 6287
rect 23388 6248 23440 6254
rect 23388 6190 23440 6196
rect 23492 5914 23520 7103
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23388 5568 23440 5574
rect 23440 5516 23520 5522
rect 23388 5510 23520 5516
rect 23400 5494 23520 5510
rect 23296 5364 23348 5370
rect 23296 5306 23348 5312
rect 23492 5030 23520 5494
rect 23480 5024 23532 5030
rect 23584 5001 23612 8350
rect 23848 8298 23900 8304
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 23754 8256 23810 8265
rect 23676 8022 23704 8230
rect 23754 8191 23810 8200
rect 23664 8016 23716 8022
rect 23664 7958 23716 7964
rect 23676 7002 23704 7958
rect 23768 7206 23796 8191
rect 23860 8090 23888 8298
rect 23848 8084 23900 8090
rect 23848 8026 23900 8032
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 23664 6996 23716 7002
rect 23664 6938 23716 6944
rect 23952 6882 23980 9930
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 24044 9586 24072 9862
rect 24122 9718 24178 9727
rect 24122 9653 24178 9662
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 23676 6854 23980 6882
rect 23480 4966 23532 4972
rect 23570 4992 23626 5001
rect 23570 4927 23626 4936
rect 23388 4752 23440 4758
rect 23388 4694 23440 4700
rect 23400 4146 23428 4694
rect 23570 4312 23626 4321
rect 23570 4247 23626 4256
rect 23388 4140 23440 4146
rect 23388 4082 23440 4088
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23388 3120 23440 3126
rect 23492 3097 23520 3674
rect 23584 3194 23612 4247
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23388 3062 23440 3068
rect 23478 3088 23534 3097
rect 23400 2961 23428 3062
rect 23478 3023 23534 3032
rect 23584 2990 23612 3130
rect 23572 2984 23624 2990
rect 23386 2952 23442 2961
rect 23572 2926 23624 2932
rect 23386 2887 23442 2896
rect 23400 2650 23428 2887
rect 23572 2848 23624 2854
rect 23572 2790 23624 2796
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 22926 776 22982 785
rect 22926 711 22982 720
rect 23584 480 23612 2790
rect 23676 2582 23704 6854
rect 23756 6656 23808 6662
rect 23756 6598 23808 6604
rect 23768 6118 23796 6598
rect 23848 6248 23900 6254
rect 23848 6190 23900 6196
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23768 4078 23796 5850
rect 23860 5778 23888 6190
rect 23940 5840 23992 5846
rect 23940 5782 23992 5788
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 23846 5536 23902 5545
rect 23846 5471 23902 5480
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23768 3777 23796 3878
rect 23754 3768 23810 3777
rect 23754 3703 23810 3712
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23664 2576 23716 2582
rect 23664 2518 23716 2524
rect 23768 1465 23796 3130
rect 23860 2854 23888 5471
rect 23952 4758 23980 5782
rect 23940 4752 23992 4758
rect 23940 4694 23992 4700
rect 24032 3052 24084 3058
rect 24032 2994 24084 3000
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 24044 1601 24072 2994
rect 24136 2836 24164 9653
rect 24228 9586 24256 10134
rect 24320 9994 24348 10406
rect 24504 10198 24532 10542
rect 24676 10532 24728 10538
rect 24676 10474 24728 10480
rect 24492 10192 24544 10198
rect 24492 10134 24544 10140
rect 24308 9988 24360 9994
rect 24308 9930 24360 9936
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24216 9580 24268 9586
rect 24216 9522 24268 9528
rect 24228 8498 24256 9522
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24228 7818 24256 8434
rect 24216 7812 24268 7818
rect 24216 7754 24268 7760
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24582 7440 24638 7449
rect 24582 7375 24584 7384
rect 24636 7375 24638 7384
rect 24584 7346 24636 7352
rect 24214 6896 24270 6905
rect 24688 6866 24716 10474
rect 24780 9217 24808 12815
rect 24860 12786 24912 12792
rect 24872 10538 24900 12786
rect 24950 12744 25006 12753
rect 24950 12679 24952 12688
rect 25004 12679 25006 12688
rect 24952 12650 25004 12656
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 24964 11257 24992 11290
rect 24950 11248 25006 11257
rect 24950 11183 25006 11192
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24860 10532 24912 10538
rect 24860 10474 24912 10480
rect 24964 10470 24992 11086
rect 24952 10464 25004 10470
rect 24952 10406 25004 10412
rect 24860 10260 24912 10266
rect 24860 10202 24912 10208
rect 24872 9722 24900 10202
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24766 9208 24822 9217
rect 24766 9143 24822 9152
rect 24860 9104 24912 9110
rect 24858 9072 24860 9081
rect 24912 9072 24914 9081
rect 24858 9007 24914 9016
rect 24858 8936 24914 8945
rect 24858 8871 24914 8880
rect 24872 8634 24900 8871
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24768 8560 24820 8566
rect 24768 8502 24820 8508
rect 24780 8129 24808 8502
rect 24766 8120 24822 8129
rect 24766 8055 24822 8064
rect 24214 6831 24216 6840
rect 24268 6831 24270 6840
rect 24676 6860 24728 6866
rect 24216 6802 24268 6808
rect 24676 6802 24728 6808
rect 24228 6338 24256 6802
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24228 6310 24348 6338
rect 24214 6216 24270 6225
rect 24214 6151 24270 6160
rect 24228 5914 24256 6151
rect 24216 5908 24268 5914
rect 24216 5850 24268 5856
rect 24320 5846 24348 6310
rect 24308 5840 24360 5846
rect 24308 5782 24360 5788
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 24228 5574 24256 5714
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 24216 5568 24268 5574
rect 24216 5510 24268 5516
rect 24228 5166 24256 5510
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5370 24716 5646
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24216 5160 24268 5166
rect 24216 5102 24268 5108
rect 24228 4758 24256 5102
rect 24216 4752 24268 4758
rect 24216 4694 24268 4700
rect 24674 4720 24730 4729
rect 24228 4486 24256 4694
rect 24780 4690 24808 8055
rect 24964 7857 24992 10406
rect 25056 8906 25084 17002
rect 25504 16652 25556 16658
rect 25504 16594 25556 16600
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25136 15564 25188 15570
rect 25136 15506 25188 15512
rect 25148 14822 25176 15506
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25136 14816 25188 14822
rect 25136 14758 25188 14764
rect 25148 13569 25176 14758
rect 25134 13560 25190 13569
rect 25134 13495 25190 13504
rect 25240 12850 25268 15302
rect 25228 12844 25280 12850
rect 25228 12786 25280 12792
rect 25136 12300 25188 12306
rect 25424 12288 25452 16390
rect 25516 15910 25544 16594
rect 25504 15904 25556 15910
rect 25504 15846 25556 15852
rect 25136 12242 25188 12248
rect 25240 12260 25452 12288
rect 25148 11558 25176 12242
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 25240 10130 25268 12260
rect 25410 12200 25466 12209
rect 25410 12135 25466 12144
rect 25424 11898 25452 12135
rect 25412 11892 25464 11898
rect 25412 11834 25464 11840
rect 25320 11688 25372 11694
rect 25320 11630 25372 11636
rect 25332 10810 25360 11630
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25228 10124 25280 10130
rect 25280 10084 25360 10112
rect 25228 10066 25280 10072
rect 25332 9722 25360 10084
rect 25412 9920 25464 9926
rect 25412 9862 25464 9868
rect 25320 9716 25372 9722
rect 25320 9658 25372 9664
rect 25228 9512 25280 9518
rect 25226 9480 25228 9489
rect 25280 9480 25282 9489
rect 25226 9415 25282 9424
rect 25136 9376 25188 9382
rect 25136 9318 25188 9324
rect 25044 8900 25096 8906
rect 25044 8842 25096 8848
rect 25042 8528 25098 8537
rect 25042 8463 25098 8472
rect 25056 8430 25084 8463
rect 25044 8424 25096 8430
rect 25148 8401 25176 9318
rect 25228 8900 25280 8906
rect 25228 8842 25280 8848
rect 25044 8366 25096 8372
rect 25134 8392 25190 8401
rect 25134 8327 25190 8336
rect 25240 8294 25268 8842
rect 25228 8288 25280 8294
rect 25228 8230 25280 8236
rect 25134 7984 25190 7993
rect 25134 7919 25190 7928
rect 25044 7880 25096 7886
rect 24950 7848 25006 7857
rect 25044 7822 25096 7828
rect 24950 7783 25006 7792
rect 25056 7546 25084 7822
rect 25148 7546 25176 7919
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25136 6996 25188 7002
rect 25136 6938 25188 6944
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24872 6118 24900 6802
rect 24860 6112 24912 6118
rect 24858 6080 24860 6089
rect 24912 6080 24914 6089
rect 24858 6015 24914 6024
rect 24950 5264 25006 5273
rect 24950 5199 25006 5208
rect 24674 4655 24730 4664
rect 24768 4684 24820 4690
rect 24216 4480 24268 4486
rect 24216 4422 24268 4428
rect 24228 4078 24256 4422
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24216 4072 24268 4078
rect 24216 4014 24268 4020
rect 24688 3641 24716 4655
rect 24768 4626 24820 4632
rect 24780 4282 24808 4626
rect 24964 4622 24992 5199
rect 25042 5128 25098 5137
rect 25042 5063 25098 5072
rect 24952 4616 25004 4622
rect 24952 4558 25004 4564
rect 24768 4276 24820 4282
rect 24768 4218 24820 4224
rect 24952 4072 25004 4078
rect 24952 4014 25004 4020
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 24674 3632 24730 3641
rect 24674 3567 24730 3576
rect 24872 3505 24900 3674
rect 24964 3670 24992 4014
rect 24952 3664 25004 3670
rect 24952 3606 25004 3612
rect 25056 3602 25084 5063
rect 25044 3596 25096 3602
rect 25044 3538 25096 3544
rect 24858 3496 24914 3505
rect 24858 3431 24914 3440
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24228 3058 24256 3334
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 25056 3194 25084 3538
rect 25044 3188 25096 3194
rect 25044 3130 25096 3136
rect 24216 3052 24268 3058
rect 24216 2994 24268 3000
rect 24136 2808 24348 2836
rect 24124 2644 24176 2650
rect 24124 2586 24176 2592
rect 24136 2553 24164 2586
rect 24122 2544 24178 2553
rect 24122 2479 24178 2488
rect 24320 2417 24348 2808
rect 24306 2408 24362 2417
rect 25148 2394 25176 6938
rect 25320 6860 25372 6866
rect 25320 6802 25372 6808
rect 25226 6352 25282 6361
rect 25226 6287 25282 6296
rect 25240 6254 25268 6287
rect 25228 6248 25280 6254
rect 25228 6190 25280 6196
rect 25332 5914 25360 6802
rect 25320 5908 25372 5914
rect 25320 5850 25372 5856
rect 25228 5160 25280 5166
rect 25228 5102 25280 5108
rect 25240 5001 25268 5102
rect 25226 4992 25282 5001
rect 25226 4927 25282 4936
rect 25332 4214 25360 5850
rect 25320 4208 25372 4214
rect 25320 4150 25372 4156
rect 25424 4049 25452 9862
rect 25516 6905 25544 15846
rect 25594 13288 25650 13297
rect 25594 13223 25650 13232
rect 25608 12986 25636 13223
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25608 12782 25636 12922
rect 25596 12776 25648 12782
rect 25596 12718 25648 12724
rect 25596 11076 25648 11082
rect 25596 11018 25648 11024
rect 25608 10470 25636 11018
rect 25596 10464 25648 10470
rect 25596 10406 25648 10412
rect 25502 6896 25558 6905
rect 25502 6831 25558 6840
rect 25608 6798 25636 10406
rect 25688 8424 25740 8430
rect 25688 8366 25740 8372
rect 25596 6792 25648 6798
rect 25596 6734 25648 6740
rect 25504 5024 25556 5030
rect 25504 4966 25556 4972
rect 25410 4040 25466 4049
rect 25410 3975 25466 3984
rect 25320 3596 25372 3602
rect 25320 3538 25372 3544
rect 25332 3194 25360 3538
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 25228 2984 25280 2990
rect 25228 2926 25280 2932
rect 25240 2689 25268 2926
rect 25226 2680 25282 2689
rect 25332 2650 25360 3130
rect 25226 2615 25282 2624
rect 25320 2644 25372 2650
rect 25320 2586 25372 2592
rect 25148 2366 25268 2394
rect 24306 2343 24362 2352
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24584 2032 24636 2038
rect 24584 1974 24636 1980
rect 24030 1592 24086 1601
rect 24030 1527 24086 1536
rect 23754 1456 23810 1465
rect 23754 1391 23810 1400
rect 24596 480 24624 1974
rect 25148 1873 25176 2246
rect 25240 2009 25268 2366
rect 25226 2000 25282 2009
rect 25226 1935 25282 1944
rect 25134 1864 25190 1873
rect 25134 1799 25190 1808
rect 25516 480 25544 4966
rect 25700 4146 25728 8366
rect 25792 7954 25820 19343
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 25780 7948 25832 7954
rect 25780 7890 25832 7896
rect 25792 7546 25820 7890
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 25884 6866 25912 11494
rect 26148 8288 26200 8294
rect 26148 8230 26200 8236
rect 25872 6860 25924 6866
rect 25872 6802 25924 6808
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 25596 3936 25648 3942
rect 25596 3878 25648 3884
rect 25608 2038 25636 3878
rect 26160 2514 26188 8230
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 26148 2508 26200 2514
rect 26148 2450 26200 2456
rect 26160 2310 26188 2450
rect 26148 2304 26200 2310
rect 26148 2246 26200 2252
rect 26160 2145 26188 2246
rect 26146 2136 26202 2145
rect 26146 2071 26202 2080
rect 25596 2032 25648 2038
rect 25596 1974 25648 1980
rect 26528 480 26556 6054
rect 27434 4040 27490 4049
rect 27434 3975 27490 3984
rect 27448 480 27476 3975
rect 478 0 534 480
rect 1398 0 1454 480
rect 2318 0 2374 480
rect 3330 0 3386 480
rect 4250 0 4306 480
rect 5262 0 5318 480
rect 6182 0 6238 480
rect 7194 0 7250 480
rect 8114 0 8170 480
rect 9126 0 9182 480
rect 10046 0 10102 480
rect 11058 0 11114 480
rect 11978 0 12034 480
rect 12990 0 13046 480
rect 13910 0 13966 480
rect 14922 0 14978 480
rect 15842 0 15898 480
rect 16854 0 16910 480
rect 17774 0 17830 480
rect 18786 0 18842 480
rect 19706 0 19762 480
rect 20718 0 20774 480
rect 21638 0 21694 480
rect 22650 0 22706 480
rect 23570 0 23626 480
rect 24582 0 24638 480
rect 25502 0 25558 480
rect 26514 0 26570 480
rect 27434 0 27490 480
<< via2 >>
rect 1398 27240 1454 27296
rect 662 23568 718 23624
rect 1582 25880 1638 25936
rect 1490 24520 1546 24576
rect 2042 23468 2044 23488
rect 2044 23468 2096 23488
rect 2096 23468 2098 23488
rect 2042 23432 2098 23468
rect 1582 23024 1638 23080
rect 2686 22616 2742 22672
rect 2134 22208 2190 22264
rect 1674 21972 1676 21992
rect 1676 21972 1728 21992
rect 1728 21972 1730 21992
rect 1674 21936 1730 21972
rect 1674 21664 1730 21720
rect 1582 20304 1638 20360
rect 1398 19624 1454 19680
rect 1582 18808 1638 18864
rect 1398 17448 1454 17504
rect 1214 9016 1270 9072
rect 1122 7792 1178 7848
rect 478 2352 534 2408
rect 1306 2080 1362 2136
rect 1582 16224 1638 16280
rect 1582 16088 1638 16144
rect 1766 16496 1822 16552
rect 2134 18808 2190 18864
rect 2042 16940 2044 16960
rect 2044 16940 2096 16960
rect 2096 16940 2098 16960
rect 2042 16904 2098 16940
rect 2042 16108 2098 16144
rect 2042 16088 2044 16108
rect 2044 16088 2096 16108
rect 2096 16088 2098 16108
rect 2042 15952 2098 16008
rect 1858 14728 1914 14784
rect 1766 13368 1822 13424
rect 1582 11212 1638 11248
rect 1582 11192 1584 11212
rect 1584 11192 1636 11212
rect 1636 11192 1638 11212
rect 1582 9696 1638 9752
rect 1858 9424 1914 9480
rect 1582 5908 1638 5944
rect 1582 5888 1584 5908
rect 1584 5888 1636 5908
rect 1636 5888 1638 5908
rect 1766 7384 1822 7440
rect 1858 6704 1914 6760
rect 1766 6296 1822 6352
rect 1490 3712 1546 3768
rect 1490 3440 1546 3496
rect 2134 10648 2190 10704
rect 2502 18672 2558 18728
rect 3146 19760 3202 19816
rect 2594 17176 2650 17232
rect 2594 16632 2650 16688
rect 2778 17040 2834 17096
rect 2686 15408 2742 15464
rect 3238 18944 3294 19000
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 4802 24792 4858 24848
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5446 23840 5502 23896
rect 5078 23704 5134 23760
rect 5078 23432 5134 23488
rect 5262 23432 5318 23488
rect 5170 22108 5172 22128
rect 5172 22108 5224 22128
rect 5224 22108 5226 22128
rect 5170 22072 5226 22108
rect 3146 14900 3148 14920
rect 3148 14900 3200 14920
rect 3200 14900 3202 14920
rect 3146 14864 3202 14900
rect 3146 14728 3202 14784
rect 3146 14476 3202 14512
rect 3146 14456 3148 14476
rect 3148 14456 3200 14476
rect 3200 14456 3202 14476
rect 2870 13368 2926 13424
rect 2318 12416 2374 12472
rect 2318 11500 2320 11520
rect 2320 11500 2372 11520
rect 2372 11500 2374 11520
rect 2318 11464 2374 11500
rect 2318 9832 2374 9888
rect 2410 9152 2466 9208
rect 2870 12144 2926 12200
rect 2870 11192 2926 11248
rect 2778 9968 2834 10024
rect 2778 9696 2834 9752
rect 2502 7112 2558 7168
rect 2410 4800 2466 4856
rect 3146 12416 3202 12472
rect 3146 8372 3148 8392
rect 3148 8372 3200 8392
rect 3200 8372 3202 8392
rect 3146 8336 3202 8372
rect 3330 15544 3386 15600
rect 3330 12316 3332 12336
rect 3332 12316 3384 12336
rect 3384 12316 3386 12336
rect 3330 12280 3386 12316
rect 3330 9288 3386 9344
rect 3238 7928 3294 7984
rect 2962 6840 3018 6896
rect 2778 5616 2834 5672
rect 2686 5072 2742 5128
rect 2962 5344 3018 5400
rect 2778 4936 2834 4992
rect 2870 4800 2926 4856
rect 2410 4120 2466 4176
rect 1582 3168 1638 3224
rect 1766 3032 1822 3088
rect 2686 4020 2688 4040
rect 2688 4020 2740 4040
rect 2740 4020 2742 4040
rect 2686 3984 2742 4020
rect 3146 7248 3202 7304
rect 3790 19624 3846 19680
rect 3882 19352 3938 19408
rect 3882 19216 3938 19272
rect 4066 19080 4122 19136
rect 3698 15972 3754 16008
rect 3698 15952 3700 15972
rect 3700 15952 3752 15972
rect 3752 15952 3754 15972
rect 3606 15680 3662 15736
rect 4066 16788 4122 16824
rect 4066 16768 4068 16788
rect 4068 16768 4120 16788
rect 4120 16768 4122 16788
rect 3974 16632 4030 16688
rect 4066 14864 4122 14920
rect 3882 8472 3938 8528
rect 3422 5616 3478 5672
rect 3698 5616 3754 5672
rect 1490 2896 1546 2952
rect 1490 2352 1546 2408
rect 2134 1808 2190 1864
rect 2502 2760 2558 2816
rect 3238 1400 3294 1456
rect 2778 720 2834 776
rect 3698 5072 3754 5128
rect 3698 4528 3754 4584
rect 4158 7928 4214 7984
rect 3882 5208 3938 5264
rect 3882 5092 3938 5128
rect 3882 5072 3884 5092
rect 3884 5072 3936 5092
rect 3936 5072 3938 5092
rect 4158 4664 4214 4720
rect 3790 3576 3846 3632
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 7654 24656 7710 24712
rect 8574 23704 8630 23760
rect 8942 23604 8944 23624
rect 8944 23604 8996 23624
rect 8996 23604 8998 23624
rect 8942 23568 8998 23604
rect 9126 23468 9128 23488
rect 9128 23468 9180 23488
rect 9180 23468 9182 23488
rect 9126 23432 9182 23468
rect 6274 22772 6330 22808
rect 6274 22752 6276 22772
rect 6276 22752 6328 22772
rect 6328 22752 6330 22772
rect 5538 21972 5540 21992
rect 5540 21972 5592 21992
rect 5592 21972 5594 21992
rect 5538 21936 5594 21972
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 6274 21412 6330 21448
rect 6274 21392 6276 21412
rect 6276 21392 6328 21412
rect 6328 21392 6330 21412
rect 5078 20304 5134 20360
rect 4710 17196 4766 17232
rect 4710 17176 4712 17196
rect 4712 17176 4764 17196
rect 4764 17176 4766 17196
rect 5354 18264 5410 18320
rect 4618 13252 4674 13288
rect 4618 13232 4620 13252
rect 4620 13232 4672 13252
rect 4672 13232 4674 13252
rect 5262 15816 5318 15872
rect 5170 13912 5226 13968
rect 4986 13368 5042 13424
rect 4710 11192 4766 11248
rect 5078 11620 5134 11656
rect 5078 11600 5080 11620
rect 5080 11600 5132 11620
rect 5132 11600 5134 11620
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5906 19896 5962 19952
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 6090 17856 6146 17912
rect 6090 16904 6146 16960
rect 5906 16632 5962 16688
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5262 10376 5318 10432
rect 5262 9832 5318 9888
rect 4986 7656 5042 7712
rect 4526 6196 4528 6216
rect 4528 6196 4580 6216
rect 4580 6196 4582 6216
rect 4526 6160 4582 6196
rect 4894 6316 4950 6352
rect 4894 6296 4896 6316
rect 4896 6296 4948 6316
rect 4948 6296 4950 6316
rect 4802 5888 4858 5944
rect 4894 5616 4950 5672
rect 4434 3712 4490 3768
rect 3882 1536 3938 1592
rect 4986 3032 5042 3088
rect 5170 2624 5226 2680
rect 4986 2488 5042 2544
rect 4526 2352 4582 2408
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6366 17448 6422 17504
rect 6182 14068 6238 14104
rect 6182 14048 6184 14068
rect 6184 14048 6236 14068
rect 6236 14048 6238 14068
rect 6090 12416 6146 12472
rect 6550 15564 6606 15600
rect 6550 15544 6552 15564
rect 6552 15544 6604 15564
rect 6604 15544 6606 15564
rect 6642 12960 6698 13016
rect 5998 10240 6054 10296
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5446 8200 5502 8256
rect 5814 8336 5870 8392
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 6366 8472 6422 8528
rect 6550 8472 6606 8528
rect 6550 7828 6552 7848
rect 6552 7828 6604 7848
rect 6604 7828 6606 7848
rect 6550 7792 6606 7828
rect 6090 6976 6146 7032
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 6274 5908 6330 5944
rect 6274 5888 6276 5908
rect 6276 5888 6328 5908
rect 6328 5888 6330 5908
rect 5906 5652 5908 5672
rect 5908 5652 5960 5672
rect 5960 5652 5962 5672
rect 5906 5616 5962 5652
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 6366 4936 6422 4992
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 7470 22072 7526 22128
rect 7010 18264 7066 18320
rect 6826 17856 6882 17912
rect 7562 19760 7618 19816
rect 7194 15408 7250 15464
rect 7010 11500 7012 11520
rect 7012 11500 7064 11520
rect 7064 11500 7066 11520
rect 7010 11464 7066 11500
rect 6918 10240 6974 10296
rect 6826 9968 6882 10024
rect 7286 9560 7342 9616
rect 7286 9152 7342 9208
rect 6918 7248 6974 7304
rect 7102 7284 7104 7304
rect 7104 7284 7156 7304
rect 7156 7284 7158 7304
rect 7102 7248 7158 7284
rect 7194 7112 7250 7168
rect 6366 4256 6422 4312
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5998 2896 6054 2952
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5446 1944 5502 2000
rect 5998 1672 6054 1728
rect 7286 6840 7342 6896
rect 7470 16768 7526 16824
rect 8298 22888 8354 22944
rect 7838 22072 7894 22128
rect 8022 20984 8078 21040
rect 7746 19080 7802 19136
rect 7746 18536 7802 18592
rect 8850 22480 8906 22536
rect 8850 22208 8906 22264
rect 8390 19352 8446 19408
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10690 24268 10746 24304
rect 10690 24248 10692 24268
rect 10692 24248 10744 24268
rect 10744 24248 10746 24268
rect 9678 19916 9734 19952
rect 9678 19896 9680 19916
rect 9680 19896 9732 19916
rect 9732 19896 9734 19916
rect 9218 19352 9274 19408
rect 8666 18944 8722 19000
rect 9494 19252 9496 19272
rect 9496 19252 9548 19272
rect 9548 19252 9550 19272
rect 9494 19216 9550 19252
rect 8390 18672 8446 18728
rect 8666 18164 8668 18184
rect 8668 18164 8720 18184
rect 8720 18164 8722 18184
rect 8666 18128 8722 18164
rect 8482 17856 8538 17912
rect 8114 17584 8170 17640
rect 9402 18808 9458 18864
rect 8666 14728 8722 14784
rect 8482 14184 8538 14240
rect 8758 14048 8814 14104
rect 7930 13132 7932 13152
rect 7932 13132 7984 13152
rect 7984 13132 7986 13152
rect 7930 13096 7986 13132
rect 8298 13268 8300 13288
rect 8300 13268 8352 13288
rect 8352 13268 8354 13288
rect 8298 13232 8354 13268
rect 7286 6296 7342 6352
rect 7838 10668 7894 10704
rect 7838 10648 7840 10668
rect 7840 10648 7892 10668
rect 7892 10648 7894 10668
rect 7470 2624 7526 2680
rect 7746 3612 7748 3632
rect 7748 3612 7800 3632
rect 7800 3612 7802 3632
rect 7746 3576 7802 3612
rect 9310 15852 9312 15872
rect 9312 15852 9364 15872
rect 9364 15852 9366 15872
rect 9310 15816 9366 15852
rect 9218 13232 9274 13288
rect 9586 15564 9642 15600
rect 9586 15544 9588 15564
rect 9588 15544 9640 15564
rect 9640 15544 9642 15564
rect 8850 12008 8906 12064
rect 8482 10648 8538 10704
rect 8758 7964 8760 7984
rect 8760 7964 8812 7984
rect 8812 7964 8814 7984
rect 8758 7928 8814 7964
rect 8298 7792 8354 7848
rect 8298 7384 8354 7440
rect 8206 7112 8262 7168
rect 8390 6976 8446 7032
rect 8574 6840 8630 6896
rect 8390 5364 8446 5400
rect 8390 5344 8392 5364
rect 8392 5344 8444 5364
rect 8444 5344 8446 5364
rect 8758 7828 8760 7848
rect 8760 7828 8812 7848
rect 8812 7828 8814 7848
rect 8758 7792 8814 7828
rect 8942 11772 8944 11792
rect 8944 11772 8996 11792
rect 8996 11772 8998 11792
rect 8942 11736 8998 11772
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 11518 24656 11574 24712
rect 11150 24384 11206 24440
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10506 20984 10562 21040
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10046 18536 10102 18592
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 9770 15680 9826 15736
rect 9954 14728 10010 14784
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10690 16360 10746 16416
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10598 15136 10654 15192
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10322 12960 10378 13016
rect 10046 12416 10102 12472
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 9678 10376 9734 10432
rect 9218 8900 9274 8936
rect 9218 8880 9220 8900
rect 9220 8880 9272 8900
rect 9272 8880 9274 8900
rect 9770 9288 9826 9344
rect 9586 8200 9642 8256
rect 9402 7384 9458 7440
rect 8850 6740 8852 6760
rect 8852 6740 8904 6760
rect 8904 6740 8906 6760
rect 8850 6704 8906 6740
rect 8666 5616 8722 5672
rect 9034 5208 9090 5264
rect 8942 4528 8998 4584
rect 8114 3984 8170 4040
rect 8574 4020 8576 4040
rect 8576 4020 8628 4040
rect 8628 4020 8630 4040
rect 8574 3984 8630 4020
rect 8114 3168 8170 3224
rect 8666 2760 8722 2816
rect 8298 2524 8300 2544
rect 8300 2524 8352 2544
rect 8352 2524 8354 2544
rect 8298 2488 8354 2524
rect 8574 2488 8630 2544
rect 8850 1400 8906 1456
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10230 9444 10286 9480
rect 10230 9424 10232 9444
rect 10232 9424 10284 9444
rect 10284 9424 10286 9444
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10046 8880 10102 8936
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10506 6296 10562 6352
rect 9862 6024 9918 6080
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10138 5752 10194 5808
rect 9402 4684 9458 4720
rect 9402 4664 9404 4684
rect 9404 4664 9456 4684
rect 9456 4664 9458 4684
rect 9954 4800 10010 4856
rect 9770 4392 9826 4448
rect 9678 4276 9734 4312
rect 9678 4256 9680 4276
rect 9680 4256 9732 4276
rect 9732 4256 9734 4276
rect 9586 3984 9642 4040
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 11334 22380 11336 22400
rect 11336 22380 11388 22400
rect 11388 22380 11390 22400
rect 11334 22344 11390 22380
rect 11334 22072 11390 22128
rect 13174 24384 13230 24440
rect 11794 24248 11850 24304
rect 12438 24248 12494 24304
rect 11150 21004 11206 21040
rect 11150 20984 11152 21004
rect 11152 20984 11204 21004
rect 11204 20984 11206 21004
rect 11058 17604 11114 17640
rect 11058 17584 11060 17604
rect 11060 17584 11112 17604
rect 11112 17584 11114 17604
rect 11058 16632 11114 16688
rect 11058 14592 11114 14648
rect 10874 13912 10930 13968
rect 10874 13504 10930 13560
rect 10874 13232 10930 13288
rect 11058 13776 11114 13832
rect 11058 13252 11114 13288
rect 11058 13232 11060 13252
rect 11060 13232 11112 13252
rect 11112 13232 11114 13252
rect 11058 13096 11114 13152
rect 11058 11636 11060 11656
rect 11060 11636 11112 11656
rect 11112 11636 11114 11656
rect 11058 11600 11114 11636
rect 10782 10648 10838 10704
rect 10874 8200 10930 8256
rect 11058 7112 11114 7168
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10690 3068 10692 3088
rect 10692 3068 10744 3088
rect 10744 3068 10746 3088
rect 10690 3032 10746 3068
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 9494 2388 9496 2408
rect 9496 2388 9548 2408
rect 9548 2388 9550 2408
rect 9494 2352 9550 2388
rect 10966 2896 11022 2952
rect 9770 1944 9826 2000
rect 9954 1944 10010 2000
rect 10782 1400 10838 1456
rect 11242 19080 11298 19136
rect 11518 21936 11574 21992
rect 11518 16632 11574 16688
rect 11518 15544 11574 15600
rect 11334 14048 11390 14104
rect 11334 13776 11390 13832
rect 11242 12144 11298 12200
rect 11426 11736 11482 11792
rect 11518 11600 11574 11656
rect 11426 11192 11482 11248
rect 11702 13368 11758 13424
rect 11610 8744 11666 8800
rect 14554 24112 14610 24168
rect 14278 23704 14334 23760
rect 12714 23568 12770 23624
rect 12162 22752 12218 22808
rect 12070 20304 12126 20360
rect 11978 17584 12034 17640
rect 12070 11328 12126 11384
rect 12070 10104 12126 10160
rect 11886 9560 11942 9616
rect 11518 5072 11574 5128
rect 11334 4020 11336 4040
rect 11336 4020 11388 4040
rect 11388 4020 11390 4040
rect 11334 3984 11390 4020
rect 11242 2760 11298 2816
rect 11150 2508 11206 2544
rect 11150 2488 11152 2508
rect 11152 2488 11204 2508
rect 11204 2488 11206 2508
rect 11426 2352 11482 2408
rect 12438 22616 12494 22672
rect 12714 21392 12770 21448
rect 12346 17040 12402 17096
rect 12438 13932 12494 13968
rect 12438 13912 12440 13932
rect 12440 13912 12492 13932
rect 12492 13912 12494 13932
rect 12622 15136 12678 15192
rect 13082 19216 13138 19272
rect 12898 17448 12954 17504
rect 13266 17076 13268 17096
rect 13268 17076 13320 17096
rect 13320 17076 13322 17096
rect 13266 17040 13322 17076
rect 12530 13776 12586 13832
rect 12346 12552 12402 12608
rect 12438 12280 12494 12336
rect 12714 12008 12770 12064
rect 12806 11056 12862 11112
rect 12714 10124 12770 10160
rect 12714 10104 12716 10124
rect 12716 10104 12768 10124
rect 12768 10104 12770 10124
rect 12530 9424 12586 9480
rect 12162 7112 12218 7168
rect 12070 6860 12126 6896
rect 12070 6840 12072 6860
rect 12072 6840 12124 6860
rect 12124 6840 12126 6860
rect 12806 7656 12862 7712
rect 12990 12144 13046 12200
rect 13542 22888 13598 22944
rect 13542 20984 13598 21040
rect 14002 22500 14058 22536
rect 14002 22480 14004 22500
rect 14004 22480 14056 22500
rect 14056 22480 14058 22500
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14738 24792 14794 24848
rect 14646 23432 14702 23488
rect 17130 24404 17186 24440
rect 17130 24384 17132 24404
rect 17132 24384 17184 24404
rect 17184 24384 17186 24404
rect 16026 24112 16082 24168
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 16210 23860 16266 23896
rect 16210 23840 16212 23860
rect 16212 23840 16264 23860
rect 16264 23840 16266 23860
rect 16026 23604 16028 23624
rect 16028 23604 16080 23624
rect 16080 23604 16082 23624
rect 16026 23568 16082 23604
rect 18234 24656 18290 24712
rect 18234 24248 18290 24304
rect 17406 23840 17462 23896
rect 16762 23432 16818 23488
rect 14462 21936 14518 21992
rect 13542 17856 13598 17912
rect 13910 17992 13966 18048
rect 13542 17176 13598 17232
rect 13358 8880 13414 8936
rect 12990 7928 13046 7984
rect 13174 7384 13230 7440
rect 12898 7248 12954 7304
rect 12162 5616 12218 5672
rect 12070 5364 12126 5400
rect 12070 5344 12072 5364
rect 12072 5344 12124 5364
rect 12124 5344 12126 5364
rect 12162 3612 12164 3632
rect 12164 3612 12216 3632
rect 12216 3612 12218 3632
rect 12162 3576 12218 3612
rect 12162 3188 12218 3224
rect 12162 3168 12164 3188
rect 12164 3168 12216 3188
rect 12216 3168 12218 3188
rect 12622 3576 12678 3632
rect 12530 2644 12586 2680
rect 12530 2624 12532 2644
rect 12532 2624 12584 2644
rect 12584 2624 12586 2644
rect 12714 1536 12770 1592
rect 12898 1536 12954 1592
rect 14278 18128 14334 18184
rect 13634 13948 13636 13968
rect 13636 13948 13688 13968
rect 13688 13948 13690 13968
rect 13634 13912 13690 13948
rect 13082 5208 13138 5264
rect 14554 18672 14610 18728
rect 15566 23180 15622 23216
rect 15566 23160 15568 23180
rect 15568 23160 15620 23180
rect 15620 23160 15622 23180
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15566 20984 15622 21040
rect 15014 20848 15070 20904
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15566 20460 15622 20496
rect 15566 20440 15568 20460
rect 15568 20440 15620 20460
rect 15620 20440 15622 20460
rect 14186 12144 14242 12200
rect 14094 10648 14150 10704
rect 13726 9052 13728 9072
rect 13728 9052 13780 9072
rect 13780 9052 13782 9072
rect 13726 9016 13782 9052
rect 14094 8880 14150 8936
rect 13634 8356 13690 8392
rect 13634 8336 13636 8356
rect 13636 8336 13688 8356
rect 13688 8336 13690 8356
rect 13910 8744 13966 8800
rect 13726 7964 13728 7984
rect 13728 7964 13780 7984
rect 13780 7964 13782 7984
rect 13726 7928 13782 7964
rect 13542 4936 13598 4992
rect 13266 1808 13322 1864
rect 14002 7404 14058 7440
rect 14002 7384 14004 7404
rect 14004 7384 14056 7404
rect 14056 7384 14058 7404
rect 14370 9152 14426 9208
rect 14646 16496 14702 16552
rect 17314 22344 17370 22400
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15658 19216 15714 19272
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14646 14184 14702 14240
rect 14554 12588 14556 12608
rect 14556 12588 14608 12608
rect 14608 12588 14610 12608
rect 14554 12552 14610 12588
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 16670 20848 16726 20904
rect 17038 17856 17094 17912
rect 16486 16768 16542 16824
rect 17222 18808 17278 18864
rect 17314 17720 17370 17776
rect 17130 17584 17186 17640
rect 15474 14456 15530 14512
rect 15382 13912 15438 13968
rect 15198 13776 15254 13832
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15474 12552 15530 12608
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14646 10376 14702 10432
rect 14462 7384 14518 7440
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15382 9424 15438 9480
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15382 7656 15438 7712
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 15014 6976 15070 7032
rect 16118 15408 16174 15464
rect 16394 15020 16450 15056
rect 17222 15544 17278 15600
rect 16394 15000 16396 15020
rect 16396 15000 16448 15020
rect 16448 15000 16450 15020
rect 15842 11056 15898 11112
rect 15566 7248 15622 7304
rect 15290 6704 15346 6760
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14738 5772 14794 5808
rect 14738 5752 14740 5772
rect 14740 5752 14792 5772
rect 14792 5752 14794 5772
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 16210 8744 16266 8800
rect 16026 7520 16082 7576
rect 15842 6432 15898 6488
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15382 4004 15438 4040
rect 15382 3984 15384 4004
rect 15384 3984 15436 4004
rect 15436 3984 15438 4004
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14554 3032 14610 3088
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15474 2760 15530 2816
rect 15658 2644 15714 2680
rect 15658 2624 15660 2644
rect 15660 2624 15712 2644
rect 15712 2624 15714 2644
rect 15382 1808 15438 1864
rect 16946 14728 17002 14784
rect 16394 12688 16450 12744
rect 16486 6568 16542 6624
rect 16486 6160 16542 6216
rect 16854 6840 16910 6896
rect 16670 4664 16726 4720
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 20166 24656 20222 24712
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 18786 24384 18842 24440
rect 21454 23976 21510 24032
rect 20350 23860 20406 23896
rect 22558 24112 22614 24168
rect 20350 23840 20352 23860
rect 20352 23840 20404 23860
rect 20404 23840 20406 23860
rect 21638 23840 21694 23896
rect 23478 27240 23534 27296
rect 24766 25880 24822 25936
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24674 24520 24730 24576
rect 24214 24112 24270 24168
rect 23018 23976 23074 24032
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 21270 23704 21326 23760
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 17590 19352 17646 19408
rect 17130 13504 17186 13560
rect 17130 12824 17186 12880
rect 17222 12588 17224 12608
rect 17224 12588 17276 12608
rect 17276 12588 17278 12608
rect 17222 12552 17278 12588
rect 17038 11600 17094 11656
rect 17314 11212 17370 11248
rect 17314 11192 17316 11212
rect 17316 11192 17368 11212
rect 17368 11192 17370 11212
rect 17406 9460 17408 9480
rect 17408 9460 17460 9480
rect 17460 9460 17462 9480
rect 17406 9424 17462 9460
rect 17958 19116 17960 19136
rect 17960 19116 18012 19136
rect 18012 19116 18014 19136
rect 17958 19080 18014 19116
rect 17774 17076 17776 17096
rect 17776 17076 17828 17096
rect 17828 17076 17830 17096
rect 17774 17040 17830 17076
rect 18234 16632 18290 16688
rect 17682 11056 17738 11112
rect 17590 6704 17646 6760
rect 17406 5616 17462 5672
rect 17590 5072 17646 5128
rect 16854 4120 16910 4176
rect 16394 3168 16450 3224
rect 16486 2216 16542 2272
rect 17130 2080 17186 2136
rect 17130 1672 17186 1728
rect 17314 1672 17370 1728
rect 18510 17176 18566 17232
rect 18602 14728 18658 14784
rect 18326 12552 18382 12608
rect 18602 12552 18658 12608
rect 17866 9444 17922 9480
rect 17866 9424 17868 9444
rect 17868 9424 17920 9444
rect 17920 9424 17922 9444
rect 18142 10648 18198 10704
rect 18050 8744 18106 8800
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19062 19352 19118 19408
rect 19062 19252 19064 19272
rect 19064 19252 19116 19272
rect 19116 19252 19118 19272
rect 19062 19216 19118 19252
rect 19890 19252 19892 19272
rect 19892 19252 19944 19272
rect 19944 19252 19946 19272
rect 19890 19216 19946 19252
rect 19246 19116 19248 19136
rect 19248 19116 19300 19136
rect 19300 19116 19302 19136
rect 19246 19080 19302 19116
rect 19246 18284 19302 18320
rect 19246 18264 19248 18284
rect 19248 18264 19300 18284
rect 19300 18264 19302 18284
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19614 18672 19670 18728
rect 19338 17992 19394 18048
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19246 17448 19302 17504
rect 18786 16224 18842 16280
rect 18970 16768 19026 16824
rect 18878 16088 18934 16144
rect 19062 15272 19118 15328
rect 18878 13232 18934 13288
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19338 14764 19340 14784
rect 19340 14764 19392 14784
rect 19392 14764 19394 14784
rect 19338 14728 19394 14764
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19798 12960 19854 13016
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19522 12280 19578 12336
rect 18970 12144 19026 12200
rect 19338 12180 19340 12200
rect 19340 12180 19392 12200
rect 19392 12180 19394 12200
rect 19338 12144 19394 12180
rect 18878 11636 18880 11656
rect 18880 11636 18932 11656
rect 18932 11636 18934 11656
rect 18878 11600 18934 11636
rect 18878 9696 18934 9752
rect 18694 8608 18750 8664
rect 18326 8200 18382 8256
rect 18050 5344 18106 5400
rect 18326 4936 18382 4992
rect 18326 3304 18382 3360
rect 18878 7792 18934 7848
rect 18970 6160 19026 6216
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19798 8744 19854 8800
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19338 6160 19394 6216
rect 19338 4120 19394 4176
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19430 3984 19486 4040
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19706 4392 19762 4448
rect 20166 13504 20222 13560
rect 20166 11056 20222 11112
rect 20074 9288 20130 9344
rect 20074 8064 20130 8120
rect 20074 7656 20130 7712
rect 20258 7656 20314 7712
rect 20258 6704 20314 6760
rect 20074 6432 20130 6488
rect 20258 6432 20314 6488
rect 20166 6296 20222 6352
rect 20074 6024 20130 6080
rect 19982 3984 20038 4040
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20166 3596 20222 3632
rect 20166 3576 20168 3596
rect 20168 3576 20220 3596
rect 20220 3576 20222 3596
rect 18142 2488 18198 2544
rect 18326 2388 18328 2408
rect 18328 2388 18380 2408
rect 18380 2388 18382 2408
rect 18326 2352 18382 2388
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20810 17740 20866 17776
rect 20810 17720 20812 17740
rect 20812 17720 20864 17740
rect 20864 17720 20866 17740
rect 20718 17176 20774 17232
rect 20810 16904 20866 16960
rect 20718 16632 20774 16688
rect 20626 16360 20682 16416
rect 20442 13096 20498 13152
rect 20534 9424 20590 9480
rect 20534 8608 20590 8664
rect 20718 9560 20774 9616
rect 20442 8064 20498 8120
rect 20626 7792 20682 7848
rect 20718 7384 20774 7440
rect 20534 3848 20590 3904
rect 21638 18672 21694 18728
rect 21270 11872 21326 11928
rect 21086 10376 21142 10432
rect 20902 6160 20958 6216
rect 21178 7148 21180 7168
rect 21180 7148 21232 7168
rect 21232 7148 21234 7168
rect 21178 7112 21234 7148
rect 20994 5752 21050 5808
rect 20902 5208 20958 5264
rect 21454 13268 21456 13288
rect 21456 13268 21508 13288
rect 21508 13268 21510 13288
rect 21454 13232 21510 13268
rect 25778 24248 25834 24304
rect 24766 23432 24822 23488
rect 27158 23432 27214 23488
rect 23386 23160 23442 23216
rect 24582 23160 24638 23216
rect 23754 22480 23810 22536
rect 23662 21528 23718 21584
rect 22190 17584 22246 17640
rect 22006 17448 22062 17504
rect 22098 16224 22154 16280
rect 22190 15544 22246 15600
rect 22098 15444 22100 15464
rect 22100 15444 22152 15464
rect 22152 15444 22154 15464
rect 22098 15408 22154 15444
rect 22282 12144 22338 12200
rect 21546 8472 21602 8528
rect 21454 7384 21510 7440
rect 21546 6196 21548 6216
rect 21548 6196 21600 6216
rect 21600 6196 21602 6216
rect 21546 6160 21602 6196
rect 21178 5072 21234 5128
rect 20810 3440 20866 3496
rect 21178 3732 21234 3768
rect 21178 3712 21180 3732
rect 21180 3712 21232 3732
rect 21232 3712 21234 3732
rect 21362 3304 21418 3360
rect 20626 2644 20682 2680
rect 20626 2624 20628 2644
rect 20628 2624 20680 2644
rect 20680 2624 20682 2644
rect 22190 12008 22246 12064
rect 22190 11328 22246 11384
rect 21914 10104 21970 10160
rect 21822 8200 21878 8256
rect 21914 7384 21970 7440
rect 22282 7112 22338 7168
rect 22466 16904 22522 16960
rect 22466 14456 22522 14512
rect 22466 12280 22522 12336
rect 22466 11328 22522 11384
rect 21822 5344 21878 5400
rect 21914 5228 21970 5264
rect 21914 5208 21916 5228
rect 21916 5208 21968 5228
rect 21968 5208 21970 5228
rect 22466 6296 22522 6352
rect 22374 5092 22430 5128
rect 22374 5072 22376 5092
rect 22376 5072 22428 5092
rect 22428 5072 22430 5092
rect 22926 15988 22928 16008
rect 22928 15988 22980 16008
rect 22980 15988 22982 16008
rect 22926 15952 22982 15988
rect 22834 13368 22890 13424
rect 22834 10512 22890 10568
rect 22834 4020 22836 4040
rect 22836 4020 22888 4040
rect 22888 4020 22890 4040
rect 22834 3984 22890 4020
rect 22374 3188 22430 3224
rect 22374 3168 22376 3188
rect 22376 3168 22428 3188
rect 22428 3168 22430 3188
rect 21546 2080 21602 2136
rect 19706 1944 19762 2000
rect 20718 1672 20774 1728
rect 23018 9696 23074 9752
rect 23018 9288 23074 9344
rect 23018 3848 23074 3904
rect 23478 15308 23480 15328
rect 23480 15308 23532 15328
rect 23532 15308 23534 15328
rect 23478 15272 23534 15308
rect 23386 14864 23442 14920
rect 23478 13776 23534 13832
rect 23478 13504 23534 13560
rect 23202 13368 23258 13424
rect 23294 9696 23350 9752
rect 23202 8780 23204 8800
rect 23204 8780 23256 8800
rect 23256 8780 23258 8800
rect 23202 8744 23258 8780
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24122 20440 24178 20496
rect 24122 19352 24178 19408
rect 24122 17448 24178 17504
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24766 23024 24822 23080
rect 24766 20304 24822 20360
rect 25778 19352 25834 19408
rect 24766 18808 24822 18864
rect 24582 18672 24638 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24582 18300 24584 18320
rect 24584 18300 24636 18320
rect 24636 18300 24638 18320
rect 24582 18264 24638 18300
rect 24674 17448 24730 17504
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 23662 12552 23718 12608
rect 24766 16088 24822 16144
rect 24858 15000 24914 15056
rect 24766 14456 24822 14512
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24030 13640 24086 13696
rect 24030 13504 24086 13560
rect 24214 13388 24270 13424
rect 24214 13368 24216 13388
rect 24216 13368 24268 13388
rect 24268 13368 24270 13388
rect 24030 13096 24086 13152
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24950 14864 25006 14920
rect 24766 12824 24822 12880
rect 24030 12552 24086 12608
rect 24030 12144 24086 12200
rect 23754 11600 23810 11656
rect 23754 10376 23810 10432
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24122 9968 24178 10024
rect 23478 7656 23534 7712
rect 23478 7112 23534 7168
rect 23202 5616 23258 5672
rect 23386 6568 23442 6624
rect 23386 6332 23388 6352
rect 23388 6332 23440 6352
rect 23440 6332 23442 6352
rect 23386 6296 23442 6332
rect 23754 8200 23810 8256
rect 24122 9662 24178 9718
rect 23570 4936 23626 4992
rect 23570 4256 23626 4312
rect 23478 3032 23534 3088
rect 23386 2896 23442 2952
rect 22926 720 22982 776
rect 23846 5480 23902 5536
rect 23754 3712 23810 3768
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24582 7404 24638 7440
rect 24582 7384 24584 7404
rect 24584 7384 24636 7404
rect 24636 7384 24638 7404
rect 24214 6860 24270 6896
rect 24950 12708 25006 12744
rect 24950 12688 24952 12708
rect 24952 12688 25004 12708
rect 25004 12688 25006 12708
rect 24950 11192 25006 11248
rect 24766 9152 24822 9208
rect 24858 9052 24860 9072
rect 24860 9052 24912 9072
rect 24912 9052 24914 9072
rect 24858 9016 24914 9052
rect 24858 8880 24914 8936
rect 24766 8064 24822 8120
rect 24214 6840 24216 6860
rect 24216 6840 24268 6860
rect 24268 6840 24270 6860
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24214 6160 24270 6216
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24674 4664 24730 4720
rect 25134 13504 25190 13560
rect 25410 12144 25466 12200
rect 25226 9460 25228 9480
rect 25228 9460 25280 9480
rect 25280 9460 25282 9480
rect 25226 9424 25282 9460
rect 25042 8472 25098 8528
rect 25134 8336 25190 8392
rect 25134 7928 25190 7984
rect 24950 7792 25006 7848
rect 24858 6060 24860 6080
rect 24860 6060 24912 6080
rect 24912 6060 24914 6080
rect 24858 6024 24914 6060
rect 24950 5208 25006 5264
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 25042 5072 25098 5128
rect 24674 3576 24730 3632
rect 24858 3440 24914 3496
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24122 2488 24178 2544
rect 24306 2352 24362 2408
rect 25226 6296 25282 6352
rect 25226 4936 25282 4992
rect 25594 13232 25650 13288
rect 25502 6840 25558 6896
rect 25410 3984 25466 4040
rect 25226 2624 25282 2680
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24030 1536 24086 1592
rect 23754 1400 23810 1456
rect 25226 1944 25282 2000
rect 25134 1808 25190 1864
rect 26146 2080 26202 2136
rect 27434 3984 27490 4040
<< metal3 >>
rect 0 27298 480 27328
rect 1393 27298 1459 27301
rect 0 27296 1459 27298
rect 0 27240 1398 27296
rect 1454 27240 1459 27296
rect 0 27238 1459 27240
rect 0 27208 480 27238
rect 1393 27235 1459 27238
rect 23473 27298 23539 27301
rect 27520 27298 28000 27328
rect 23473 27296 28000 27298
rect 23473 27240 23478 27296
rect 23534 27240 28000 27296
rect 23473 27238 28000 27240
rect 23473 27235 23539 27238
rect 27520 27208 28000 27238
rect 0 25938 480 25968
rect 1577 25938 1643 25941
rect 0 25936 1643 25938
rect 0 25880 1582 25936
rect 1638 25880 1643 25936
rect 0 25878 1643 25880
rect 0 25848 480 25878
rect 1577 25875 1643 25878
rect 24761 25938 24827 25941
rect 27520 25938 28000 25968
rect 24761 25936 28000 25938
rect 24761 25880 24766 25936
rect 24822 25880 28000 25936
rect 24761 25878 28000 25880
rect 24761 25875 24827 25878
rect 27520 25848 28000 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 4797 24850 4863 24853
rect 14733 24850 14799 24853
rect 4797 24848 14799 24850
rect 4797 24792 4802 24848
rect 4858 24792 14738 24848
rect 14794 24792 14799 24848
rect 4797 24790 14799 24792
rect 4797 24787 4863 24790
rect 14733 24787 14799 24790
rect 7649 24714 7715 24717
rect 11513 24714 11579 24717
rect 7649 24712 11579 24714
rect 7649 24656 7654 24712
rect 7710 24656 11518 24712
rect 11574 24656 11579 24712
rect 7649 24654 11579 24656
rect 7649 24651 7715 24654
rect 11513 24651 11579 24654
rect 18229 24714 18295 24717
rect 20161 24714 20227 24717
rect 18229 24712 20227 24714
rect 18229 24656 18234 24712
rect 18290 24656 20166 24712
rect 20222 24656 20227 24712
rect 18229 24654 20227 24656
rect 18229 24651 18295 24654
rect 20161 24651 20227 24654
rect 0 24578 480 24608
rect 1485 24578 1551 24581
rect 0 24576 1551 24578
rect 0 24520 1490 24576
rect 1546 24520 1551 24576
rect 0 24518 1551 24520
rect 0 24488 480 24518
rect 1485 24515 1551 24518
rect 24669 24578 24735 24581
rect 27520 24578 28000 24608
rect 24669 24576 28000 24578
rect 24669 24520 24674 24576
rect 24730 24520 28000 24576
rect 24669 24518 28000 24520
rect 24669 24515 24735 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 27520 24488 28000 24518
rect 19610 24447 19930 24448
rect 11145 24442 11211 24445
rect 13169 24442 13235 24445
rect 11145 24440 13235 24442
rect 11145 24384 11150 24440
rect 11206 24384 13174 24440
rect 13230 24384 13235 24440
rect 11145 24382 13235 24384
rect 11145 24379 11211 24382
rect 13169 24379 13235 24382
rect 17125 24442 17191 24445
rect 18781 24442 18847 24445
rect 17125 24440 18847 24442
rect 17125 24384 17130 24440
rect 17186 24384 18786 24440
rect 18842 24384 18847 24440
rect 17125 24382 18847 24384
rect 17125 24379 17191 24382
rect 18781 24379 18847 24382
rect 10685 24306 10751 24309
rect 11789 24306 11855 24309
rect 12433 24306 12499 24309
rect 10685 24304 12499 24306
rect 10685 24248 10690 24304
rect 10746 24248 11794 24304
rect 11850 24248 12438 24304
rect 12494 24248 12499 24304
rect 10685 24246 12499 24248
rect 10685 24243 10751 24246
rect 11789 24243 11855 24246
rect 12433 24243 12499 24246
rect 18229 24306 18295 24309
rect 25773 24306 25839 24309
rect 18229 24304 25839 24306
rect 18229 24248 18234 24304
rect 18290 24248 25778 24304
rect 25834 24248 25839 24304
rect 18229 24246 25839 24248
rect 18229 24243 18295 24246
rect 25773 24243 25839 24246
rect 14549 24170 14615 24173
rect 16021 24170 16087 24173
rect 14549 24168 16087 24170
rect 14549 24112 14554 24168
rect 14610 24112 16026 24168
rect 16082 24112 16087 24168
rect 14549 24110 16087 24112
rect 14549 24107 14615 24110
rect 16021 24107 16087 24110
rect 22553 24170 22619 24173
rect 24209 24170 24275 24173
rect 22553 24168 24275 24170
rect 22553 24112 22558 24168
rect 22614 24112 24214 24168
rect 24270 24112 24275 24168
rect 22553 24110 24275 24112
rect 22553 24107 22619 24110
rect 24209 24107 24275 24110
rect 21449 24034 21515 24037
rect 23013 24034 23079 24037
rect 21449 24032 23079 24034
rect 21449 23976 21454 24032
rect 21510 23976 23018 24032
rect 23074 23976 23079 24032
rect 21449 23974 23079 23976
rect 21449 23971 21515 23974
rect 23013 23971 23079 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 5441 23898 5507 23901
rect 2822 23896 5507 23898
rect 2822 23840 5446 23896
rect 5502 23840 5507 23896
rect 2822 23838 5507 23840
rect 657 23626 723 23629
rect 2822 23626 2882 23838
rect 5441 23835 5507 23838
rect 16205 23898 16271 23901
rect 17401 23898 17467 23901
rect 16205 23896 17467 23898
rect 16205 23840 16210 23896
rect 16266 23840 17406 23896
rect 17462 23840 17467 23896
rect 16205 23838 17467 23840
rect 16205 23835 16271 23838
rect 17401 23835 17467 23838
rect 20345 23898 20411 23901
rect 21633 23898 21699 23901
rect 20345 23896 21699 23898
rect 20345 23840 20350 23896
rect 20406 23840 21638 23896
rect 21694 23840 21699 23896
rect 20345 23838 21699 23840
rect 20345 23835 20411 23838
rect 21633 23835 21699 23838
rect 5073 23762 5139 23765
rect 8569 23762 8635 23765
rect 5073 23760 8635 23762
rect 5073 23704 5078 23760
rect 5134 23704 8574 23760
rect 8630 23704 8635 23760
rect 5073 23702 8635 23704
rect 5073 23699 5139 23702
rect 8569 23699 8635 23702
rect 14273 23762 14339 23765
rect 21265 23762 21331 23765
rect 14273 23760 21331 23762
rect 14273 23704 14278 23760
rect 14334 23704 21270 23760
rect 21326 23704 21331 23760
rect 14273 23702 21331 23704
rect 14273 23699 14339 23702
rect 21265 23699 21331 23702
rect 657 23624 2882 23626
rect 657 23568 662 23624
rect 718 23568 2882 23624
rect 657 23566 2882 23568
rect 657 23563 723 23566
rect 2998 23564 3004 23628
rect 3068 23626 3074 23628
rect 8937 23626 9003 23629
rect 3068 23624 9003 23626
rect 3068 23568 8942 23624
rect 8998 23568 9003 23624
rect 3068 23566 9003 23568
rect 3068 23564 3074 23566
rect 8937 23563 9003 23566
rect 12709 23626 12775 23629
rect 16021 23626 16087 23629
rect 12709 23624 16087 23626
rect 12709 23568 12714 23624
rect 12770 23568 16026 23624
rect 16082 23568 16087 23624
rect 12709 23566 16087 23568
rect 12709 23563 12775 23566
rect 16021 23563 16087 23566
rect 2037 23490 2103 23493
rect 5073 23490 5139 23493
rect 2037 23488 5139 23490
rect 2037 23432 2042 23488
rect 2098 23432 5078 23488
rect 5134 23432 5139 23488
rect 2037 23430 5139 23432
rect 2037 23427 2103 23430
rect 5073 23427 5139 23430
rect 5257 23490 5323 23493
rect 9121 23490 9187 23493
rect 5257 23488 9187 23490
rect 5257 23432 5262 23488
rect 5318 23432 9126 23488
rect 9182 23432 9187 23488
rect 5257 23430 9187 23432
rect 5257 23427 5323 23430
rect 9121 23427 9187 23430
rect 14641 23490 14707 23493
rect 16757 23490 16823 23493
rect 14641 23488 16823 23490
rect 14641 23432 14646 23488
rect 14702 23432 16762 23488
rect 16818 23432 16823 23488
rect 14641 23430 16823 23432
rect 14641 23427 14707 23430
rect 16757 23427 16823 23430
rect 24761 23490 24827 23493
rect 27153 23490 27219 23493
rect 24761 23488 27219 23490
rect 24761 23432 24766 23488
rect 24822 23432 27158 23488
rect 27214 23432 27219 23488
rect 24761 23430 27219 23432
rect 24761 23427 24827 23430
rect 27153 23427 27219 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 15561 23218 15627 23221
rect 23381 23218 23447 23221
rect 24577 23218 24643 23221
rect 15561 23216 24643 23218
rect 15561 23160 15566 23216
rect 15622 23160 23386 23216
rect 23442 23160 24582 23216
rect 24638 23160 24643 23216
rect 15561 23158 24643 23160
rect 15561 23155 15627 23158
rect 23381 23155 23447 23158
rect 24577 23155 24643 23158
rect 0 23082 480 23112
rect 1577 23082 1643 23085
rect 0 23080 1643 23082
rect 0 23024 1582 23080
rect 1638 23024 1643 23080
rect 0 23022 1643 23024
rect 0 22992 480 23022
rect 1577 23019 1643 23022
rect 24761 23082 24827 23085
rect 27520 23082 28000 23112
rect 24761 23080 28000 23082
rect 24761 23024 24766 23080
rect 24822 23024 28000 23080
rect 24761 23022 28000 23024
rect 24761 23019 24827 23022
rect 27520 22992 28000 23022
rect 8293 22946 8359 22949
rect 13537 22946 13603 22949
rect 8293 22944 13603 22946
rect 8293 22888 8298 22944
rect 8354 22888 13542 22944
rect 13598 22888 13603 22944
rect 8293 22886 13603 22888
rect 8293 22883 8359 22886
rect 13537 22883 13603 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 6269 22810 6335 22813
rect 12157 22810 12223 22813
rect 6269 22808 12223 22810
rect 6269 22752 6274 22808
rect 6330 22752 12162 22808
rect 12218 22752 12223 22808
rect 6269 22750 12223 22752
rect 6269 22747 6335 22750
rect 12157 22747 12223 22750
rect 2681 22674 2747 22677
rect 12433 22674 12499 22677
rect 2681 22672 12499 22674
rect 2681 22616 2686 22672
rect 2742 22616 12438 22672
rect 12494 22616 12499 22672
rect 2681 22614 12499 22616
rect 2681 22611 2747 22614
rect 12433 22611 12499 22614
rect 8845 22538 8911 22541
rect 13997 22538 14063 22541
rect 23749 22538 23815 22541
rect 8845 22536 23815 22538
rect 8845 22480 8850 22536
rect 8906 22480 14002 22536
rect 14058 22480 23754 22536
rect 23810 22480 23815 22536
rect 8845 22478 23815 22480
rect 8845 22475 8911 22478
rect 13997 22475 14063 22478
rect 23749 22475 23815 22478
rect 11329 22402 11395 22405
rect 17309 22402 17375 22405
rect 11329 22400 17375 22402
rect 11329 22344 11334 22400
rect 11390 22344 17314 22400
rect 17370 22344 17375 22400
rect 11329 22342 17375 22344
rect 11329 22339 11395 22342
rect 17309 22339 17375 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 2129 22266 2195 22269
rect 8845 22266 8911 22269
rect 2129 22264 8911 22266
rect 2129 22208 2134 22264
rect 2190 22208 8850 22264
rect 8906 22208 8911 22264
rect 2129 22206 8911 22208
rect 2129 22203 2195 22206
rect 8845 22203 8911 22206
rect 5165 22130 5231 22133
rect 7465 22130 7531 22133
rect 5165 22128 7531 22130
rect 5165 22072 5170 22128
rect 5226 22072 7470 22128
rect 7526 22072 7531 22128
rect 5165 22070 7531 22072
rect 5165 22067 5231 22070
rect 7465 22067 7531 22070
rect 7833 22130 7899 22133
rect 11329 22130 11395 22133
rect 7833 22128 11395 22130
rect 7833 22072 7838 22128
rect 7894 22072 11334 22128
rect 11390 22072 11395 22128
rect 7833 22070 11395 22072
rect 7833 22067 7899 22070
rect 11329 22067 11395 22070
rect 1669 21994 1735 21997
rect 5533 21994 5599 21997
rect 1669 21992 5599 21994
rect 1669 21936 1674 21992
rect 1730 21936 5538 21992
rect 5594 21936 5599 21992
rect 1669 21934 5599 21936
rect 1669 21931 1735 21934
rect 5533 21931 5599 21934
rect 11513 21994 11579 21997
rect 14457 21994 14523 21997
rect 11513 21992 14523 21994
rect 11513 21936 11518 21992
rect 11574 21936 14462 21992
rect 14518 21936 14523 21992
rect 11513 21934 14523 21936
rect 11513 21931 11579 21934
rect 14457 21931 14523 21934
rect 5610 21792 5930 21793
rect 0 21722 480 21752
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 1669 21722 1735 21725
rect 27520 21722 28000 21752
rect 0 21720 1735 21722
rect 0 21664 1674 21720
rect 1730 21664 1735 21720
rect 0 21662 1735 21664
rect 0 21632 480 21662
rect 1669 21659 1735 21662
rect 24718 21662 28000 21722
rect 23657 21586 23723 21589
rect 24718 21586 24778 21662
rect 27520 21632 28000 21662
rect 23657 21584 24778 21586
rect 23657 21528 23662 21584
rect 23718 21528 24778 21584
rect 23657 21526 24778 21528
rect 23657 21523 23723 21526
rect 6269 21450 6335 21453
rect 12709 21450 12775 21453
rect 6269 21448 12775 21450
rect 6269 21392 6274 21448
rect 6330 21392 12714 21448
rect 12770 21392 12775 21448
rect 6269 21390 12775 21392
rect 6269 21387 6335 21390
rect 12709 21387 12775 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 8017 21042 8083 21045
rect 10501 21042 10567 21045
rect 11145 21042 11211 21045
rect 8017 21040 11211 21042
rect 8017 20984 8022 21040
rect 8078 20984 10506 21040
rect 10562 20984 11150 21040
rect 11206 20984 11211 21040
rect 8017 20982 11211 20984
rect 8017 20979 8083 20982
rect 10501 20979 10567 20982
rect 11145 20979 11211 20982
rect 13537 21042 13603 21045
rect 15561 21042 15627 21045
rect 13537 21040 15627 21042
rect 13537 20984 13542 21040
rect 13598 20984 15566 21040
rect 15622 20984 15627 21040
rect 13537 20982 15627 20984
rect 13537 20979 13603 20982
rect 15561 20979 15627 20982
rect 15009 20906 15075 20909
rect 16665 20906 16731 20909
rect 15009 20904 16731 20906
rect 15009 20848 15014 20904
rect 15070 20848 16670 20904
rect 16726 20848 16731 20904
rect 15009 20846 16731 20848
rect 15009 20843 15075 20846
rect 16665 20843 16731 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 15561 20498 15627 20501
rect 24117 20498 24183 20501
rect 15561 20496 24183 20498
rect 15561 20440 15566 20496
rect 15622 20440 24122 20496
rect 24178 20440 24183 20496
rect 15561 20438 24183 20440
rect 15561 20435 15627 20438
rect 24117 20435 24183 20438
rect 0 20362 480 20392
rect 1577 20362 1643 20365
rect 0 20360 1643 20362
rect 0 20304 1582 20360
rect 1638 20304 1643 20360
rect 0 20302 1643 20304
rect 0 20272 480 20302
rect 1577 20299 1643 20302
rect 5073 20362 5139 20365
rect 12065 20362 12131 20365
rect 5073 20360 12131 20362
rect 5073 20304 5078 20360
rect 5134 20304 12070 20360
rect 12126 20304 12131 20360
rect 5073 20302 12131 20304
rect 5073 20299 5139 20302
rect 12065 20299 12131 20302
rect 24761 20362 24827 20365
rect 27520 20362 28000 20392
rect 24761 20360 28000 20362
rect 24761 20304 24766 20360
rect 24822 20304 28000 20360
rect 24761 20302 28000 20304
rect 24761 20299 24827 20302
rect 27520 20272 28000 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 5901 19954 5967 19957
rect 9673 19954 9739 19957
rect 5901 19952 9739 19954
rect 5901 19896 5906 19952
rect 5962 19896 9678 19952
rect 9734 19896 9739 19952
rect 5901 19894 9739 19896
rect 5901 19891 5967 19894
rect 9673 19891 9739 19894
rect 3141 19818 3207 19821
rect 7557 19818 7623 19821
rect 3141 19816 7623 19818
rect 3141 19760 3146 19816
rect 3202 19760 7562 19816
rect 7618 19760 7623 19816
rect 3141 19758 7623 19760
rect 3141 19755 3207 19758
rect 7557 19755 7623 19758
rect 1393 19682 1459 19685
rect 3785 19682 3851 19685
rect 1393 19680 3851 19682
rect 1393 19624 1398 19680
rect 1454 19624 3790 19680
rect 3846 19624 3851 19680
rect 1393 19622 3851 19624
rect 1393 19619 1459 19622
rect 3785 19619 3851 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 3877 19412 3943 19413
rect 3877 19408 3924 19412
rect 3988 19410 3994 19412
rect 8385 19410 8451 19413
rect 9213 19410 9279 19413
rect 17585 19410 17651 19413
rect 19057 19410 19123 19413
rect 3877 19352 3882 19408
rect 3877 19348 3924 19352
rect 3988 19350 4034 19410
rect 8385 19408 19123 19410
rect 8385 19352 8390 19408
rect 8446 19352 9218 19408
rect 9274 19352 17590 19408
rect 17646 19352 19062 19408
rect 19118 19352 19123 19408
rect 8385 19350 19123 19352
rect 3988 19348 3994 19350
rect 3877 19347 3943 19348
rect 8385 19347 8451 19350
rect 9213 19347 9279 19350
rect 17585 19347 17651 19350
rect 19057 19347 19123 19350
rect 24117 19410 24183 19413
rect 25773 19410 25839 19413
rect 24117 19408 25839 19410
rect 24117 19352 24122 19408
rect 24178 19352 25778 19408
rect 25834 19352 25839 19408
rect 24117 19350 25839 19352
rect 24117 19347 24183 19350
rect 25773 19347 25839 19350
rect 3877 19274 3943 19277
rect 9489 19274 9555 19277
rect 3877 19272 9555 19274
rect 3877 19216 3882 19272
rect 3938 19216 9494 19272
rect 9550 19216 9555 19272
rect 3877 19214 9555 19216
rect 3877 19211 3943 19214
rect 9489 19211 9555 19214
rect 13077 19274 13143 19277
rect 15653 19274 15719 19277
rect 19057 19274 19123 19277
rect 19885 19274 19951 19277
rect 13077 19272 19951 19274
rect 13077 19216 13082 19272
rect 13138 19216 15658 19272
rect 15714 19216 19062 19272
rect 19118 19216 19890 19272
rect 19946 19216 19951 19272
rect 13077 19214 19951 19216
rect 13077 19211 13143 19214
rect 15653 19211 15719 19214
rect 19057 19211 19123 19214
rect 19885 19211 19951 19214
rect 4061 19138 4127 19141
rect 7741 19138 7807 19141
rect 4061 19136 7807 19138
rect 4061 19080 4066 19136
rect 4122 19080 7746 19136
rect 7802 19080 7807 19136
rect 4061 19078 7807 19080
rect 4061 19075 4127 19078
rect 7741 19075 7807 19078
rect 11237 19138 11303 19141
rect 17953 19138 18019 19141
rect 19241 19140 19307 19141
rect 19190 19138 19196 19140
rect 11237 19136 18019 19138
rect 11237 19080 11242 19136
rect 11298 19080 17958 19136
rect 18014 19080 18019 19136
rect 11237 19078 18019 19080
rect 19150 19078 19196 19138
rect 19260 19136 19307 19140
rect 19302 19080 19307 19136
rect 11237 19075 11303 19078
rect 17953 19075 18019 19078
rect 19190 19076 19196 19078
rect 19260 19076 19307 19080
rect 19241 19075 19307 19076
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 3233 19002 3299 19005
rect 8661 19002 8727 19005
rect 3233 19000 8727 19002
rect 3233 18944 3238 19000
rect 3294 18944 8666 19000
rect 8722 18944 8727 19000
rect 3233 18942 8727 18944
rect 3233 18939 3299 18942
rect 8661 18939 8727 18942
rect 0 18866 480 18896
rect 1577 18866 1643 18869
rect 0 18864 1643 18866
rect 0 18808 1582 18864
rect 1638 18808 1643 18864
rect 0 18806 1643 18808
rect 0 18776 480 18806
rect 1577 18803 1643 18806
rect 2129 18866 2195 18869
rect 9397 18866 9463 18869
rect 2129 18864 9463 18866
rect 2129 18808 2134 18864
rect 2190 18808 9402 18864
rect 9458 18808 9463 18864
rect 2129 18806 9463 18808
rect 2129 18803 2195 18806
rect 9397 18803 9463 18806
rect 17217 18866 17283 18869
rect 24761 18866 24827 18869
rect 27520 18866 28000 18896
rect 17217 18864 19810 18866
rect 17217 18808 17222 18864
rect 17278 18808 19810 18864
rect 17217 18806 19810 18808
rect 17217 18803 17283 18806
rect 2497 18730 2563 18733
rect 8385 18730 8451 18733
rect 2497 18728 8451 18730
rect 2497 18672 2502 18728
rect 2558 18672 8390 18728
rect 8446 18672 8451 18728
rect 2497 18670 8451 18672
rect 2497 18667 2563 18670
rect 8385 18667 8451 18670
rect 14549 18730 14615 18733
rect 19609 18730 19675 18733
rect 14549 18728 19675 18730
rect 14549 18672 14554 18728
rect 14610 18672 19614 18728
rect 19670 18672 19675 18728
rect 14549 18670 19675 18672
rect 19750 18730 19810 18806
rect 24761 18864 28000 18866
rect 24761 18808 24766 18864
rect 24822 18808 28000 18864
rect 24761 18806 28000 18808
rect 24761 18803 24827 18806
rect 27520 18776 28000 18806
rect 21633 18730 21699 18733
rect 24577 18730 24643 18733
rect 19750 18728 24643 18730
rect 19750 18672 21638 18728
rect 21694 18672 24582 18728
rect 24638 18672 24643 18728
rect 19750 18670 24643 18672
rect 14549 18667 14615 18670
rect 19609 18667 19675 18670
rect 21633 18667 21699 18670
rect 24577 18667 24643 18670
rect 7741 18594 7807 18597
rect 10041 18594 10107 18597
rect 7741 18592 10107 18594
rect 7741 18536 7746 18592
rect 7802 18536 10046 18592
rect 10102 18536 10107 18592
rect 7741 18534 10107 18536
rect 7741 18531 7807 18534
rect 10041 18531 10107 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 5349 18322 5415 18325
rect 7005 18322 7071 18325
rect 5349 18320 7071 18322
rect 5349 18264 5354 18320
rect 5410 18264 7010 18320
rect 7066 18264 7071 18320
rect 5349 18262 7071 18264
rect 5349 18259 5415 18262
rect 7005 18259 7071 18262
rect 19241 18322 19307 18325
rect 24577 18322 24643 18325
rect 19241 18320 24643 18322
rect 19241 18264 19246 18320
rect 19302 18264 24582 18320
rect 24638 18264 24643 18320
rect 19241 18262 24643 18264
rect 19241 18259 19307 18262
rect 24577 18259 24643 18262
rect 8661 18186 8727 18189
rect 14273 18186 14339 18189
rect 8661 18184 14339 18186
rect 8661 18128 8666 18184
rect 8722 18128 14278 18184
rect 14334 18128 14339 18184
rect 8661 18126 14339 18128
rect 8661 18123 8727 18126
rect 14273 18123 14339 18126
rect 13905 18050 13971 18053
rect 19333 18050 19399 18053
rect 13905 18048 19399 18050
rect 13905 17992 13910 18048
rect 13966 17992 19338 18048
rect 19394 17992 19399 18048
rect 13905 17990 19399 17992
rect 13905 17987 13971 17990
rect 19333 17987 19399 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 6085 17914 6151 17917
rect 6821 17914 6887 17917
rect 8477 17914 8543 17917
rect 6085 17912 8543 17914
rect 6085 17856 6090 17912
rect 6146 17856 6826 17912
rect 6882 17856 8482 17912
rect 8538 17856 8543 17912
rect 6085 17854 8543 17856
rect 6085 17851 6151 17854
rect 6821 17851 6887 17854
rect 8477 17851 8543 17854
rect 13537 17914 13603 17917
rect 17033 17914 17099 17917
rect 13537 17912 17099 17914
rect 13537 17856 13542 17912
rect 13598 17856 17038 17912
rect 17094 17856 17099 17912
rect 13537 17854 17099 17856
rect 13537 17851 13603 17854
rect 17033 17851 17099 17854
rect 17309 17778 17375 17781
rect 20805 17778 20871 17781
rect 17309 17776 20871 17778
rect 17309 17720 17314 17776
rect 17370 17720 20810 17776
rect 20866 17720 20871 17776
rect 17309 17718 20871 17720
rect 17309 17715 17375 17718
rect 20805 17715 20871 17718
rect 8109 17642 8175 17645
rect 11053 17642 11119 17645
rect 8109 17640 11119 17642
rect 8109 17584 8114 17640
rect 8170 17584 11058 17640
rect 11114 17584 11119 17640
rect 8109 17582 11119 17584
rect 8109 17579 8175 17582
rect 11053 17579 11119 17582
rect 11973 17642 12039 17645
rect 17125 17642 17191 17645
rect 22185 17642 22251 17645
rect 11973 17640 22251 17642
rect 11973 17584 11978 17640
rect 12034 17584 17130 17640
rect 17186 17584 22190 17640
rect 22246 17584 22251 17640
rect 11973 17582 22251 17584
rect 11973 17579 12039 17582
rect 17125 17579 17191 17582
rect 22185 17579 22251 17582
rect 0 17506 480 17536
rect 1393 17506 1459 17509
rect 0 17504 1459 17506
rect 0 17448 1398 17504
rect 1454 17448 1459 17504
rect 0 17446 1459 17448
rect 0 17416 480 17446
rect 1393 17443 1459 17446
rect 6361 17506 6427 17509
rect 12893 17506 12959 17509
rect 6361 17504 12959 17506
rect 6361 17448 6366 17504
rect 6422 17448 12898 17504
rect 12954 17448 12959 17504
rect 6361 17446 12959 17448
rect 6361 17443 6427 17446
rect 12893 17443 12959 17446
rect 19241 17506 19307 17509
rect 22001 17506 22067 17509
rect 24117 17506 24183 17509
rect 19241 17504 24183 17506
rect 19241 17448 19246 17504
rect 19302 17448 22006 17504
rect 22062 17448 24122 17504
rect 24178 17448 24183 17504
rect 19241 17446 24183 17448
rect 19241 17443 19307 17446
rect 22001 17443 22067 17446
rect 24117 17443 24183 17446
rect 24669 17506 24735 17509
rect 27520 17506 28000 17536
rect 24669 17504 28000 17506
rect 24669 17448 24674 17504
rect 24730 17448 28000 17504
rect 24669 17446 28000 17448
rect 24669 17443 24735 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 27520 17416 28000 17446
rect 24277 17375 24597 17376
rect 2589 17234 2655 17237
rect 4705 17234 4771 17237
rect 2589 17232 4771 17234
rect 2589 17176 2594 17232
rect 2650 17176 4710 17232
rect 4766 17176 4771 17232
rect 2589 17174 4771 17176
rect 2589 17171 2655 17174
rect 4705 17171 4771 17174
rect 13537 17234 13603 17237
rect 18505 17234 18571 17237
rect 20713 17234 20779 17237
rect 13537 17232 20779 17234
rect 13537 17176 13542 17232
rect 13598 17176 18510 17232
rect 18566 17176 20718 17232
rect 20774 17176 20779 17232
rect 13537 17174 20779 17176
rect 13537 17171 13603 17174
rect 18505 17171 18571 17174
rect 20713 17171 20779 17174
rect 2773 17098 2839 17101
rect 12341 17098 12407 17101
rect 2773 17096 12407 17098
rect 2773 17040 2778 17096
rect 2834 17040 12346 17096
rect 12402 17040 12407 17096
rect 2773 17038 12407 17040
rect 2773 17035 2839 17038
rect 12341 17035 12407 17038
rect 13261 17098 13327 17101
rect 17769 17098 17835 17101
rect 13261 17096 17835 17098
rect 13261 17040 13266 17096
rect 13322 17040 17774 17096
rect 17830 17040 17835 17096
rect 13261 17038 17835 17040
rect 13261 17035 13327 17038
rect 17769 17035 17835 17038
rect 2037 16962 2103 16965
rect 6085 16962 6151 16965
rect 2037 16960 6151 16962
rect 2037 16904 2042 16960
rect 2098 16904 6090 16960
rect 6146 16904 6151 16960
rect 2037 16902 6151 16904
rect 2037 16899 2103 16902
rect 6085 16899 6151 16902
rect 20805 16962 20871 16965
rect 22461 16962 22527 16965
rect 20805 16960 22527 16962
rect 20805 16904 20810 16960
rect 20866 16904 22466 16960
rect 22522 16904 22527 16960
rect 20805 16902 22527 16904
rect 20805 16899 20871 16902
rect 22461 16899 22527 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 4061 16826 4127 16829
rect 7465 16826 7531 16829
rect 4061 16824 7531 16826
rect 4061 16768 4066 16824
rect 4122 16768 7470 16824
rect 7526 16768 7531 16824
rect 4061 16766 7531 16768
rect 4061 16763 4127 16766
rect 7465 16763 7531 16766
rect 16481 16826 16547 16829
rect 18965 16826 19031 16829
rect 16481 16824 19031 16826
rect 16481 16768 16486 16824
rect 16542 16768 18970 16824
rect 19026 16768 19031 16824
rect 16481 16766 19031 16768
rect 16481 16763 16547 16766
rect 18965 16763 19031 16766
rect 2589 16690 2655 16693
rect 3969 16690 4035 16693
rect 5901 16690 5967 16693
rect 2589 16688 3802 16690
rect 2589 16632 2594 16688
rect 2650 16632 3802 16688
rect 2589 16630 3802 16632
rect 2589 16627 2655 16630
rect 1761 16554 1827 16557
rect 3742 16554 3802 16630
rect 3969 16688 5967 16690
rect 3969 16632 3974 16688
rect 4030 16632 5906 16688
rect 5962 16632 5967 16688
rect 3969 16630 5967 16632
rect 3969 16627 4035 16630
rect 5901 16627 5967 16630
rect 11053 16690 11119 16693
rect 11513 16690 11579 16693
rect 11053 16688 11579 16690
rect 11053 16632 11058 16688
rect 11114 16632 11518 16688
rect 11574 16632 11579 16688
rect 11053 16630 11579 16632
rect 11053 16627 11119 16630
rect 11513 16627 11579 16630
rect 18229 16690 18295 16693
rect 20713 16690 20779 16693
rect 18229 16688 20779 16690
rect 18229 16632 18234 16688
rect 18290 16632 20718 16688
rect 20774 16632 20779 16688
rect 18229 16630 20779 16632
rect 18229 16627 18295 16630
rect 20713 16627 20779 16630
rect 14641 16554 14707 16557
rect 1761 16552 1962 16554
rect 1761 16496 1766 16552
rect 1822 16496 1962 16552
rect 1761 16494 1962 16496
rect 3742 16494 6194 16554
rect 1761 16491 1827 16494
rect 1577 16284 1643 16285
rect 1526 16282 1532 16284
rect 1486 16222 1532 16282
rect 1596 16280 1643 16284
rect 1638 16224 1643 16280
rect 1526 16220 1532 16222
rect 1596 16220 1643 16224
rect 1577 16219 1643 16220
rect 0 16146 480 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 480 16086
rect 1577 16083 1643 16086
rect 1902 16010 1962 16494
rect 6134 16418 6194 16494
rect 14641 16552 15394 16554
rect 14641 16496 14646 16552
rect 14702 16496 15394 16552
rect 14641 16494 15394 16496
rect 14641 16491 14707 16494
rect 10685 16418 10751 16421
rect 6134 16416 10751 16418
rect 6134 16360 10690 16416
rect 10746 16360 10751 16416
rect 6134 16358 10751 16360
rect 15334 16418 15394 16494
rect 20621 16418 20687 16421
rect 15334 16416 20687 16418
rect 15334 16360 20626 16416
rect 20682 16360 20687 16416
rect 15334 16358 20687 16360
rect 10685 16355 10751 16358
rect 20621 16355 20687 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 18781 16282 18847 16285
rect 22093 16282 22159 16285
rect 18781 16280 22159 16282
rect 18781 16224 18786 16280
rect 18842 16224 22098 16280
rect 22154 16224 22159 16280
rect 18781 16222 22159 16224
rect 18781 16219 18847 16222
rect 22093 16219 22159 16222
rect 2037 16146 2103 16149
rect 18873 16146 18939 16149
rect 2037 16144 18939 16146
rect 2037 16088 2042 16144
rect 2098 16088 18878 16144
rect 18934 16088 18939 16144
rect 2037 16086 18939 16088
rect 2037 16083 2103 16086
rect 18873 16083 18939 16086
rect 24761 16146 24827 16149
rect 27520 16146 28000 16176
rect 24761 16144 28000 16146
rect 24761 16088 24766 16144
rect 24822 16088 28000 16144
rect 24761 16086 28000 16088
rect 24761 16083 24827 16086
rect 27520 16056 28000 16086
rect 2037 16010 2103 16013
rect 1902 16008 2103 16010
rect 1902 15952 2042 16008
rect 2098 15952 2103 16008
rect 1902 15950 2103 15952
rect 2037 15947 2103 15950
rect 3693 16010 3759 16013
rect 22921 16010 22987 16013
rect 3693 16008 22987 16010
rect 3693 15952 3698 16008
rect 3754 15952 22926 16008
rect 22982 15952 22987 16008
rect 3693 15950 22987 15952
rect 3693 15947 3759 15950
rect 22921 15947 22987 15950
rect 5257 15874 5323 15877
rect 9305 15874 9371 15877
rect 5257 15872 9371 15874
rect 5257 15816 5262 15872
rect 5318 15816 9310 15872
rect 9366 15816 9371 15872
rect 5257 15814 9371 15816
rect 5257 15811 5323 15814
rect 9305 15811 9371 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 3601 15738 3667 15741
rect 9765 15738 9831 15741
rect 3601 15736 9831 15738
rect 3601 15680 3606 15736
rect 3662 15680 9770 15736
rect 9826 15680 9831 15736
rect 3601 15678 9831 15680
rect 3601 15675 3667 15678
rect 9765 15675 9831 15678
rect 3325 15602 3391 15605
rect 6545 15602 6611 15605
rect 3325 15600 6611 15602
rect 3325 15544 3330 15600
rect 3386 15544 6550 15600
rect 6606 15544 6611 15600
rect 3325 15542 6611 15544
rect 3325 15539 3391 15542
rect 6545 15539 6611 15542
rect 9581 15602 9647 15605
rect 11513 15602 11579 15605
rect 9581 15600 11579 15602
rect 9581 15544 9586 15600
rect 9642 15544 11518 15600
rect 11574 15544 11579 15600
rect 9581 15542 11579 15544
rect 9581 15539 9647 15542
rect 11513 15539 11579 15542
rect 17217 15602 17283 15605
rect 22185 15602 22251 15605
rect 17217 15600 22251 15602
rect 17217 15544 17222 15600
rect 17278 15544 22190 15600
rect 22246 15544 22251 15600
rect 17217 15542 22251 15544
rect 17217 15539 17283 15542
rect 22185 15539 22251 15542
rect 2681 15466 2747 15469
rect 7189 15466 7255 15469
rect 2681 15464 7255 15466
rect 2681 15408 2686 15464
rect 2742 15408 7194 15464
rect 7250 15408 7255 15464
rect 2681 15406 7255 15408
rect 2681 15403 2747 15406
rect 7189 15403 7255 15406
rect 16113 15466 16179 15469
rect 22093 15466 22159 15469
rect 16113 15464 22159 15466
rect 16113 15408 16118 15464
rect 16174 15408 22098 15464
rect 22154 15408 22159 15464
rect 16113 15406 22159 15408
rect 16113 15403 16179 15406
rect 22093 15403 22159 15406
rect 19057 15330 19123 15333
rect 23473 15330 23539 15333
rect 19057 15328 23539 15330
rect 19057 15272 19062 15328
rect 19118 15272 23478 15328
rect 23534 15272 23539 15328
rect 19057 15270 23539 15272
rect 19057 15267 19123 15270
rect 23473 15267 23539 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 10593 15194 10659 15197
rect 12617 15194 12683 15197
rect 10593 15192 12683 15194
rect 10593 15136 10598 15192
rect 10654 15136 12622 15192
rect 12678 15136 12683 15192
rect 10593 15134 12683 15136
rect 10593 15131 10659 15134
rect 12617 15131 12683 15134
rect 16389 15058 16455 15061
rect 24853 15058 24919 15061
rect 16389 15056 24919 15058
rect 16389 15000 16394 15056
rect 16450 15000 24858 15056
rect 24914 15000 24919 15056
rect 16389 14998 24919 15000
rect 16389 14995 16455 14998
rect 24853 14995 24919 14998
rect 3141 14922 3207 14925
rect 4061 14922 4127 14925
rect 21398 14922 21404 14924
rect 3141 14920 21404 14922
rect 3141 14864 3146 14920
rect 3202 14864 4066 14920
rect 4122 14864 21404 14920
rect 3141 14862 21404 14864
rect 3141 14859 3207 14862
rect 4061 14859 4127 14862
rect 21398 14860 21404 14862
rect 21468 14922 21474 14924
rect 23381 14922 23447 14925
rect 24945 14922 25011 14925
rect 21468 14920 25011 14922
rect 21468 14864 23386 14920
rect 23442 14864 24950 14920
rect 25006 14864 25011 14920
rect 21468 14862 25011 14864
rect 21468 14860 21474 14862
rect 23381 14859 23447 14862
rect 24945 14859 25011 14862
rect 0 14786 480 14816
rect 1853 14786 1919 14789
rect 0 14784 1919 14786
rect 0 14728 1858 14784
rect 1914 14728 1919 14784
rect 0 14726 1919 14728
rect 0 14696 480 14726
rect 1853 14723 1919 14726
rect 3141 14786 3207 14789
rect 8661 14786 8727 14789
rect 3141 14784 8727 14786
rect 3141 14728 3146 14784
rect 3202 14728 8666 14784
rect 8722 14728 8727 14784
rect 3141 14726 8727 14728
rect 3141 14723 3207 14726
rect 8661 14723 8727 14726
rect 9806 14724 9812 14788
rect 9876 14786 9882 14788
rect 9949 14786 10015 14789
rect 9876 14784 10015 14786
rect 9876 14728 9954 14784
rect 10010 14728 10015 14784
rect 9876 14726 10015 14728
rect 9876 14724 9882 14726
rect 9949 14723 10015 14726
rect 16941 14786 17007 14789
rect 18597 14786 18663 14789
rect 19333 14786 19399 14789
rect 27520 14786 28000 14816
rect 16941 14784 19399 14786
rect 16941 14728 16946 14784
rect 17002 14728 18602 14784
rect 18658 14728 19338 14784
rect 19394 14728 19399 14784
rect 16941 14726 19399 14728
rect 16941 14723 17007 14726
rect 18597 14723 18663 14726
rect 19333 14723 19399 14726
rect 24902 14726 28000 14786
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 11053 14650 11119 14653
rect 10734 14648 11119 14650
rect 10734 14592 11058 14648
rect 11114 14592 11119 14648
rect 10734 14590 11119 14592
rect 3141 14514 3207 14517
rect 3734 14514 3740 14516
rect 3141 14512 3740 14514
rect 3141 14456 3146 14512
rect 3202 14456 3740 14512
rect 3141 14454 3740 14456
rect 3141 14451 3207 14454
rect 3734 14452 3740 14454
rect 3804 14514 3810 14516
rect 10734 14514 10794 14590
rect 11053 14587 11119 14590
rect 3804 14454 10794 14514
rect 15469 14514 15535 14517
rect 22461 14514 22527 14517
rect 15469 14512 22527 14514
rect 15469 14456 15474 14512
rect 15530 14456 22466 14512
rect 22522 14456 22527 14512
rect 15469 14454 22527 14456
rect 3804 14452 3810 14454
rect 15469 14451 15535 14454
rect 22461 14451 22527 14454
rect 24761 14514 24827 14517
rect 24902 14514 24962 14726
rect 27520 14696 28000 14726
rect 24761 14512 24962 14514
rect 24761 14456 24766 14512
rect 24822 14456 24962 14512
rect 24761 14454 24962 14456
rect 24761 14451 24827 14454
rect 8477 14242 8543 14245
rect 14641 14242 14707 14245
rect 8477 14240 14707 14242
rect 8477 14184 8482 14240
rect 8538 14184 14646 14240
rect 14702 14184 14707 14240
rect 8477 14182 14707 14184
rect 8477 14179 8543 14182
rect 14641 14179 14707 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 6177 14106 6243 14109
rect 8753 14106 8819 14109
rect 11329 14106 11395 14109
rect 6177 14104 11395 14106
rect 6177 14048 6182 14104
rect 6238 14048 8758 14104
rect 8814 14048 11334 14104
rect 11390 14048 11395 14104
rect 6177 14046 11395 14048
rect 6177 14043 6243 14046
rect 8753 14043 8819 14046
rect 11329 14043 11395 14046
rect 5165 13970 5231 13973
rect 10869 13970 10935 13973
rect 12433 13970 12499 13973
rect 5165 13968 9322 13970
rect 5165 13912 5170 13968
rect 5226 13912 9322 13968
rect 5165 13910 9322 13912
rect 5165 13907 5231 13910
rect 9262 13834 9322 13910
rect 10869 13968 12499 13970
rect 10869 13912 10874 13968
rect 10930 13912 12438 13968
rect 12494 13912 12499 13968
rect 10869 13910 12499 13912
rect 10869 13907 10935 13910
rect 12433 13907 12499 13910
rect 13629 13970 13695 13973
rect 15377 13970 15443 13973
rect 13629 13968 15443 13970
rect 13629 13912 13634 13968
rect 13690 13912 15382 13968
rect 15438 13912 15443 13968
rect 13629 13910 15443 13912
rect 13629 13907 13695 13910
rect 15377 13907 15443 13910
rect 11053 13834 11119 13837
rect 9262 13832 11119 13834
rect 9262 13776 11058 13832
rect 11114 13776 11119 13832
rect 9262 13774 11119 13776
rect 11053 13771 11119 13774
rect 11329 13834 11395 13837
rect 12525 13834 12591 13837
rect 11329 13832 12591 13834
rect 11329 13776 11334 13832
rect 11390 13776 12530 13832
rect 12586 13776 12591 13832
rect 11329 13774 12591 13776
rect 11329 13771 11395 13774
rect 12525 13771 12591 13774
rect 15193 13834 15259 13837
rect 23473 13834 23539 13837
rect 15193 13832 23539 13834
rect 15193 13776 15198 13832
rect 15254 13776 23478 13832
rect 23534 13776 23539 13832
rect 15193 13774 23539 13776
rect 15193 13771 15259 13774
rect 23473 13771 23539 13774
rect 23606 13636 23612 13700
rect 23676 13698 23682 13700
rect 24025 13698 24091 13701
rect 23676 13696 24091 13698
rect 23676 13640 24030 13696
rect 24086 13640 24091 13696
rect 23676 13638 24091 13640
rect 23676 13636 23682 13638
rect 24025 13635 24091 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 10869 13562 10935 13565
rect 17125 13562 17191 13565
rect 10869 13560 17191 13562
rect 10869 13504 10874 13560
rect 10930 13504 17130 13560
rect 17186 13504 17191 13560
rect 10869 13502 17191 13504
rect 10869 13499 10935 13502
rect 17125 13499 17191 13502
rect 20161 13562 20227 13565
rect 23473 13562 23539 13565
rect 20161 13560 23539 13562
rect 20161 13504 20166 13560
rect 20222 13504 23478 13560
rect 23534 13504 23539 13560
rect 20161 13502 23539 13504
rect 20161 13499 20227 13502
rect 23473 13499 23539 13502
rect 24025 13562 24091 13565
rect 25129 13562 25195 13565
rect 24025 13560 25195 13562
rect 24025 13504 24030 13560
rect 24086 13504 25134 13560
rect 25190 13504 25195 13560
rect 24025 13502 25195 13504
rect 24025 13499 24091 13502
rect 25129 13499 25195 13502
rect 1761 13426 1827 13429
rect 2865 13426 2931 13429
rect 1761 13424 2931 13426
rect 1761 13368 1766 13424
rect 1822 13368 2870 13424
rect 2926 13368 2931 13424
rect 1761 13366 2931 13368
rect 1761 13363 1827 13366
rect 2865 13363 2931 13366
rect 4981 13426 5047 13429
rect 11697 13426 11763 13429
rect 22829 13426 22895 13429
rect 23197 13426 23263 13429
rect 24209 13426 24275 13429
rect 4981 13424 22754 13426
rect 4981 13368 4986 13424
rect 5042 13368 11702 13424
rect 11758 13368 22754 13424
rect 4981 13366 22754 13368
rect 4981 13363 5047 13366
rect 11697 13363 11763 13366
rect 0 13290 480 13320
rect 4613 13290 4679 13293
rect 8293 13290 8359 13293
rect 0 13230 4032 13290
rect 0 13200 480 13230
rect 3972 12882 4032 13230
rect 4613 13288 8359 13290
rect 4613 13232 4618 13288
rect 4674 13232 8298 13288
rect 8354 13232 8359 13288
rect 4613 13230 8359 13232
rect 4613 13227 4679 13230
rect 8293 13227 8359 13230
rect 9213 13290 9279 13293
rect 10869 13290 10935 13293
rect 9213 13288 10935 13290
rect 9213 13232 9218 13288
rect 9274 13232 10874 13288
rect 10930 13232 10935 13288
rect 9213 13230 10935 13232
rect 9213 13227 9279 13230
rect 10869 13227 10935 13230
rect 11053 13290 11119 13293
rect 18873 13290 18939 13293
rect 21449 13290 21515 13293
rect 11053 13288 18706 13290
rect 11053 13232 11058 13288
rect 11114 13232 18706 13288
rect 11053 13230 18706 13232
rect 11053 13227 11119 13230
rect 7925 13154 7991 13157
rect 11053 13154 11119 13157
rect 7925 13152 11119 13154
rect 7925 13096 7930 13152
rect 7986 13096 11058 13152
rect 11114 13096 11119 13152
rect 7925 13094 11119 13096
rect 7925 13091 7991 13094
rect 11053 13091 11119 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 6637 13018 6703 13021
rect 10317 13018 10383 13021
rect 6637 13016 10383 13018
rect 6637 12960 6642 13016
rect 6698 12960 10322 13016
rect 10378 12960 10383 13016
rect 6637 12958 10383 12960
rect 18646 13018 18706 13230
rect 18873 13288 21515 13290
rect 18873 13232 18878 13288
rect 18934 13232 21454 13288
rect 21510 13232 21515 13288
rect 18873 13230 21515 13232
rect 18873 13227 18939 13230
rect 21449 13227 21515 13230
rect 19190 13092 19196 13156
rect 19260 13154 19266 13156
rect 20437 13154 20503 13157
rect 19260 13152 20503 13154
rect 19260 13096 20442 13152
rect 20498 13096 20503 13152
rect 19260 13094 20503 13096
rect 22694 13154 22754 13366
rect 22829 13424 24275 13426
rect 22829 13368 22834 13424
rect 22890 13368 23202 13424
rect 23258 13368 24214 13424
rect 24270 13368 24275 13424
rect 22829 13366 24275 13368
rect 22829 13363 22895 13366
rect 23197 13363 23263 13366
rect 24209 13363 24275 13366
rect 25589 13290 25655 13293
rect 27520 13290 28000 13320
rect 25589 13288 28000 13290
rect 25589 13232 25594 13288
rect 25650 13232 28000 13288
rect 25589 13230 28000 13232
rect 25589 13227 25655 13230
rect 27520 13200 28000 13230
rect 24025 13154 24091 13157
rect 22694 13152 24091 13154
rect 22694 13096 24030 13152
rect 24086 13096 24091 13152
rect 22694 13094 24091 13096
rect 19260 13092 19266 13094
rect 20437 13091 20503 13094
rect 24025 13091 24091 13094
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 19793 13018 19859 13021
rect 23606 13018 23612 13020
rect 18646 13016 23612 13018
rect 18646 12960 19798 13016
rect 19854 12960 23612 13016
rect 18646 12958 23612 12960
rect 6637 12955 6703 12958
rect 10317 12955 10383 12958
rect 19793 12955 19859 12958
rect 23606 12956 23612 12958
rect 23676 12956 23682 13020
rect 17125 12882 17191 12885
rect 24761 12882 24827 12885
rect 3972 12822 10794 12882
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 2313 12474 2379 12477
rect 3141 12474 3207 12477
rect 2313 12472 3207 12474
rect 2313 12416 2318 12472
rect 2374 12416 3146 12472
rect 3202 12416 3207 12472
rect 2313 12414 3207 12416
rect 2313 12411 2379 12414
rect 3141 12411 3207 12414
rect 6085 12474 6151 12477
rect 10041 12474 10107 12477
rect 6085 12472 10107 12474
rect 6085 12416 6090 12472
rect 6146 12416 10046 12472
rect 10102 12416 10107 12472
rect 6085 12414 10107 12416
rect 10734 12474 10794 12822
rect 17125 12880 24827 12882
rect 17125 12824 17130 12880
rect 17186 12824 24766 12880
rect 24822 12824 24827 12880
rect 17125 12822 24827 12824
rect 17125 12819 17191 12822
rect 24761 12819 24827 12822
rect 16389 12746 16455 12749
rect 24945 12746 25011 12749
rect 16389 12744 25011 12746
rect 16389 12688 16394 12744
rect 16450 12688 24950 12744
rect 25006 12688 25011 12744
rect 16389 12686 25011 12688
rect 16389 12683 16455 12686
rect 24945 12683 25011 12686
rect 12341 12610 12407 12613
rect 14549 12610 14615 12613
rect 12341 12608 14615 12610
rect 12341 12552 12346 12608
rect 12402 12552 14554 12608
rect 14610 12552 14615 12608
rect 12341 12550 14615 12552
rect 12341 12547 12407 12550
rect 14549 12547 14615 12550
rect 15469 12610 15535 12613
rect 17217 12610 17283 12613
rect 15469 12608 17283 12610
rect 15469 12552 15474 12608
rect 15530 12552 17222 12608
rect 17278 12552 17283 12608
rect 15469 12550 17283 12552
rect 15469 12547 15535 12550
rect 17217 12547 17283 12550
rect 18321 12610 18387 12613
rect 18597 12610 18663 12613
rect 18321 12608 18663 12610
rect 18321 12552 18326 12608
rect 18382 12552 18602 12608
rect 18658 12552 18663 12608
rect 18321 12550 18663 12552
rect 18321 12547 18387 12550
rect 18597 12547 18663 12550
rect 23657 12610 23723 12613
rect 24025 12610 24091 12613
rect 23657 12608 24091 12610
rect 23657 12552 23662 12608
rect 23718 12552 24030 12608
rect 24086 12552 24091 12608
rect 23657 12550 24091 12552
rect 23657 12547 23723 12550
rect 24025 12547 24091 12550
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 10734 12414 19442 12474
rect 6085 12411 6151 12414
rect 10041 12411 10107 12414
rect 3325 12338 3391 12341
rect 12433 12338 12499 12341
rect 3325 12336 12499 12338
rect 3325 12280 3330 12336
rect 3386 12280 12438 12336
rect 12494 12280 12499 12336
rect 3325 12278 12499 12280
rect 19382 12338 19442 12414
rect 19517 12338 19583 12341
rect 22461 12338 22527 12341
rect 19382 12336 22527 12338
rect 19382 12280 19522 12336
rect 19578 12280 22466 12336
rect 22522 12280 22527 12336
rect 19382 12278 22527 12280
rect 3325 12275 3391 12278
rect 12433 12275 12499 12278
rect 19517 12275 19583 12278
rect 22461 12275 22527 12278
rect 2865 12202 2931 12205
rect 9806 12202 9812 12204
rect 2865 12200 9812 12202
rect 2865 12144 2870 12200
rect 2926 12144 9812 12200
rect 2865 12142 9812 12144
rect 2865 12139 2931 12142
rect 9806 12140 9812 12142
rect 9876 12202 9882 12204
rect 11237 12202 11303 12205
rect 12985 12202 13051 12205
rect 9876 12200 13051 12202
rect 9876 12144 11242 12200
rect 11298 12144 12990 12200
rect 13046 12144 13051 12200
rect 9876 12142 13051 12144
rect 9876 12140 9882 12142
rect 11237 12139 11303 12142
rect 12985 12139 13051 12142
rect 14181 12202 14247 12205
rect 18965 12202 19031 12205
rect 14181 12200 19031 12202
rect 14181 12144 14186 12200
rect 14242 12144 18970 12200
rect 19026 12144 19031 12200
rect 14181 12142 19031 12144
rect 14181 12139 14247 12142
rect 18965 12139 19031 12142
rect 19333 12202 19399 12205
rect 22277 12202 22343 12205
rect 19333 12200 22343 12202
rect 19333 12144 19338 12200
rect 19394 12144 22282 12200
rect 22338 12144 22343 12200
rect 19333 12142 22343 12144
rect 19333 12139 19399 12142
rect 22277 12139 22343 12142
rect 24025 12202 24091 12205
rect 25405 12202 25471 12205
rect 24025 12200 25471 12202
rect 24025 12144 24030 12200
rect 24086 12144 25410 12200
rect 25466 12144 25471 12200
rect 24025 12142 25471 12144
rect 24025 12139 24091 12142
rect 25405 12139 25471 12142
rect 8845 12066 8911 12069
rect 12709 12066 12775 12069
rect 22185 12066 22251 12069
rect 6180 12064 12775 12066
rect 6180 12008 8850 12064
rect 8906 12008 12714 12064
rect 12770 12008 12775 12064
rect 6180 12006 12775 12008
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 0 11870 5458 11930
rect 0 11840 480 11870
rect 5398 11794 5458 11870
rect 6180 11794 6240 12006
rect 8845 12003 8911 12006
rect 12709 12003 12775 12006
rect 16990 12064 22251 12066
rect 16990 12008 22190 12064
rect 22246 12008 22251 12064
rect 16990 12006 22251 12008
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 5398 11734 6240 11794
rect 8937 11794 9003 11797
rect 11421 11794 11487 11797
rect 16990 11794 17050 12006
rect 22185 12003 22251 12006
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 21265 11930 21331 11933
rect 21398 11930 21404 11932
rect 21265 11928 21404 11930
rect 21265 11872 21270 11928
rect 21326 11872 21404 11928
rect 21265 11870 21404 11872
rect 21265 11867 21331 11870
rect 21398 11868 21404 11870
rect 21468 11868 21474 11932
rect 27520 11930 28000 11960
rect 24902 11870 28000 11930
rect 24902 11794 24962 11870
rect 27520 11840 28000 11870
rect 8937 11792 11346 11794
rect 8937 11736 8942 11792
rect 8998 11736 11346 11792
rect 8937 11734 11346 11736
rect 8937 11731 9003 11734
rect 5073 11658 5139 11661
rect 11053 11658 11119 11661
rect 5073 11656 11119 11658
rect 5073 11600 5078 11656
rect 5134 11600 11058 11656
rect 11114 11600 11119 11656
rect 5073 11598 11119 11600
rect 11286 11658 11346 11734
rect 11421 11792 17050 11794
rect 11421 11736 11426 11792
rect 11482 11736 17050 11792
rect 11421 11734 17050 11736
rect 17220 11734 24962 11794
rect 11421 11731 11487 11734
rect 11513 11658 11579 11661
rect 17033 11658 17099 11661
rect 11286 11656 17099 11658
rect 11286 11600 11518 11656
rect 11574 11600 17038 11656
rect 17094 11600 17099 11656
rect 11286 11598 17099 11600
rect 5073 11595 5139 11598
rect 11053 11595 11119 11598
rect 11513 11595 11579 11598
rect 17033 11595 17099 11598
rect 2313 11522 2379 11525
rect 7005 11522 7071 11525
rect 2313 11520 7071 11522
rect 2313 11464 2318 11520
rect 2374 11464 7010 11520
rect 7066 11464 7071 11520
rect 2313 11462 7071 11464
rect 2313 11459 2379 11462
rect 7005 11459 7071 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 12065 11386 12131 11389
rect 17220 11386 17280 11734
rect 18873 11658 18939 11661
rect 23749 11658 23815 11661
rect 18873 11656 23815 11658
rect 18873 11600 18878 11656
rect 18934 11600 23754 11656
rect 23810 11600 23815 11656
rect 18873 11598 23815 11600
rect 18873 11595 18939 11598
rect 23749 11595 23815 11598
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 12065 11384 17280 11386
rect 12065 11328 12070 11384
rect 12126 11328 17280 11384
rect 12065 11326 17280 11328
rect 22185 11386 22251 11389
rect 22461 11386 22527 11389
rect 22185 11384 22527 11386
rect 22185 11328 22190 11384
rect 22246 11328 22466 11384
rect 22522 11328 22527 11384
rect 22185 11326 22527 11328
rect 12065 11323 12131 11326
rect 22185 11323 22251 11326
rect 22461 11323 22527 11326
rect 1577 11250 1643 11253
rect 2865 11250 2931 11253
rect 1577 11248 2931 11250
rect 1577 11192 1582 11248
rect 1638 11192 2870 11248
rect 2926 11192 2931 11248
rect 1577 11190 2931 11192
rect 1577 11187 1643 11190
rect 2865 11187 2931 11190
rect 4705 11250 4771 11253
rect 11421 11250 11487 11253
rect 4705 11248 11487 11250
rect 4705 11192 4710 11248
rect 4766 11192 11426 11248
rect 11482 11192 11487 11248
rect 4705 11190 11487 11192
rect 4705 11187 4771 11190
rect 11421 11187 11487 11190
rect 17309 11250 17375 11253
rect 24945 11250 25011 11253
rect 17309 11248 25011 11250
rect 17309 11192 17314 11248
rect 17370 11192 24950 11248
rect 25006 11192 25011 11248
rect 17309 11190 25011 11192
rect 17309 11187 17375 11190
rect 24945 11187 25011 11190
rect 12801 11114 12867 11117
rect 15837 11114 15903 11117
rect 12801 11112 15903 11114
rect 12801 11056 12806 11112
rect 12862 11056 15842 11112
rect 15898 11056 15903 11112
rect 12801 11054 15903 11056
rect 12801 11051 12867 11054
rect 15837 11051 15903 11054
rect 17677 11114 17743 11117
rect 20161 11114 20227 11117
rect 17677 11112 20227 11114
rect 17677 11056 17682 11112
rect 17738 11056 20166 11112
rect 20222 11056 20227 11112
rect 17677 11054 20227 11056
rect 17677 11051 17743 11054
rect 20161 11051 20227 11054
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 2129 10706 2195 10709
rect 7833 10706 7899 10709
rect 2129 10704 7899 10706
rect 2129 10648 2134 10704
rect 2190 10648 7838 10704
rect 7894 10648 7899 10704
rect 2129 10646 7899 10648
rect 2129 10643 2195 10646
rect 7833 10643 7899 10646
rect 8477 10706 8543 10709
rect 10777 10706 10843 10709
rect 8477 10704 10843 10706
rect 8477 10648 8482 10704
rect 8538 10648 10782 10704
rect 10838 10648 10843 10704
rect 8477 10646 10843 10648
rect 8477 10643 8543 10646
rect 10777 10643 10843 10646
rect 14089 10706 14155 10709
rect 18137 10706 18203 10709
rect 14089 10704 18203 10706
rect 14089 10648 14094 10704
rect 14150 10648 18142 10704
rect 18198 10648 18203 10704
rect 14089 10646 18203 10648
rect 14089 10643 14155 10646
rect 18137 10643 18203 10646
rect 0 10570 480 10600
rect 22829 10570 22895 10573
rect 27520 10570 28000 10600
rect 0 10510 10794 10570
rect 0 10480 480 10510
rect 5257 10434 5323 10437
rect 9673 10434 9739 10437
rect 5257 10432 9739 10434
rect 5257 10376 5262 10432
rect 5318 10376 9678 10432
rect 9734 10376 9739 10432
rect 5257 10374 9739 10376
rect 10734 10434 10794 10510
rect 15702 10568 22895 10570
rect 15702 10512 22834 10568
rect 22890 10512 22895 10568
rect 15702 10510 22895 10512
rect 14641 10434 14707 10437
rect 15702 10434 15762 10510
rect 22829 10507 22895 10510
rect 24902 10510 28000 10570
rect 10734 10432 15762 10434
rect 10734 10376 14646 10432
rect 14702 10376 15762 10432
rect 10734 10374 15762 10376
rect 21081 10434 21147 10437
rect 23749 10434 23815 10437
rect 21081 10432 23815 10434
rect 21081 10376 21086 10432
rect 21142 10376 23754 10432
rect 23810 10376 23815 10432
rect 21081 10374 23815 10376
rect 5257 10371 5323 10374
rect 9673 10371 9739 10374
rect 14641 10371 14707 10374
rect 21081 10371 21147 10374
rect 23749 10371 23815 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 5993 10298 6059 10301
rect 6913 10298 6979 10301
rect 5993 10296 10104 10298
rect 5993 10240 5998 10296
rect 6054 10240 6918 10296
rect 6974 10240 10104 10296
rect 5993 10238 10104 10240
rect 5993 10235 6059 10238
rect 6913 10235 6979 10238
rect 10044 10162 10104 10238
rect 12065 10162 12131 10165
rect 10044 10160 12131 10162
rect 10044 10104 12070 10160
rect 12126 10104 12131 10160
rect 10044 10102 12131 10104
rect 12065 10099 12131 10102
rect 12709 10162 12775 10165
rect 21909 10162 21975 10165
rect 24902 10162 24962 10510
rect 27520 10480 28000 10510
rect 12709 10160 24962 10162
rect 12709 10104 12714 10160
rect 12770 10104 21914 10160
rect 21970 10104 24962 10160
rect 12709 10102 24962 10104
rect 12709 10099 12775 10102
rect 21909 10099 21975 10102
rect 2773 10026 2839 10029
rect 3182 10026 3188 10028
rect 2773 10024 3188 10026
rect 2773 9968 2778 10024
rect 2834 9968 3188 10024
rect 2773 9966 3188 9968
rect 2773 9963 2839 9966
rect 3182 9964 3188 9966
rect 3252 9964 3258 10028
rect 6821 10026 6887 10029
rect 5398 10024 6887 10026
rect 5398 9968 6826 10024
rect 6882 9968 6887 10024
rect 5398 9966 6887 9968
rect 2313 9890 2379 9893
rect 5257 9890 5323 9893
rect 5398 9890 5458 9966
rect 6821 9963 6887 9966
rect 24117 10024 24183 10029
rect 24117 9968 24122 10024
rect 24178 9968 24183 10024
rect 24117 9963 24183 9968
rect 2313 9888 5458 9890
rect 2313 9832 2318 9888
rect 2374 9832 5262 9888
rect 5318 9832 5458 9888
rect 2313 9830 5458 9832
rect 2313 9827 2379 9830
rect 5257 9827 5323 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 1577 9754 1643 9757
rect 2773 9754 2839 9757
rect 1577 9752 2839 9754
rect 1577 9696 1582 9752
rect 1638 9696 2778 9752
rect 2834 9696 2839 9752
rect 1577 9694 2839 9696
rect 1577 9691 1643 9694
rect 2773 9691 2839 9694
rect 18873 9754 18939 9757
rect 23013 9754 23079 9757
rect 23289 9754 23355 9757
rect 18873 9752 23355 9754
rect 18873 9696 18878 9752
rect 18934 9696 23018 9752
rect 23074 9696 23294 9752
rect 23350 9696 23355 9752
rect 24120 9723 24180 9963
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 18873 9694 23355 9696
rect 18873 9691 18939 9694
rect 23013 9691 23079 9694
rect 23289 9691 23355 9694
rect 24117 9718 24183 9723
rect 24117 9662 24122 9718
rect 24178 9662 24183 9718
rect 24117 9657 24183 9662
rect 7281 9618 7347 9621
rect 11881 9618 11947 9621
rect 20713 9618 20779 9621
rect 7281 9616 11947 9618
rect 7281 9560 7286 9616
rect 7342 9560 11886 9616
rect 11942 9560 11947 9616
rect 7281 9558 11947 9560
rect 7281 9555 7347 9558
rect 11881 9555 11947 9558
rect 15150 9616 20779 9618
rect 15150 9560 20718 9616
rect 20774 9560 20779 9616
rect 15150 9558 20779 9560
rect 1853 9482 1919 9485
rect 10225 9482 10291 9485
rect 1853 9480 10291 9482
rect 1853 9424 1858 9480
rect 1914 9424 10230 9480
rect 10286 9424 10291 9480
rect 1853 9422 10291 9424
rect 1853 9419 1919 9422
rect 10225 9419 10291 9422
rect 12525 9482 12591 9485
rect 15150 9482 15210 9558
rect 20713 9555 20779 9558
rect 12525 9480 15210 9482
rect 12525 9424 12530 9480
rect 12586 9424 15210 9480
rect 12525 9422 15210 9424
rect 15377 9482 15443 9485
rect 17401 9482 17467 9485
rect 15377 9480 17467 9482
rect 15377 9424 15382 9480
rect 15438 9424 17406 9480
rect 17462 9424 17467 9480
rect 15377 9422 17467 9424
rect 12525 9419 12591 9422
rect 15377 9419 15443 9422
rect 17401 9419 17467 9422
rect 17861 9482 17927 9485
rect 20529 9482 20595 9485
rect 25221 9482 25287 9485
rect 17861 9480 20178 9482
rect 17861 9424 17866 9480
rect 17922 9424 20178 9480
rect 17861 9422 20178 9424
rect 17861 9419 17927 9422
rect 20118 9349 20178 9422
rect 20529 9480 25287 9482
rect 20529 9424 20534 9480
rect 20590 9424 25226 9480
rect 25282 9424 25287 9480
rect 20529 9422 25287 9424
rect 20529 9419 20595 9422
rect 25221 9419 25287 9422
rect 3325 9346 3391 9349
rect 9765 9346 9831 9349
rect 3325 9344 9831 9346
rect 3325 9288 3330 9344
rect 3386 9288 9770 9344
rect 9826 9288 9831 9344
rect 3325 9286 9831 9288
rect 3325 9283 3391 9286
rect 9765 9283 9831 9286
rect 20069 9346 20178 9349
rect 23013 9346 23079 9349
rect 20069 9344 23079 9346
rect 20069 9288 20074 9344
rect 20130 9288 23018 9344
rect 23074 9288 23079 9344
rect 20069 9286 23079 9288
rect 20069 9283 20135 9286
rect 23013 9283 23079 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 2405 9210 2471 9213
rect 7281 9210 7347 9213
rect 14365 9210 14431 9213
rect 1166 9150 1548 9210
rect 0 9074 480 9104
rect 1166 9077 1226 9150
rect 1166 9074 1275 9077
rect 1488 9074 1548 9150
rect 2405 9208 7347 9210
rect 2405 9152 2410 9208
rect 2466 9152 7286 9208
rect 7342 9152 7347 9208
rect 2405 9150 7347 9152
rect 2405 9147 2471 9150
rect 7281 9147 7347 9150
rect 11976 9208 14431 9210
rect 11976 9152 14370 9208
rect 14426 9152 14431 9208
rect 11976 9150 14431 9152
rect 11976 9074 12036 9150
rect 14365 9147 14431 9150
rect 24761 9210 24827 9213
rect 24761 9208 25146 9210
rect 24761 9152 24766 9208
rect 24822 9152 25146 9208
rect 24761 9150 25146 9152
rect 24761 9147 24827 9150
rect 0 9072 1356 9074
rect 0 9016 1214 9072
rect 1270 9016 1356 9072
rect 0 9014 1356 9016
rect 1488 9014 12036 9074
rect 13721 9074 13787 9077
rect 24853 9074 24919 9077
rect 13721 9072 24919 9074
rect 13721 9016 13726 9072
rect 13782 9016 24858 9072
rect 24914 9016 24919 9072
rect 13721 9014 24919 9016
rect 25086 9074 25146 9150
rect 27520 9074 28000 9104
rect 25086 9014 28000 9074
rect 0 8984 480 9014
rect 1209 9011 1275 9014
rect 13721 9011 13787 9014
rect 24853 9011 24919 9014
rect 27520 8984 28000 9014
rect 9213 8938 9279 8941
rect 10041 8938 10107 8941
rect 13353 8938 13419 8941
rect 9213 8936 13419 8938
rect 9213 8880 9218 8936
rect 9274 8880 10046 8936
rect 10102 8880 13358 8936
rect 13414 8880 13419 8936
rect 9213 8878 13419 8880
rect 9213 8875 9279 8878
rect 10041 8875 10107 8878
rect 13353 8875 13419 8878
rect 14089 8938 14155 8941
rect 24853 8938 24919 8941
rect 14089 8936 24919 8938
rect 14089 8880 14094 8936
rect 14150 8880 24858 8936
rect 24914 8880 24919 8936
rect 14089 8878 24919 8880
rect 14089 8875 14155 8878
rect 24853 8875 24919 8878
rect 11605 8802 11671 8805
rect 13905 8802 13971 8805
rect 11605 8800 13971 8802
rect 11605 8744 11610 8800
rect 11666 8744 13910 8800
rect 13966 8744 13971 8800
rect 11605 8742 13971 8744
rect 11605 8739 11671 8742
rect 13905 8739 13971 8742
rect 16205 8802 16271 8805
rect 18045 8802 18111 8805
rect 19793 8802 19859 8805
rect 23197 8802 23263 8805
rect 16205 8800 23263 8802
rect 16205 8744 16210 8800
rect 16266 8744 18050 8800
rect 18106 8744 19798 8800
rect 19854 8744 23202 8800
rect 23258 8744 23263 8800
rect 16205 8742 23263 8744
rect 16205 8739 16271 8742
rect 18045 8739 18111 8742
rect 19793 8739 19859 8742
rect 23197 8739 23263 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 18689 8666 18755 8669
rect 20529 8666 20595 8669
rect 18689 8664 20595 8666
rect 18689 8608 18694 8664
rect 18750 8608 20534 8664
rect 20590 8608 20595 8664
rect 18689 8606 20595 8608
rect 18689 8603 18755 8606
rect 20529 8603 20595 8606
rect 3877 8530 3943 8533
rect 6361 8530 6427 8533
rect 3877 8528 6427 8530
rect 3877 8472 3882 8528
rect 3938 8472 6366 8528
rect 6422 8472 6427 8528
rect 3877 8470 6427 8472
rect 3877 8467 3943 8470
rect 6361 8467 6427 8470
rect 6545 8530 6611 8533
rect 21541 8530 21607 8533
rect 25037 8530 25103 8533
rect 6545 8528 25103 8530
rect 6545 8472 6550 8528
rect 6606 8472 21546 8528
rect 21602 8472 25042 8528
rect 25098 8472 25103 8528
rect 6545 8470 25103 8472
rect 6545 8467 6611 8470
rect 21541 8467 21607 8470
rect 25037 8467 25103 8470
rect 3141 8394 3207 8397
rect 5809 8394 5875 8397
rect 3141 8392 5875 8394
rect 3141 8336 3146 8392
rect 3202 8336 5814 8392
rect 5870 8336 5875 8392
rect 3141 8334 5875 8336
rect 3141 8331 3207 8334
rect 5809 8331 5875 8334
rect 13629 8394 13695 8397
rect 25129 8394 25195 8397
rect 13629 8392 25195 8394
rect 13629 8336 13634 8392
rect 13690 8336 25134 8392
rect 25190 8336 25195 8392
rect 13629 8334 25195 8336
rect 13629 8331 13695 8334
rect 25129 8331 25195 8334
rect 5441 8258 5507 8261
rect 9581 8258 9647 8261
rect 5441 8256 9647 8258
rect 5441 8200 5446 8256
rect 5502 8200 9586 8256
rect 9642 8200 9647 8256
rect 5441 8198 9647 8200
rect 5441 8195 5507 8198
rect 9581 8195 9647 8198
rect 10869 8258 10935 8261
rect 18321 8258 18387 8261
rect 10869 8256 18387 8258
rect 10869 8200 10874 8256
rect 10930 8200 18326 8256
rect 18382 8200 18387 8256
rect 10869 8198 18387 8200
rect 10869 8195 10935 8198
rect 18321 8195 18387 8198
rect 21817 8258 21883 8261
rect 23749 8258 23815 8261
rect 21817 8256 23815 8258
rect 21817 8200 21822 8256
rect 21878 8200 23754 8256
rect 23810 8200 23815 8256
rect 21817 8198 23815 8200
rect 21817 8195 21883 8198
rect 23749 8195 23815 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 20069 8122 20135 8125
rect 20437 8122 20503 8125
rect 24761 8122 24827 8125
rect 20069 8120 24827 8122
rect 20069 8064 20074 8120
rect 20130 8064 20442 8120
rect 20498 8064 24766 8120
rect 24822 8064 24827 8120
rect 20069 8062 24827 8064
rect 20069 8059 20135 8062
rect 20437 8059 20503 8062
rect 24761 8059 24827 8062
rect 3233 7986 3299 7989
rect 4153 7986 4219 7989
rect 3233 7984 4219 7986
rect 3233 7928 3238 7984
rect 3294 7928 4158 7984
rect 4214 7928 4219 7984
rect 3233 7926 4219 7928
rect 3233 7923 3299 7926
rect 4153 7923 4219 7926
rect 8753 7986 8819 7989
rect 12985 7986 13051 7989
rect 8753 7984 13051 7986
rect 8753 7928 8758 7984
rect 8814 7928 12990 7984
rect 13046 7928 13051 7984
rect 8753 7926 13051 7928
rect 8753 7923 8819 7926
rect 12985 7923 13051 7926
rect 13721 7986 13787 7989
rect 25129 7986 25195 7989
rect 13721 7984 25195 7986
rect 13721 7928 13726 7984
rect 13782 7928 25134 7984
rect 25190 7928 25195 7984
rect 13721 7926 25195 7928
rect 13721 7923 13787 7926
rect 25129 7923 25195 7926
rect 1117 7850 1183 7853
rect 1526 7850 1532 7852
rect 1117 7848 1532 7850
rect 1117 7792 1122 7848
rect 1178 7792 1532 7848
rect 1117 7790 1532 7792
rect 1117 7787 1183 7790
rect 1526 7788 1532 7790
rect 1596 7850 1602 7852
rect 6545 7850 6611 7853
rect 8293 7850 8359 7853
rect 1596 7790 6056 7850
rect 1596 7788 1602 7790
rect 0 7714 480 7744
rect 4981 7714 5047 7717
rect 0 7712 5047 7714
rect 0 7656 4986 7712
rect 5042 7656 5047 7712
rect 0 7654 5047 7656
rect 5996 7714 6056 7790
rect 6545 7848 8359 7850
rect 6545 7792 6550 7848
rect 6606 7792 8298 7848
rect 8354 7792 8359 7848
rect 6545 7790 8359 7792
rect 6545 7787 6611 7790
rect 8293 7787 8359 7790
rect 8753 7850 8819 7853
rect 18873 7850 18939 7853
rect 8753 7848 18939 7850
rect 8753 7792 8758 7848
rect 8814 7792 18878 7848
rect 18934 7792 18939 7848
rect 8753 7790 18939 7792
rect 8753 7787 8819 7790
rect 18873 7787 18939 7790
rect 20621 7850 20687 7853
rect 24945 7850 25011 7853
rect 20621 7848 25011 7850
rect 20621 7792 20626 7848
rect 20682 7792 24950 7848
rect 25006 7792 25011 7848
rect 20621 7790 25011 7792
rect 20621 7787 20687 7790
rect 24945 7787 25011 7790
rect 12801 7714 12867 7717
rect 5996 7712 12867 7714
rect 5996 7656 12806 7712
rect 12862 7656 12867 7712
rect 5996 7654 12867 7656
rect 0 7624 480 7654
rect 4981 7651 5047 7654
rect 12801 7651 12867 7654
rect 15377 7714 15443 7717
rect 20069 7714 20135 7717
rect 15377 7712 20135 7714
rect 15377 7656 15382 7712
rect 15438 7656 20074 7712
rect 20130 7656 20135 7712
rect 15377 7654 20135 7656
rect 15377 7651 15443 7654
rect 20069 7651 20135 7654
rect 20253 7714 20319 7717
rect 23473 7714 23539 7717
rect 27520 7714 28000 7744
rect 20253 7712 23539 7714
rect 20253 7656 20258 7712
rect 20314 7656 23478 7712
rect 23534 7656 23539 7712
rect 20253 7654 23539 7656
rect 20253 7651 20319 7654
rect 23473 7651 23539 7654
rect 24902 7654 28000 7714
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 16021 7578 16087 7581
rect 16021 7576 20914 7578
rect 16021 7520 16026 7576
rect 16082 7520 20914 7576
rect 16021 7518 20914 7520
rect 16021 7515 16087 7518
rect 1761 7442 1827 7445
rect 8293 7442 8359 7445
rect 1761 7440 8359 7442
rect 1761 7384 1766 7440
rect 1822 7384 8298 7440
rect 8354 7384 8359 7440
rect 1761 7382 8359 7384
rect 1761 7379 1827 7382
rect 8293 7379 8359 7382
rect 9397 7442 9463 7445
rect 13169 7442 13235 7445
rect 13997 7442 14063 7445
rect 9397 7440 14063 7442
rect 9397 7384 9402 7440
rect 9458 7384 13174 7440
rect 13230 7384 14002 7440
rect 14058 7384 14063 7440
rect 9397 7382 14063 7384
rect 9397 7379 9463 7382
rect 13169 7379 13235 7382
rect 13997 7379 14063 7382
rect 14457 7442 14523 7445
rect 20713 7442 20779 7445
rect 14457 7440 20779 7442
rect 14457 7384 14462 7440
rect 14518 7384 20718 7440
rect 20774 7384 20779 7440
rect 14457 7382 20779 7384
rect 14457 7379 14523 7382
rect 20713 7379 20779 7382
rect 3141 7308 3207 7309
rect 3141 7306 3188 7308
rect 3096 7304 3188 7306
rect 3252 7306 3258 7308
rect 6913 7306 6979 7309
rect 3252 7304 6979 7306
rect 3096 7248 3146 7304
rect 3252 7248 6918 7304
rect 6974 7248 6979 7304
rect 3096 7246 3188 7248
rect 3141 7244 3188 7246
rect 3252 7246 6979 7248
rect 3252 7244 3258 7246
rect 3141 7243 3207 7244
rect 6913 7243 6979 7246
rect 7097 7306 7163 7309
rect 12893 7306 12959 7309
rect 15561 7306 15627 7309
rect 20854 7306 20914 7518
rect 21449 7442 21515 7445
rect 21909 7442 21975 7445
rect 24577 7442 24643 7445
rect 21449 7440 24643 7442
rect 21449 7384 21454 7440
rect 21510 7384 21914 7440
rect 21970 7384 24582 7440
rect 24638 7384 24643 7440
rect 21449 7382 24643 7384
rect 21449 7379 21515 7382
rect 21909 7379 21975 7382
rect 24577 7379 24643 7382
rect 24902 7306 24962 7654
rect 27520 7624 28000 7654
rect 7097 7304 10794 7306
rect 7097 7248 7102 7304
rect 7158 7248 10794 7304
rect 7097 7246 10794 7248
rect 7097 7243 7163 7246
rect 2497 7170 2563 7173
rect 7189 7170 7255 7173
rect 8201 7170 8267 7173
rect 2497 7168 8267 7170
rect 2497 7112 2502 7168
rect 2558 7112 7194 7168
rect 7250 7112 8206 7168
rect 8262 7112 8267 7168
rect 2497 7110 8267 7112
rect 2497 7107 2563 7110
rect 7189 7107 7255 7110
rect 8201 7107 8267 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 6085 7034 6151 7037
rect 8385 7034 8451 7037
rect 6085 7032 8451 7034
rect 6085 6976 6090 7032
rect 6146 6976 8390 7032
rect 8446 6976 8451 7032
rect 6085 6974 8451 6976
rect 10734 7034 10794 7246
rect 11102 7304 15627 7306
rect 11102 7248 12898 7304
rect 12954 7248 15566 7304
rect 15622 7248 15627 7304
rect 11102 7246 15627 7248
rect 11102 7173 11162 7246
rect 12893 7243 12959 7246
rect 15561 7243 15627 7246
rect 19382 7246 20178 7306
rect 20854 7246 24962 7306
rect 11053 7168 11162 7173
rect 11053 7112 11058 7168
rect 11114 7112 11162 7168
rect 11053 7110 11162 7112
rect 12157 7170 12223 7173
rect 19382 7170 19442 7246
rect 12157 7168 19442 7170
rect 12157 7112 12162 7168
rect 12218 7112 19442 7168
rect 12157 7110 19442 7112
rect 20118 7170 20178 7246
rect 21173 7170 21239 7173
rect 22277 7170 22343 7173
rect 23473 7170 23539 7173
rect 20118 7168 23539 7170
rect 20118 7112 21178 7168
rect 21234 7112 22282 7168
rect 22338 7112 23478 7168
rect 23534 7112 23539 7168
rect 20118 7110 23539 7112
rect 11053 7107 11119 7110
rect 12157 7107 12223 7110
rect 21173 7107 21239 7110
rect 22277 7107 22343 7110
rect 23473 7107 23539 7110
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 15009 7034 15075 7037
rect 10734 7032 15075 7034
rect 10734 6976 15014 7032
rect 15070 6976 15075 7032
rect 10734 6974 15075 6976
rect 6085 6971 6151 6974
rect 8385 6971 8451 6974
rect 15009 6971 15075 6974
rect 2957 6900 3023 6901
rect 2957 6896 3004 6900
rect 3068 6898 3074 6900
rect 7281 6898 7347 6901
rect 8569 6898 8635 6901
rect 2957 6840 2962 6896
rect 2957 6836 3004 6840
rect 3068 6838 3114 6898
rect 7281 6896 8635 6898
rect 7281 6840 7286 6896
rect 7342 6840 8574 6896
rect 8630 6840 8635 6896
rect 7281 6838 8635 6840
rect 3068 6836 3074 6838
rect 2957 6835 3023 6836
rect 7281 6835 7347 6838
rect 8569 6835 8635 6838
rect 12065 6898 12131 6901
rect 16849 6898 16915 6901
rect 12065 6896 16915 6898
rect 12065 6840 12070 6896
rect 12126 6840 16854 6896
rect 16910 6840 16915 6896
rect 12065 6838 16915 6840
rect 12065 6835 12131 6838
rect 16849 6835 16915 6838
rect 24209 6898 24275 6901
rect 25497 6898 25563 6901
rect 24209 6896 25563 6898
rect 24209 6840 24214 6896
rect 24270 6840 25502 6896
rect 25558 6840 25563 6896
rect 24209 6838 25563 6840
rect 24209 6835 24275 6838
rect 25497 6835 25563 6838
rect 1853 6762 1919 6765
rect 8845 6762 8911 6765
rect 1853 6760 8911 6762
rect 1853 6704 1858 6760
rect 1914 6704 8850 6760
rect 8906 6704 8911 6760
rect 1853 6702 8911 6704
rect 1853 6699 1919 6702
rect 8845 6699 8911 6702
rect 15285 6762 15351 6765
rect 17585 6762 17651 6765
rect 20253 6762 20319 6765
rect 15285 6760 20319 6762
rect 15285 6704 15290 6760
rect 15346 6704 17590 6760
rect 17646 6704 20258 6760
rect 20314 6704 20319 6760
rect 15285 6702 20319 6704
rect 15285 6699 15351 6702
rect 17585 6699 17651 6702
rect 20253 6699 20319 6702
rect 16481 6626 16547 6629
rect 23381 6626 23447 6629
rect 16481 6624 23447 6626
rect 16481 6568 16486 6624
rect 16542 6568 23386 6624
rect 23442 6568 23447 6624
rect 16481 6566 23447 6568
rect 16481 6563 16547 6566
rect 23381 6563 23447 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 3734 6490 3740 6492
rect 1350 6430 3740 6490
rect 0 6354 480 6384
rect 1350 6354 1410 6430
rect 3734 6428 3740 6430
rect 3804 6428 3810 6492
rect 15837 6490 15903 6493
rect 20069 6490 20135 6493
rect 15334 6488 20135 6490
rect 15334 6432 15842 6488
rect 15898 6432 20074 6488
rect 20130 6432 20135 6488
rect 15334 6430 20135 6432
rect 0 6294 1410 6354
rect 1761 6354 1827 6357
rect 4889 6354 4955 6357
rect 7281 6354 7347 6357
rect 1761 6352 7347 6354
rect 1761 6296 1766 6352
rect 1822 6296 4894 6352
rect 4950 6296 7286 6352
rect 7342 6296 7347 6352
rect 1761 6294 7347 6296
rect 0 6264 480 6294
rect 1761 6291 1827 6294
rect 4889 6291 4955 6294
rect 7281 6291 7347 6294
rect 10501 6354 10567 6357
rect 15334 6354 15394 6430
rect 15837 6427 15903 6430
rect 20069 6427 20135 6430
rect 20253 6490 20319 6493
rect 20253 6488 24180 6490
rect 20253 6432 20258 6488
rect 20314 6432 24180 6488
rect 20253 6430 24180 6432
rect 20253 6427 20319 6430
rect 10501 6352 15394 6354
rect 10501 6296 10506 6352
rect 10562 6296 15394 6352
rect 10501 6294 15394 6296
rect 20161 6354 20227 6357
rect 22461 6354 22527 6357
rect 23381 6354 23447 6357
rect 20161 6352 23447 6354
rect 20161 6296 20166 6352
rect 20222 6296 22466 6352
rect 22522 6296 23386 6352
rect 23442 6296 23447 6352
rect 20161 6294 23447 6296
rect 24120 6354 24180 6430
rect 25221 6354 25287 6357
rect 27520 6354 28000 6384
rect 24120 6352 25287 6354
rect 24120 6296 25226 6352
rect 25282 6296 25287 6352
rect 24120 6294 25287 6296
rect 10501 6291 10567 6294
rect 20161 6291 20227 6294
rect 22461 6291 22527 6294
rect 23381 6291 23447 6294
rect 25221 6291 25287 6294
rect 25454 6294 28000 6354
rect 4521 6218 4587 6221
rect 16481 6218 16547 6221
rect 4521 6216 16547 6218
rect 4521 6160 4526 6216
rect 4582 6160 16486 6216
rect 16542 6160 16547 6216
rect 4521 6158 16547 6160
rect 4521 6155 4587 6158
rect 16481 6155 16547 6158
rect 18965 6218 19031 6221
rect 19333 6218 19399 6221
rect 20897 6218 20963 6221
rect 18965 6216 20963 6218
rect 18965 6160 18970 6216
rect 19026 6160 19338 6216
rect 19394 6160 20902 6216
rect 20958 6160 20963 6216
rect 18965 6158 20963 6160
rect 18965 6155 19031 6158
rect 19333 6155 19399 6158
rect 20897 6155 20963 6158
rect 21541 6218 21607 6221
rect 24209 6218 24275 6221
rect 21541 6216 24275 6218
rect 21541 6160 21546 6216
rect 21602 6160 24214 6216
rect 24270 6160 24275 6216
rect 21541 6158 24275 6160
rect 21541 6155 21607 6158
rect 24209 6155 24275 6158
rect 9857 6082 9923 6085
rect 1580 6080 9923 6082
rect 1580 6024 9862 6080
rect 9918 6024 9923 6080
rect 1580 6022 9923 6024
rect 1580 5949 1640 6022
rect 9857 6019 9923 6022
rect 20069 6082 20135 6085
rect 24853 6082 24919 6085
rect 20069 6080 24919 6082
rect 20069 6024 20074 6080
rect 20130 6024 24858 6080
rect 24914 6024 24919 6080
rect 20069 6022 24919 6024
rect 20069 6019 20135 6022
rect 24853 6019 24919 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 1577 5944 1643 5949
rect 1577 5888 1582 5944
rect 1638 5888 1643 5944
rect 1577 5883 1643 5888
rect 3918 5884 3924 5948
rect 3988 5946 3994 5948
rect 4797 5946 4863 5949
rect 6269 5946 6335 5949
rect 3988 5944 6335 5946
rect 3988 5888 4802 5944
rect 4858 5888 6274 5944
rect 6330 5888 6335 5944
rect 3988 5886 6335 5888
rect 3988 5884 3994 5886
rect 4797 5883 4863 5886
rect 6269 5883 6335 5886
rect 10133 5810 10199 5813
rect 3558 5808 10199 5810
rect 3558 5752 10138 5808
rect 10194 5752 10199 5808
rect 3558 5750 10199 5752
rect 2773 5674 2839 5677
rect 3417 5674 3483 5677
rect 3558 5674 3618 5750
rect 10133 5747 10199 5750
rect 14733 5810 14799 5813
rect 20989 5810 21055 5813
rect 14733 5808 21055 5810
rect 14733 5752 14738 5808
rect 14794 5752 20994 5808
rect 21050 5752 21055 5808
rect 14733 5750 21055 5752
rect 14733 5747 14799 5750
rect 20989 5747 21055 5750
rect 2773 5672 3618 5674
rect 2773 5616 2778 5672
rect 2834 5616 3422 5672
rect 3478 5616 3618 5672
rect 2773 5614 3618 5616
rect 3693 5674 3759 5677
rect 4889 5674 4955 5677
rect 5901 5674 5967 5677
rect 3693 5672 5967 5674
rect 3693 5616 3698 5672
rect 3754 5616 4894 5672
rect 4950 5616 5906 5672
rect 5962 5616 5967 5672
rect 3693 5614 5967 5616
rect 2773 5611 2839 5614
rect 3417 5611 3483 5614
rect 3693 5611 3759 5614
rect 4889 5611 4955 5614
rect 5901 5611 5967 5614
rect 8661 5674 8727 5677
rect 12157 5674 12223 5677
rect 8661 5672 12223 5674
rect 8661 5616 8666 5672
rect 8722 5616 12162 5672
rect 12218 5616 12223 5672
rect 8661 5614 12223 5616
rect 8661 5611 8727 5614
rect 12157 5611 12223 5614
rect 17401 5674 17467 5677
rect 23197 5674 23263 5677
rect 25454 5674 25514 6294
rect 27520 6264 28000 6294
rect 17401 5672 25514 5674
rect 17401 5616 17406 5672
rect 17462 5616 23202 5672
rect 23258 5616 25514 5672
rect 17401 5614 25514 5616
rect 17401 5611 17467 5614
rect 23197 5611 23263 5614
rect 23841 5538 23907 5541
rect 15334 5536 23907 5538
rect 15334 5480 23846 5536
rect 23902 5480 23907 5536
rect 15334 5478 23907 5480
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 2957 5402 3023 5405
rect 2822 5400 3023 5402
rect 2822 5344 2962 5400
rect 3018 5344 3023 5400
rect 2822 5342 3023 5344
rect 2681 5130 2747 5133
rect 2822 5130 2882 5342
rect 2957 5339 3023 5342
rect 8385 5402 8451 5405
rect 12065 5402 12131 5405
rect 8385 5400 12131 5402
rect 8385 5344 8390 5400
rect 8446 5344 12070 5400
rect 12126 5344 12131 5400
rect 8385 5342 12131 5344
rect 8385 5339 8451 5342
rect 12065 5339 12131 5342
rect 3877 5266 3943 5269
rect 9029 5266 9095 5269
rect 3877 5264 9095 5266
rect 3877 5208 3882 5264
rect 3938 5208 9034 5264
rect 9090 5208 9095 5264
rect 3877 5206 9095 5208
rect 3877 5203 3943 5206
rect 9029 5203 9095 5206
rect 13077 5266 13143 5269
rect 15334 5266 15394 5478
rect 23841 5475 23907 5478
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 18045 5402 18111 5405
rect 21817 5402 21883 5405
rect 18045 5400 21883 5402
rect 18045 5344 18050 5400
rect 18106 5344 21822 5400
rect 21878 5344 21883 5400
rect 18045 5342 21883 5344
rect 18045 5339 18111 5342
rect 21817 5339 21883 5342
rect 20897 5266 20963 5269
rect 21909 5266 21975 5269
rect 24945 5266 25011 5269
rect 13077 5264 15394 5266
rect 13077 5208 13082 5264
rect 13138 5208 15394 5264
rect 13077 5206 15394 5208
rect 17358 5264 21466 5266
rect 17358 5208 20902 5264
rect 20958 5208 21466 5264
rect 17358 5206 21466 5208
rect 13077 5203 13143 5206
rect 3693 5130 3759 5133
rect 2681 5128 3759 5130
rect 2681 5072 2686 5128
rect 2742 5072 3698 5128
rect 3754 5072 3759 5128
rect 2681 5070 3759 5072
rect 2681 5067 2747 5070
rect 3693 5067 3759 5070
rect 3877 5130 3943 5133
rect 11513 5130 11579 5133
rect 17358 5130 17418 5206
rect 20897 5203 20963 5206
rect 3877 5128 17418 5130
rect 3877 5072 3882 5128
rect 3938 5072 11518 5128
rect 11574 5072 17418 5128
rect 3877 5070 17418 5072
rect 17585 5130 17651 5133
rect 21173 5130 21239 5133
rect 17585 5128 21239 5130
rect 17585 5072 17590 5128
rect 17646 5072 21178 5128
rect 21234 5072 21239 5128
rect 17585 5070 21239 5072
rect 21406 5130 21466 5206
rect 21909 5264 25011 5266
rect 21909 5208 21914 5264
rect 21970 5208 24950 5264
rect 25006 5208 25011 5264
rect 21909 5206 25011 5208
rect 21909 5203 21975 5206
rect 24945 5203 25011 5206
rect 22369 5130 22435 5133
rect 25037 5130 25103 5133
rect 21406 5128 25103 5130
rect 21406 5072 22374 5128
rect 22430 5072 25042 5128
rect 25098 5072 25103 5128
rect 21406 5070 25103 5072
rect 3877 5067 3943 5070
rect 11513 5067 11579 5070
rect 17585 5067 17651 5070
rect 21173 5067 21239 5070
rect 22369 5067 22435 5070
rect 25037 5067 25103 5070
rect 2773 4994 2839 4997
rect 6361 4994 6427 4997
rect 2773 4992 6427 4994
rect 2773 4936 2778 4992
rect 2834 4936 6366 4992
rect 6422 4936 6427 4992
rect 2773 4934 6427 4936
rect 2773 4931 2839 4934
rect 6361 4931 6427 4934
rect 13537 4994 13603 4997
rect 18321 4994 18387 4997
rect 13537 4992 18387 4994
rect 13537 4936 13542 4992
rect 13598 4936 18326 4992
rect 18382 4936 18387 4992
rect 13537 4934 18387 4936
rect 13537 4931 13603 4934
rect 18321 4931 18387 4934
rect 23565 4994 23631 4997
rect 25221 4994 25287 4997
rect 23565 4992 25287 4994
rect 23565 4936 23570 4992
rect 23626 4936 25226 4992
rect 25282 4936 25287 4992
rect 23565 4934 25287 4936
rect 23565 4931 23631 4934
rect 25221 4931 25287 4934
rect 10277 4928 10597 4929
rect 0 4858 480 4888
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 2405 4858 2471 4861
rect 0 4856 2471 4858
rect 0 4800 2410 4856
rect 2466 4800 2471 4856
rect 0 4798 2471 4800
rect 0 4768 480 4798
rect 2405 4795 2471 4798
rect 2865 4858 2931 4861
rect 9949 4858 10015 4861
rect 2865 4856 10015 4858
rect 2865 4800 2870 4856
rect 2926 4800 9954 4856
rect 10010 4800 10015 4856
rect 2865 4798 10015 4800
rect 2865 4795 2931 4798
rect 9949 4795 10015 4798
rect 23606 4796 23612 4860
rect 23676 4858 23682 4860
rect 27520 4858 28000 4888
rect 23676 4798 28000 4858
rect 23676 4796 23682 4798
rect 27520 4768 28000 4798
rect 4153 4722 4219 4725
rect 9397 4722 9463 4725
rect 4153 4720 9463 4722
rect 4153 4664 4158 4720
rect 4214 4664 9402 4720
rect 9458 4664 9463 4720
rect 4153 4662 9463 4664
rect 4153 4659 4219 4662
rect 9397 4659 9463 4662
rect 16665 4722 16731 4725
rect 24669 4722 24735 4725
rect 16665 4720 24735 4722
rect 16665 4664 16670 4720
rect 16726 4664 24674 4720
rect 24730 4664 24735 4720
rect 16665 4662 24735 4664
rect 16665 4659 16731 4662
rect 24669 4659 24735 4662
rect 3693 4586 3759 4589
rect 8937 4586 9003 4589
rect 3693 4584 8770 4586
rect 3693 4528 3698 4584
rect 3754 4528 8770 4584
rect 3693 4526 8770 4528
rect 3693 4523 3759 4526
rect 8710 4450 8770 4526
rect 8937 4584 19994 4586
rect 8937 4528 8942 4584
rect 8998 4528 19994 4584
rect 8937 4526 19994 4528
rect 8937 4523 9003 4526
rect 9765 4450 9831 4453
rect 19701 4450 19767 4453
rect 8710 4448 9831 4450
rect 8710 4392 9770 4448
rect 9826 4392 9831 4448
rect 8710 4390 9831 4392
rect 9765 4387 9831 4390
rect 16622 4448 19767 4450
rect 16622 4392 19706 4448
rect 19762 4392 19767 4448
rect 16622 4390 19767 4392
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 6361 4314 6427 4317
rect 9673 4314 9739 4317
rect 6361 4312 9739 4314
rect 6361 4256 6366 4312
rect 6422 4256 9678 4312
rect 9734 4256 9739 4312
rect 6361 4254 9739 4256
rect 6361 4251 6427 4254
rect 9673 4251 9739 4254
rect 2405 4178 2471 4181
rect 16622 4178 16682 4390
rect 19701 4387 19767 4390
rect 19934 4314 19994 4526
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 23565 4314 23631 4317
rect 19934 4312 23631 4314
rect 19934 4256 23570 4312
rect 23626 4256 23631 4312
rect 19934 4254 23631 4256
rect 23565 4251 23631 4254
rect 2405 4176 16682 4178
rect 2405 4120 2410 4176
rect 2466 4120 16682 4176
rect 2405 4118 16682 4120
rect 16849 4178 16915 4181
rect 19333 4178 19399 4181
rect 16849 4176 19399 4178
rect 16849 4120 16854 4176
rect 16910 4120 19338 4176
rect 19394 4120 19399 4176
rect 16849 4118 19399 4120
rect 2405 4115 2471 4118
rect 16849 4115 16915 4118
rect 19333 4115 19399 4118
rect 2681 4042 2747 4045
rect 8109 4042 8175 4045
rect 8569 4042 8635 4045
rect 2681 4040 8635 4042
rect 2681 3984 2686 4040
rect 2742 3984 8114 4040
rect 8170 3984 8574 4040
rect 8630 3984 8635 4040
rect 2681 3982 8635 3984
rect 2681 3979 2747 3982
rect 8109 3979 8175 3982
rect 8569 3979 8635 3982
rect 9581 4042 9647 4045
rect 11329 4042 11395 4045
rect 9581 4040 11395 4042
rect 9581 3984 9586 4040
rect 9642 3984 11334 4040
rect 11390 3984 11395 4040
rect 9581 3982 11395 3984
rect 9581 3979 9647 3982
rect 11329 3979 11395 3982
rect 15377 4042 15443 4045
rect 19425 4042 19491 4045
rect 15377 4040 19491 4042
rect 15377 3984 15382 4040
rect 15438 3984 19430 4040
rect 19486 3984 19491 4040
rect 15377 3982 19491 3984
rect 15377 3979 15443 3982
rect 19425 3979 19491 3982
rect 19977 4042 20043 4045
rect 22829 4042 22895 4045
rect 19977 4040 22895 4042
rect 19977 3984 19982 4040
rect 20038 3984 22834 4040
rect 22890 3984 22895 4040
rect 19977 3982 22895 3984
rect 19977 3979 20043 3982
rect 22829 3979 22895 3982
rect 25405 4042 25471 4045
rect 27429 4042 27495 4045
rect 25405 4040 27495 4042
rect 25405 3984 25410 4040
rect 25466 3984 27434 4040
rect 27490 3984 27495 4040
rect 25405 3982 27495 3984
rect 25405 3979 25471 3982
rect 27429 3979 27495 3982
rect 20529 3906 20595 3909
rect 23013 3906 23079 3909
rect 20529 3904 23079 3906
rect 20529 3848 20534 3904
rect 20590 3848 23018 3904
rect 23074 3848 23079 3904
rect 20529 3846 23079 3848
rect 20529 3843 20595 3846
rect 23013 3843 23079 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 1485 3770 1551 3773
rect 4429 3770 4495 3773
rect 21173 3770 21239 3773
rect 23749 3770 23815 3773
rect 1485 3768 8034 3770
rect 1485 3712 1490 3768
rect 1546 3712 4434 3768
rect 4490 3712 8034 3768
rect 1485 3710 8034 3712
rect 1485 3707 1551 3710
rect 4429 3707 4495 3710
rect 3785 3634 3851 3637
rect 7741 3634 7807 3637
rect 3785 3632 7807 3634
rect 3785 3576 3790 3632
rect 3846 3576 7746 3632
rect 7802 3576 7807 3632
rect 3785 3574 7807 3576
rect 7974 3634 8034 3710
rect 21173 3768 23815 3770
rect 21173 3712 21178 3768
rect 21234 3712 23754 3768
rect 23810 3712 23815 3768
rect 21173 3710 23815 3712
rect 21173 3707 21239 3710
rect 23749 3707 23815 3710
rect 12157 3634 12223 3637
rect 7974 3632 12223 3634
rect 7974 3576 12162 3632
rect 12218 3576 12223 3632
rect 7974 3574 12223 3576
rect 3785 3571 3851 3574
rect 7741 3571 7807 3574
rect 12157 3571 12223 3574
rect 12617 3634 12683 3637
rect 20161 3634 20227 3637
rect 12617 3632 20227 3634
rect 12617 3576 12622 3632
rect 12678 3576 20166 3632
rect 20222 3576 20227 3632
rect 12617 3574 20227 3576
rect 12617 3571 12683 3574
rect 20161 3571 20227 3574
rect 24669 3634 24735 3637
rect 24669 3632 25146 3634
rect 24669 3576 24674 3632
rect 24730 3576 25146 3632
rect 24669 3574 25146 3576
rect 24669 3571 24735 3574
rect 0 3498 480 3528
rect 1485 3498 1551 3501
rect 0 3496 1551 3498
rect 0 3440 1490 3496
rect 1546 3440 1551 3496
rect 0 3438 1551 3440
rect 0 3408 480 3438
rect 1485 3435 1551 3438
rect 20805 3498 20871 3501
rect 24853 3498 24919 3501
rect 20805 3496 24919 3498
rect 20805 3440 20810 3496
rect 20866 3440 24858 3496
rect 24914 3440 24919 3496
rect 20805 3438 24919 3440
rect 25086 3498 25146 3574
rect 27520 3498 28000 3528
rect 25086 3438 28000 3498
rect 20805 3435 20871 3438
rect 24853 3435 24919 3438
rect 27520 3408 28000 3438
rect 18321 3362 18387 3365
rect 21357 3362 21423 3365
rect 18321 3360 21423 3362
rect 18321 3304 18326 3360
rect 18382 3304 21362 3360
rect 21418 3304 21423 3360
rect 18321 3302 21423 3304
rect 18321 3299 18387 3302
rect 21357 3299 21423 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 1577 3226 1643 3229
rect 8109 3226 8175 3229
rect 12157 3226 12223 3229
rect 1577 3224 5458 3226
rect 1577 3168 1582 3224
rect 1638 3168 5458 3224
rect 1577 3166 5458 3168
rect 1577 3163 1643 3166
rect 1761 3090 1827 3093
rect 4981 3090 5047 3093
rect 1761 3088 5047 3090
rect 1761 3032 1766 3088
rect 1822 3032 4986 3088
rect 5042 3032 5047 3088
rect 1761 3030 5047 3032
rect 5398 3090 5458 3166
rect 8109 3224 12223 3226
rect 8109 3168 8114 3224
rect 8170 3168 12162 3224
rect 12218 3168 12223 3224
rect 8109 3166 12223 3168
rect 8109 3163 8175 3166
rect 12157 3163 12223 3166
rect 16389 3226 16455 3229
rect 22369 3226 22435 3229
rect 16389 3224 22435 3226
rect 16389 3168 16394 3224
rect 16450 3168 22374 3224
rect 22430 3168 22435 3224
rect 16389 3166 22435 3168
rect 16389 3163 16455 3166
rect 22369 3163 22435 3166
rect 10685 3090 10751 3093
rect 5398 3088 10751 3090
rect 5398 3032 10690 3088
rect 10746 3032 10751 3088
rect 5398 3030 10751 3032
rect 1761 3027 1827 3030
rect 4981 3027 5047 3030
rect 10685 3027 10751 3030
rect 14549 3090 14615 3093
rect 23473 3090 23539 3093
rect 14549 3088 23539 3090
rect 14549 3032 14554 3088
rect 14610 3032 23478 3088
rect 23534 3032 23539 3088
rect 14549 3030 23539 3032
rect 14549 3027 14615 3030
rect 23473 3027 23539 3030
rect 1485 2954 1551 2957
rect 5993 2954 6059 2957
rect 1485 2952 6059 2954
rect 1485 2896 1490 2952
rect 1546 2896 5998 2952
rect 6054 2896 6059 2952
rect 1485 2894 6059 2896
rect 1485 2891 1551 2894
rect 5993 2891 6059 2894
rect 10961 2954 11027 2957
rect 23381 2954 23447 2957
rect 10961 2952 23447 2954
rect 10961 2896 10966 2952
rect 11022 2896 23386 2952
rect 23442 2896 23447 2952
rect 10961 2894 23447 2896
rect 10961 2891 11027 2894
rect 23381 2891 23447 2894
rect 2497 2818 2563 2821
rect 8661 2818 8727 2821
rect 2497 2816 8727 2818
rect 2497 2760 2502 2816
rect 2558 2760 8666 2816
rect 8722 2760 8727 2816
rect 2497 2758 8727 2760
rect 2497 2755 2563 2758
rect 8661 2755 8727 2758
rect 11237 2818 11303 2821
rect 15469 2818 15535 2821
rect 11237 2816 15535 2818
rect 11237 2760 11242 2816
rect 11298 2760 15474 2816
rect 15530 2760 15535 2816
rect 11237 2758 15535 2760
rect 11237 2755 11303 2758
rect 15469 2755 15535 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 5165 2682 5231 2685
rect 7465 2682 7531 2685
rect 5165 2680 7531 2682
rect 5165 2624 5170 2680
rect 5226 2624 7470 2680
rect 7526 2624 7531 2680
rect 5165 2622 7531 2624
rect 5165 2619 5231 2622
rect 7465 2619 7531 2622
rect 12525 2682 12591 2685
rect 15653 2682 15719 2685
rect 12525 2680 15719 2682
rect 12525 2624 12530 2680
rect 12586 2624 15658 2680
rect 15714 2624 15719 2680
rect 12525 2622 15719 2624
rect 12525 2619 12591 2622
rect 15653 2619 15719 2622
rect 20621 2682 20687 2685
rect 25221 2682 25287 2685
rect 20621 2680 25287 2682
rect 20621 2624 20626 2680
rect 20682 2624 25226 2680
rect 25282 2624 25287 2680
rect 20621 2622 25287 2624
rect 20621 2619 20687 2622
rect 25221 2619 25287 2622
rect 4981 2546 5047 2549
rect 8293 2546 8359 2549
rect 4981 2544 8359 2546
rect 4981 2488 4986 2544
rect 5042 2488 8298 2544
rect 8354 2488 8359 2544
rect 4981 2486 8359 2488
rect 4981 2483 5047 2486
rect 8293 2483 8359 2486
rect 8569 2546 8635 2549
rect 11145 2546 11211 2549
rect 8569 2544 11211 2546
rect 8569 2488 8574 2544
rect 8630 2488 11150 2544
rect 11206 2488 11211 2544
rect 8569 2486 11211 2488
rect 8569 2483 8635 2486
rect 11145 2483 11211 2486
rect 18137 2546 18203 2549
rect 24117 2546 24183 2549
rect 18137 2544 24183 2546
rect 18137 2488 18142 2544
rect 18198 2488 24122 2544
rect 24178 2488 24183 2544
rect 18137 2486 24183 2488
rect 18137 2483 18203 2486
rect 24117 2483 24183 2486
rect 473 2410 539 2413
rect 1485 2410 1551 2413
rect 473 2408 1551 2410
rect 473 2352 478 2408
rect 534 2352 1490 2408
rect 1546 2352 1551 2408
rect 473 2350 1551 2352
rect 473 2347 539 2350
rect 1485 2347 1551 2350
rect 4521 2410 4587 2413
rect 9489 2410 9555 2413
rect 11421 2410 11487 2413
rect 4521 2408 11487 2410
rect 4521 2352 4526 2408
rect 4582 2352 9494 2408
rect 9550 2352 11426 2408
rect 11482 2352 11487 2408
rect 4521 2350 11487 2352
rect 4521 2347 4587 2350
rect 9489 2347 9555 2350
rect 11421 2347 11487 2350
rect 18321 2410 18387 2413
rect 24301 2410 24367 2413
rect 18321 2408 24367 2410
rect 18321 2352 18326 2408
rect 18382 2352 24306 2408
rect 24362 2352 24367 2408
rect 18321 2350 24367 2352
rect 18321 2347 18387 2350
rect 24301 2347 24367 2350
rect 16481 2274 16547 2277
rect 16481 2272 21834 2274
rect 16481 2216 16486 2272
rect 16542 2216 21834 2272
rect 16481 2214 21834 2216
rect 16481 2211 16547 2214
rect 5610 2208 5930 2209
rect 0 2138 480 2168
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 1301 2138 1367 2141
rect 0 2136 1367 2138
rect 0 2080 1306 2136
rect 1362 2080 1367 2136
rect 0 2078 1367 2080
rect 0 2048 480 2078
rect 1301 2075 1367 2078
rect 17125 2138 17191 2141
rect 21541 2138 21607 2141
rect 17125 2136 21607 2138
rect 17125 2080 17130 2136
rect 17186 2080 21546 2136
rect 21602 2080 21607 2136
rect 17125 2078 21607 2080
rect 17125 2075 17191 2078
rect 21541 2075 21607 2078
rect 5441 2002 5507 2005
rect 9765 2002 9831 2005
rect 5441 2000 9831 2002
rect 5441 1944 5446 2000
rect 5502 1944 9770 2000
rect 9826 1944 9831 2000
rect 5441 1942 9831 1944
rect 5441 1939 5507 1942
rect 9765 1939 9831 1942
rect 9949 2002 10015 2005
rect 19701 2002 19767 2005
rect 9949 2000 19767 2002
rect 9949 1944 9954 2000
rect 10010 1944 19706 2000
rect 19762 1944 19767 2000
rect 9949 1942 19767 1944
rect 21774 2002 21834 2214
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 26141 2138 26207 2141
rect 27520 2138 28000 2168
rect 26141 2136 28000 2138
rect 26141 2080 26146 2136
rect 26202 2080 28000 2136
rect 26141 2078 28000 2080
rect 26141 2075 26207 2078
rect 27520 2048 28000 2078
rect 25221 2002 25287 2005
rect 21774 2000 25287 2002
rect 21774 1944 25226 2000
rect 25282 1944 25287 2000
rect 21774 1942 25287 1944
rect 9949 1939 10015 1942
rect 19701 1939 19767 1942
rect 25221 1939 25287 1942
rect 2129 1866 2195 1869
rect 13261 1866 13327 1869
rect 2129 1864 13327 1866
rect 2129 1808 2134 1864
rect 2190 1808 13266 1864
rect 13322 1808 13327 1864
rect 2129 1806 13327 1808
rect 2129 1803 2195 1806
rect 13261 1803 13327 1806
rect 15377 1866 15443 1869
rect 25129 1866 25195 1869
rect 15377 1864 25195 1866
rect 15377 1808 15382 1864
rect 15438 1808 25134 1864
rect 25190 1808 25195 1864
rect 15377 1806 25195 1808
rect 15377 1803 15443 1806
rect 25129 1803 25195 1806
rect 5993 1730 6059 1733
rect 17125 1730 17191 1733
rect 5993 1728 17191 1730
rect 5993 1672 5998 1728
rect 6054 1672 17130 1728
rect 17186 1672 17191 1728
rect 5993 1670 17191 1672
rect 5993 1667 6059 1670
rect 17125 1667 17191 1670
rect 17309 1730 17375 1733
rect 20713 1730 20779 1733
rect 17309 1728 20779 1730
rect 17309 1672 17314 1728
rect 17370 1672 20718 1728
rect 20774 1672 20779 1728
rect 17309 1670 20779 1672
rect 17309 1667 17375 1670
rect 20713 1667 20779 1670
rect 3877 1594 3943 1597
rect 12709 1594 12775 1597
rect 3877 1592 12775 1594
rect 3877 1536 3882 1592
rect 3938 1536 12714 1592
rect 12770 1536 12775 1592
rect 3877 1534 12775 1536
rect 3877 1531 3943 1534
rect 12709 1531 12775 1534
rect 12893 1594 12959 1597
rect 24025 1594 24091 1597
rect 12893 1592 24091 1594
rect 12893 1536 12898 1592
rect 12954 1536 24030 1592
rect 24086 1536 24091 1592
rect 12893 1534 24091 1536
rect 12893 1531 12959 1534
rect 24025 1531 24091 1534
rect 3233 1458 3299 1461
rect 8845 1458 8911 1461
rect 3233 1456 8911 1458
rect 3233 1400 3238 1456
rect 3294 1400 8850 1456
rect 8906 1400 8911 1456
rect 3233 1398 8911 1400
rect 3233 1395 3299 1398
rect 8845 1395 8911 1398
rect 10777 1458 10843 1461
rect 23749 1458 23815 1461
rect 10777 1456 23815 1458
rect 10777 1400 10782 1456
rect 10838 1400 23754 1456
rect 23810 1400 23815 1456
rect 10777 1398 23815 1400
rect 10777 1395 10843 1398
rect 23749 1395 23815 1398
rect 0 778 480 808
rect 2773 778 2839 781
rect 0 776 2839 778
rect 0 720 2778 776
rect 2834 720 2839 776
rect 0 718 2839 720
rect 0 688 480 718
rect 2773 715 2839 718
rect 22921 778 22987 781
rect 27520 778 28000 808
rect 22921 776 28000 778
rect 22921 720 22926 776
rect 22982 720 28000 776
rect 22921 718 28000 720
rect 22921 715 22987 718
rect 27520 688 28000 718
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 3004 23564 3068 23628
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 3924 19408 3988 19412
rect 3924 19352 3938 19408
rect 3938 19352 3988 19408
rect 3924 19348 3988 19352
rect 19196 19136 19260 19140
rect 19196 19080 19246 19136
rect 19246 19080 19260 19136
rect 19196 19076 19260 19080
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 1532 16280 1596 16284
rect 1532 16224 1582 16280
rect 1582 16224 1596 16280
rect 1532 16220 1596 16224
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 21404 14860 21468 14924
rect 9812 14724 9876 14788
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 3740 14452 3804 14516
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 23612 13636 23676 13700
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 19196 13092 19260 13156
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 23612 12956 23676 13020
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 9812 12140 9876 12204
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 21404 11868 21468 11932
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 3188 9964 3252 10028
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 1532 7788 1596 7852
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 3188 7304 3252 7308
rect 3188 7248 3202 7304
rect 3202 7248 3252 7304
rect 3188 7244 3252 7248
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 3004 6896 3068 6900
rect 3004 6840 3018 6896
rect 3018 6840 3068 6896
rect 3004 6836 3068 6840
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 3740 6428 3804 6492
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 3924 5884 3988 5948
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 23612 4796 23676 4860
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 3003 23628 3069 23629
rect 3003 23564 3004 23628
rect 3068 23564 3069 23628
rect 3003 23563 3069 23564
rect 1531 16284 1597 16285
rect 1531 16220 1532 16284
rect 1596 16220 1597 16284
rect 1531 16219 1597 16220
rect 1534 7853 1594 16219
rect 1531 7852 1597 7853
rect 1531 7788 1532 7852
rect 1596 7788 1597 7852
rect 1531 7787 1597 7788
rect 3006 6901 3066 23563
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 3923 19412 3989 19413
rect 3923 19348 3924 19412
rect 3988 19348 3989 19412
rect 3923 19347 3989 19348
rect 3739 14516 3805 14517
rect 3739 14452 3740 14516
rect 3804 14452 3805 14516
rect 3739 14451 3805 14452
rect 3187 10028 3253 10029
rect 3187 9964 3188 10028
rect 3252 9964 3253 10028
rect 3187 9963 3253 9964
rect 3190 7309 3250 9963
rect 3187 7308 3253 7309
rect 3187 7244 3188 7308
rect 3252 7244 3253 7308
rect 3187 7243 3253 7244
rect 3003 6900 3069 6901
rect 3003 6836 3004 6900
rect 3068 6836 3069 6900
rect 3003 6835 3069 6836
rect 3742 6493 3802 14451
rect 3739 6492 3805 6493
rect 3739 6428 3740 6492
rect 3804 6428 3805 6492
rect 3739 6427 3805 6428
rect 3926 5949 3986 19347
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 9811 14788 9877 14789
rect 9811 14724 9812 14788
rect 9876 14724 9877 14788
rect 9811 14723 9877 14724
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 9814 12205 9874 14723
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 9811 12204 9877 12205
rect 9811 12140 9812 12204
rect 9876 12140 9877 12204
rect 9811 12139 9877 12140
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 3923 5948 3989 5949
rect 3923 5884 3924 5948
rect 3988 5884 3989 5948
rect 3923 5883 3989 5884
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19195 19140 19261 19141
rect 19195 19076 19196 19140
rect 19260 19076 19261 19140
rect 19195 19075 19261 19076
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 19198 13157 19258 19075
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 21403 14924 21469 14925
rect 21403 14860 21404 14924
rect 21468 14860 21469 14924
rect 21403 14859 21469 14860
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19195 13156 19261 13157
rect 19195 13092 19196 13156
rect 19260 13092 19261 13156
rect 19195 13091 19261 13092
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 21406 11933 21466 14859
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 23611 13700 23677 13701
rect 23611 13636 23612 13700
rect 23676 13636 23677 13700
rect 23611 13635 23677 13636
rect 23614 13021 23674 13635
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 23611 13020 23677 13021
rect 23611 12956 23612 13020
rect 23676 12956 23677 13020
rect 23611 12955 23677 12956
rect 21403 11932 21469 11933
rect 21403 11868 21404 11932
rect 21468 11868 21469 11932
rect 21403 11867 21469 11868
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 23614 4861 23674 12955
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 23611 4860 23677 4861
rect 23611 4796 23612 4860
rect 23676 4796 23677 4860
rect 23611 4795 23677 4796
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _090_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _172_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _183_
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__C
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_16
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_20
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__B
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_35
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_33
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_38
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_39
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_50 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_54 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6072 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6900 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_76
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _119_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _173_
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_80
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_78
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_91
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__B
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__B
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _278_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__C
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_or4_4  _186_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _184_
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_108
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_116
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_141
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_148
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_152
timestamp 1586364061
transform 1 0 15088 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_159
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _175_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_161
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_163
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__277__A
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_188
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_198 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_200
timestamp 1586364061
transform 1 0 19504 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_205
timestamp 1586364061
transform 1 0 19964 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_228
timestamp 1586364061
transform 1 0 22080 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_225
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_232
timestamp 1586364061
transform 1 0 22448 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _276_
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__276__A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_or4_4  _139_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_254
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_258
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_266
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_2  _274_
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__274__A
timestamp 1586364061
transform 1 0 26128 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_270
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_274
timestamp 1586364061
transform 1 0 26312 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _118_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_47
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_51
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_1  _089_
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_58
timestamp 1586364061
transform 1 0 6440 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_62
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_65
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_75
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_79
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_101
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use scs8hd_or4_4  _174_
timestamp 1586364061
transform 1 0 10580 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__D
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_112
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 222 592
use scs8hd_or2_4  _185_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__186__D
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_116
timestamp 1586364061
transform 1 0 11776 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__185__B
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_2  _277_
timestamp 1586364061
transform 1 0 17112 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_172
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_1  _141_
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_195
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_219
timestamp 1586364061
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _182_
timestamp 1586364061
transform 1 0 23184 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 23000 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22632 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_232
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_236
timestamp 1586364061
transform 1 0 22816 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_249
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_253
timestamp 1586364061
transform 1 0 24380 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _146_
timestamp 1586364061
transform 1 0 24748 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_266
timestamp 1586364061
transform 1 0 25576 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_nand2_4  _151_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _171_
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__D
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_17
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_21
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_55
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_or2_4  _092_
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__197__B
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _091_
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__197__C
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _140_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__B
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_126
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13892 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_130
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_148
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_152
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_164
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_212
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_216
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_223
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_235
timestamp 1586364061
transform 1 0 22724 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_254
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _273_
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__273__A
timestamp 1586364061
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_266
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_3_270 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25944 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_276
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_or4_4  _120_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__C
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_40
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_75
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__D
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_79
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_or4_4  _197_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _193_
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__224__C
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__B
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__278__A
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_123
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_147
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_160
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_171
timestamp 1586364061
transform 1 0 16836 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_175
timestamp 1586364061
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_179
timestamp 1586364061
transform 1 0 17572 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_183
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_195
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 21068 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_228
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22816 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22540 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_232
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_235
timestamp 1586364061
transform 1 0 22724 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 24380 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_245
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_249
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_252
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_262 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25208 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_or4_4  _093_
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__B
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_32
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_37
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_49
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_73
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_77
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_or4_4  _216_
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__A
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__224__B
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_90
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__C
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_115
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use scs8hd_buf_1  _176_
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_131
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_150
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_169
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_199
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_203
timestamp 1586364061
transform 1 0 19780 0 1 4896
box -38 -48 314 592
use scs8hd_buf_2  _275_
timestamp 1586364061
transform 1 0 20056 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__275__A
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_210
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_214
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_229
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_233
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_237
timestamp 1586364061
transform 1 0 22908 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_241
timestamp 1586364061
transform 1 0 23276 0 1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _272_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__272__A
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_266
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_5_270
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use scs8hd_inv_8  _138_
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__C
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_10
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_nor2_4  _190_
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 866 592
use scs8hd_or4_4  _208_
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__232__C
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__D
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__B
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_19
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4324 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_32
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_46
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_50
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_49
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_54
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_58
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_75
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__B
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_79
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_78
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_82
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_1  _088_
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_97
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__224__D
timestamp 1586364061
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use scs8hd_or4_4  _224_
timestamp 1586364061
transform 1 0 10304 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _195_
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__D
timestamp 1586364061
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_109
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_113
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_111
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_115
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _179_
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12696 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_128
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13708 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13156 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_129
timestamp 1586364061
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_133
timestamp 1586364061
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_146
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_150
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_165
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_163
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_167
timestamp 1586364061
transform 1 0 16468 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_7_.latch
timestamp 1586364061
transform 1 0 18124 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_182
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _177_
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_200
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_203
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _181_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_213
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_218
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_228
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22540 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_242
timestamp 1586364061
transform 1 0 23368 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_233
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_237
timestamp 1586364061
transform 1 0 22908 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 24104 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _155_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_247
timestamp 1586364061
transform 1 0 23828 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_254
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 406 592
use scs8hd_buf_2  _271_
timestamp 1586364061
transform 1 0 25208 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__271__A
timestamp 1586364061
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 25116 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_259
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_260
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_266
timestamp 1586364061
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_7_270
timestamp 1586364061
transform 1 0 25944 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_276
timestamp 1586364061
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__D
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _232_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 4140 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__232__D
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_42
timestamp 1586364061
transform 1 0 4968 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_61
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__B
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_78
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_82
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_86
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _196_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__B
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_113
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_6  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_123
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _178_
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_157
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_161
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_174
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_6_.latch
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_197
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 20148 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_209
timestamp 1586364061
transform 1 0 20332 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 21528 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21344 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_219
timestamp 1586364061
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23276 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22724 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_233
timestamp 1586364061
transform 1 0 22540 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_237
timestamp 1586364061
transform 1 0 22908 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_250
timestamp 1586364061
transform 1 0 24104 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_254
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 24840 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_267
timestamp 1586364061
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_8
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_13
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__190__B
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_29
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_33
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_37
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_82
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _225_
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_104
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_108
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_116
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_120
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_126
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_145
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_162
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_166
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_9_189
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_216
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 21528 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_233
timestamp 1586364061
transform 1 0 22540 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_237
timestamp 1586364061
transform 1 0 22908 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_265
timestamp 1586364061
transform 1 0 25484 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_273
timestamp 1586364061
transform 1 0 26220 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_20
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_24
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_28
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_49
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _194_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_72
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_10_104
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_123
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_131
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_3  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_160
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_164
timestamp 1586364061
transform 1 0 16192 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_10_179
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_200
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_212
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_7_.latch
timestamp 1586364061
transform 1 0 21804 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 21620 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_221
timestamp 1586364061
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_236
timestamp 1586364061
transform 1 0 22816 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23552 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_253
timestamp 1586364061
transform 1 0 24380 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25116 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_264
timestamp 1586364061
transform 1 0 25392 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_272
timestamp 1586364061
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_8  _150_
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_14
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_18
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_37
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__191__B
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_81
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_85
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_102
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_106
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_144
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_148
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_152
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_167
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_188
timestamp 1586364061
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_192
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_205
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_209
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_216
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_6_.latch
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_236
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_254
timestamp 1586364061
transform 1 0 24472 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_258
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_261
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_265
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_buf_1  _086_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _084_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__189__B
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _082_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__C
timestamp 1586364061
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_49
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _191_
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_62
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__192__B
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_66
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_81
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_85
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_89
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_12_118
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_130
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_134
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_138
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_164
timestamp 1586364061
transform 1 0 16192 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16928 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_12_168
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_12_181
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_189
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_201
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 21620 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_219
timestamp 1586364061
transform 1 0 21252 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 23368 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23184 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_234
timestamp 1586364061
transform 1 0 22632 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_238
timestamp 1586364061
transform 1 0 23000 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_255
timestamp 1586364061
transform 1 0 24564 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_262
timestamp 1586364061
transform 1 0 25208 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_1  _134_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_or4_4  _152_
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__C
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_or3_4  _085_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _189_
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_14
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_or3_4  _112_
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 866 592
use scs8hd_or3_4  _115_
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_13_49
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_14_49
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 590 592
use scs8hd_or3_4  _103_
timestamp 1586364061
transform 1 0 6348 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _192_
timestamp 1586364061
transform 1 0 6900 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__C
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_55
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _206_
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_72
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_66
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_14_74
timestamp 1586364061
transform 1 0 7912 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__206__B
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_90
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_107
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_111
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_112
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_120
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_121
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_142
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_154
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _121_
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_6  FILLER_13_142
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 590 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_158
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_167
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_171
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_189
timestamp 1586364061
transform 1 0 18492 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_185
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_187
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__B
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_191
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_195
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_205
timestamp 1586364061
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_209
timestamp 1586364061
transform 1 0 20332 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_212
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_216
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20700 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_218
timestamp 1586364061
transform 1 0 21160 0 -1 10336
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_224
timestamp 1586364061
transform 1 0 21712 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23276 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_237
timestamp 1586364061
transform 1 0 22908 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_243
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_254
timestamp 1586364061
transform 1 0 24472 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _270_
timestamp 1586364061
transform 1 0 25208 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_265
timestamp 1586364061
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_266
timestamp 1586364061
transform 1 0 25576 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__270__A
timestamp 1586364061
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_273
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_or3_4  _100_
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__097__C
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_21
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_25
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _083_
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _126_
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__109__C
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__B
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_42
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_46
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_68
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_81
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_85
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_100
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _116_
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_104
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_140
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_15_154
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _227_
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__227__B
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_158
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_178
timestamp 1586364061
transform 1 0 17480 0 1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _228_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_203
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_207
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_219
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_223
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_260
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_265
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_273
timestamp 1586364061
transform 1 0 26220 0 1 10336
box -38 -48 406 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__D
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__B
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_or3_4  _097_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_or3_4  _109_
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__200__B
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_45
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _207_
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_6  FILLER_16_62
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_81
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_6  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 590 592
use scs8hd_buf_1  _104_
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_124
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_128
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_132
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_165
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17296 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_16_173
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_187
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_195
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_212
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_229
timestamp 1586364061
transform 1 0 22172 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_233
timestamp 1586364061
transform 1 0 22540 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_236
timestamp 1586364061
transform 1 0 22816 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_240
timestamp 1586364061
transform 1 0 23184 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_250
timestamp 1586364061
transform 1 0 24104 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_254
timestamp 1586364061
transform 1 0 24472 0 -1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 24840 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_267
timestamp 1586364061
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 406 592
use scs8hd_buf_1  _124_
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 314 592
use scs8hd_buf_1  _130_
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _106_
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_31
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_44
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _113_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__203__B
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_55
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__B
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_65
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_69
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _107_
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_103
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_107
timestamp 1586364061
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _226_
timestamp 1586364061
transform 1 0 12512 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__B
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_133
timestamp 1586364061
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_137
timestamp 1586364061
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_169
timestamp 1586364061
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_173
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_177
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_189
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_6_.latch
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_17_204
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_209
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_224
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_228
timestamp 1586364061
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_235
timestamp 1586364061
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_239
timestamp 1586364061
transform 1 0 23092 0 1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _265_
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__265__A
timestamp 1586364061
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_266
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_17_270
timestamp 1586364061
transform 1 0 25944 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_276
timestamp 1586364061
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__100__C
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _230_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_6  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 590 592
use scs8hd_nor2_4  _200_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _203_
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_45
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_58
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _204_
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_101
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_111
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_135
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_139
timestamp 1586364061
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_143
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_151
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_186
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_18_194
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_226
timestamp 1586364061
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_230
timestamp 1586364061
transform 1 0 22264 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_18_243
timestamp 1586364061
transform 1 0 23460 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 23644 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_247
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_260
timestamp 1586364061
transform 1 0 25024 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_272
timestamp 1586364061
transform 1 0 26128 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__260__A
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_10
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _110_
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 866 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_14
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_21
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_25
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_21
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_25
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_7_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__201__B
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_38
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_46
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_43
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_20_51
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_58
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_73
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_67
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_1  _101_
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_84
timestamp 1586364061
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__B
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_103
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_104
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_115
timestamp 1586364061
transform 1 0 11684 0 -1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_127
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_131
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_136
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_140
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_148
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_152
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_168
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_184
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_197
timestamp 1586364061
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_201
timestamp 1586364061
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_205
timestamp 1586364061
transform 1 0 19964 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_210
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_206
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20792 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_225
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_229
timestamp 1586364061
transform 1 0 22172 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_219
timestamp 1586364061
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_229
timestamp 1586364061
transform 1 0 22172 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22908 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24472 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_252
timestamp 1586364061
transform 1 0 24288 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_256
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_246
timestamp 1586364061
transform 1 0 23736 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_267
timestamp 1586364061
transform 1 0 25668 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_257
timestamp 1586364061
transform 1 0 24748 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_269
timestamp 1586364061
transform 1 0 25852 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_1  _199_
timestamp 1586364061
transform 1 0 1840 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_6_.latch
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_34
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_47
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__B
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_55
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_78
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_85
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_89
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__214__A
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__214__B
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_105
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_109
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_112
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_116
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_134
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_148
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_161
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_165
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_169
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_212
timestamp 1586364061
transform 1 0 20608 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_217
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  FILLER_21_229
timestamp 1586364061
transform 1 0 22172 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_234
timestamp 1586364061
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_238
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__269__A
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_254
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_265
timestamp 1586364061
transform 1 0 25484 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_buf_2  _260_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _201_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_29
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _202_
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_60
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_79
timestamp 1586364061
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_87
timestamp 1586364061
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _205_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _214_
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__213__B
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_107
timestamp 1586364061
transform 1 0 10948 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_119
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_136
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_150
timestamp 1586364061
transform 1 0 14904 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_171
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_176
timestamp 1586364061
transform 1 0 17296 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_187
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_210
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_228
timestamp 1586364061
transform 1 0 22080 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_22_241
timestamp 1586364061
transform 1 0 23276 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_2  _269_
timestamp 1586364061
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_247
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_259
timestamp 1586364061
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_271
timestamp 1586364061
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_1  _188_
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_8
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_12
timestamp 1586364061
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__256__A
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_19
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__B
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_90
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_94
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_97
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _213_
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__213__A
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_114
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__215__A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__215__B
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_126
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_130
timestamp 1586364061
transform 1 0 13064 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_134
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_146
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_163
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_201
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_7_.latch
timestamp 1586364061
transform 1 0 20516 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22264 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_222
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_226
timestamp 1586364061
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23092 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_233
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_237
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_241
timestamp 1586364061
transform 1 0 23276 0 1 14688
box -38 -48 314 592
use scs8hd_conb_1  _248_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_248
timestamp 1586364061
transform 1 0 23920 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_252
timestamp 1586364061
transform 1 0 24288 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_259
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_263
timestamp 1586364061
transform 1 0 25300 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_275
timestamp 1586364061
transform 1 0 26404 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _256_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_7
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_11
timestamp 1586364061
transform 1 0 2116 0 -1 15776
box -38 -48 406 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_18
timestamp 1586364061
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_29
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_24_40
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_51
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_74
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_78
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 590 592
use scs8hd_nor2_4  _229_
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _215_
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_104
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_121
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_24_140
timestamp 1586364061
transform 1 0 13984 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_148
timestamp 1586364061
transform 1 0 14720 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_151
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_6  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18124 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_183
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_187
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_200
timestamp 1586364061
transform 1 0 19504 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_204
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_212
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22080 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_226
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_230
timestamp 1586364061
transform 1 0 22264 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22632 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_237
timestamp 1586364061
transform 1 0 22908 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_248
timestamp 1586364061
transform 1 0 23920 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _259_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__259__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_25
timestamp 1586364061
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_44
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_48
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_67
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_84
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_87
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_91
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_106
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_112
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_116
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13064 0 1 15776
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_25_141
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_210
timestamp 1586364061
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_221
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_225
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_239
timestamp 1586364061
transform 1 0 23092 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_243
timestamp 1586364061
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use scs8hd_buf_2  _268_
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_253
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__268__A
timestamp 1586364061
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_259
timestamp 1586364061
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_263
timestamp 1586364061
transform 1 0 25300 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_267
timestamp 1586364061
transform 1 0 25668 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_275
timestamp 1586364061
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _187_
timestamp 1586364061
transform 1 0 1932 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _258_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__258__A
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_8  FILLER_26_12
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _209_
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 2300 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_23
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_34
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_43
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_47
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_60
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_55
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__221__B
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_106
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_109
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_113
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _210_
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__221__A
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__210__B
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_116
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_120
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__219__A
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_140
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__219__B
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_142
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_146
timestamp 1586364061
transform 1 0 14536 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16100 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_155
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_170
timestamp 1586364061
transform 1 0 16744 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_176
timestamp 1586364061
transform 1 0 17296 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_174
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_178
timestamp 1586364061
transform 1 0 17480 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__212__B
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_188
timestamp 1586364061
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_192
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__212__A
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_205
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_197
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_204
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20608 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_213
timestamp 1586364061
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_218
timestamp 1586364061
transform 1 0 21160 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_215
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22080 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_229
timestamp 1586364061
transform 1 0 22172 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_219
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_226
timestamp 1586364061
transform 1 0 21896 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_230
timestamp 1586364061
transform 1 0 22264 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22908 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_240
timestamp 1586364061
transform 1 0 23184 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_6  FILLER_27_234
timestamp 1586364061
transform 1 0 22632 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_242
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _246_
timestamp 1586364061
transform 1 0 23920 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _267_
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_253
timestamp 1586364061
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24932 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__267__A
timestamp 1586364061
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_262
timestamp 1586364061
transform 1 0 25208 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_259
timestamp 1586364061
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_263
timestamp 1586364061
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_274
timestamp 1586364061
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_275
timestamp 1586364061
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _198_
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_8  FILLER_28_12
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 774 592
use scs8hd_conb_1  _243_
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__238__B
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_29
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__B
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_45
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_49
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5980 0 -1 17952
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__231__B
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_81
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_87
timestamp 1586364061
transform 1 0 9108 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_100
timestamp 1586364061
transform 1 0 10304 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_110
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 774 592
use scs8hd_nor2_4  _221_
timestamp 1586364061
transform 1 0 11960 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_28_127
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _219_
timestamp 1586364061
transform 1 0 13524 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_131
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_144
timestamp 1586364061
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_148
timestamp 1586364061
transform 1 0 14720 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_152
timestamp 1586364061
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16008 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_160
timestamp 1586364061
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_164
timestamp 1586364061
transform 1 0 16192 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_28_179
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _212_
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_183
timestamp 1586364061
transform 1 0 17940 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_196
timestamp 1586364061
transform 1 0 19136 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_208
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_8  FILLER_28_218
timestamp 1586364061
transform 1 0 21160 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_226
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23184 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_232
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_243
timestamp 1586364061
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_255
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_267
timestamp 1586364061
transform 1 0 25668 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_8
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_12
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _249_
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_19
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _238_
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 866 592
use scs8hd_decap_6  FILLER_29_36
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 590 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 866 592
use scs8hd_fill_1  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_76
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 406 592
use scs8hd_nor2_4  _231_
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_83
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__222__B
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _222_
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _223_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _218_
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__218__A
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_149
timestamp 1586364061
transform 1 0 14812 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_153
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_156
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__211__B
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_204
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _250_
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_215
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 774 592
use scs8hd_conb_1  _251_
timestamp 1586364061
transform 1 0 21620 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_226
timestamp 1586364061
transform 1 0 21896 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_29_238
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__279__A
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_253
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_12
timestamp 1586364061
transform 1 0 2208 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 406 592
use scs8hd_conb_1  _245_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__237__B
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_29
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_35
timestamp 1586364061
transform 1 0 4324 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _235_
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__B
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_39
timestamp 1586364061
transform 1 0 4692 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_42
timestamp 1586364061
transform 1 0 4968 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_55
timestamp 1586364061
transform 1 0 6164 0 -1 19040
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_72
timestamp 1586364061
transform 1 0 7728 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_76
timestamp 1586364061
transform 1 0 8096 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9844 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_97
timestamp 1586364061
transform 1 0 10028 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_111
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__223__B
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_118
timestamp 1586364061
transform 1 0 11960 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_122
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__218__B
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_138
timestamp 1586364061
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_142
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_165
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _211_
timestamp 1586364061
transform 1 0 17020 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_169
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_182
timestamp 1586364061
transform 1 0 17848 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_186
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_193
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_8  FILLER_30_204
timestamp 1586364061
transform 1 0 19872 0 -1 19040
box -38 -48 774 592
use scs8hd_conb_1  _242_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_212
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_218
timestamp 1586364061
transform 1 0 21160 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_230
timestamp 1586364061
transform 1 0 22264 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_242
timestamp 1586364061
transform 1 0 23368 0 -1 19040
box -38 -48 1142 592
use scs8hd_buf_2  _279_
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_254
timestamp 1586364061
transform 1 0 24472 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_259
timestamp 1586364061
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_271
timestamp 1586364061
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_2  _257_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__257__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_23
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _237_
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _234_
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7728 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_66
timestamp 1586364061
transform 1 0 7176 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_83
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_87
timestamp 1586364061
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_31_102
timestamp 1586364061
transform 1 0 10488 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _217_
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__217__A
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_106
timestamp 1586364061
transform 1 0 10856 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12512 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_139
timestamp 1586364061
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_161
timestamp 1586364061
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_165
timestamp 1586364061
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_172
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_176
timestamp 1586364061
transform 1 0 17296 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_181
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_187
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_191
timestamp 1586364061
transform 1 0 18676 0 1 19040
box -38 -48 406 592
use scs8hd_buf_1  _154_
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 19872 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_198
timestamp 1586364061
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_202
timestamp 1586364061
transform 1 0 19688 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _241_
timestamp 1586364061
transform 1 0 20056 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_209
timestamp 1586364061
transform 1 0 20332 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_221
timestamp 1586364061
transform 1 0 21436 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_233
timestamp 1586364061
transform 1 0 22540 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_241
timestamp 1586364061
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use scs8hd_buf_2  _266_
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__266__A
timestamp 1586364061
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_259
timestamp 1586364061
transform 1 0 24932 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_263
timestamp 1586364061
transform 1 0 25300 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_275
timestamp 1586364061
transform 1 0 26404 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 1142 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 774 592
use scs8hd_nor2_4  _236_
timestamp 1586364061
transform 1 0 4784 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__234__B
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_49
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6348 0 -1 20128
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_32_53
timestamp 1586364061
transform 1 0 5980 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_6  FILLER_32_74
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_104
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_32_115
timestamp 1586364061
transform 1 0 11684 0 -1 20128
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_123
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_126
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_139
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_143
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_151
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_171
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_32_188
timestamp 1586364061
transform 1 0 18400 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19136 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_199
timestamp 1586364061
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_211
timestamp 1586364061
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_9
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_13
timestamp 1586364061
transform 1 0 2300 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_17
timestamp 1586364061
transform 1 0 2668 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_21
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_25
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_1  _164_
timestamp 1586364061
transform 1 0 4416 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3772 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_32
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_36
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use scs8hd_nor2_4  _239_
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__B
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_40
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_39
timestamp 1586364061
transform 1 0 4692 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_43
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_46
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_34_50
timestamp 1586364061
transform 1 0 5704 0 -1 21216
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6440 0 -1 21216
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_73
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_77
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_69
timestamp 1586364061
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_73
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_77
timestamp 1586364061
transform 1 0 8188 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_94
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_90
timestamp 1586364061
transform 1 0 9384 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_100
timestamp 1586364061
transform 1 0 10304 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_97
timestamp 1586364061
transform 1 0 10028 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_107
timestamp 1586364061
transform 1 0 10948 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_111
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 774 592
use scs8hd_decap_8  FILLER_34_110
timestamp 1586364061
transform 1 0 11224 0 -1 21216
box -38 -48 774 592
use scs8hd_nor2_4  _220_
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__220__A
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__220__B
timestamp 1586364061
transform 1 0 12604 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_121
timestamp 1586364061
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_127
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_118
timestamp 1586364061
transform 1 0 11960 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_34_128
timestamp 1586364061
transform 1 0 12880 0 -1 21216
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13064 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_134
timestamp 1586364061
transform 1 0 13432 0 -1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14996 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_154
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_158
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_162
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17388 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_172
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_176
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_169
timestamp 1586364061
transform 1 0 16652 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_173
timestamp 1586364061
transform 1 0 17020 0 -1 21216
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_187
timestamp 1586364061
transform 1 0 18308 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_191
timestamp 1586364061
transform 1 0 18676 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_186
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_198
timestamp 1586364061
transform 1 0 19320 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_202
timestamp 1586364061
transform 1 0 19688 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_198
timestamp 1586364061
transform 1 0 19320 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_214
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_210
timestamp 1586364061
transform 1 0 20424 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_226
timestamp 1586364061
transform 1 0 21896 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_238
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_2  _255_
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__255__A
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_11
timestamp 1586364061
transform 1 0 2116 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_23
timestamp 1586364061
transform 1 0 3220 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_35
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_40
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8740 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_79
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_92
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_96
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_109
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_35_115
timestamp 1586364061
transform 1 0 11684 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_119
timestamp 1586364061
transform 1 0 12052 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_139
timestamp 1586364061
transform 1 0 13892 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_152
timestamp 1586364061
transform 1 0 15088 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_169
timestamp 1586364061
transform 1 0 16652 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_173
timestamp 1586364061
transform 1 0 17020 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_177
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_191
timestamp 1586364061
transform 1 0 18676 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_203
timestamp 1586364061
transform 1 0 19780 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_215
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_227
timestamp 1586364061
transform 1 0 21988 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_35_239
timestamp 1586364061
transform 1 0 23092 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_243
timestamp 1586364061
transform 1 0 23460 0 1 21216
box -38 -48 130 592
use scs8hd_buf_2  _264_
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_253
timestamp 1586364061
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__264__A
timestamp 1586364061
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_259
timestamp 1586364061
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_263
timestamp 1586364061
transform 1 0 25300 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_275
timestamp 1586364061
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__252__A
timestamp 1586364061
transform 1 0 1564 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_7
timestamp 1586364061
transform 1 0 1748 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_19
timestamp 1586364061
transform 1 0 2852 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_conb_1  _240_
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_47
timestamp 1586364061
transform 1 0 5428 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6164 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_58
timestamp 1586364061
transform 1 0 6440 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_8  FILLER_36_75
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_85
timestamp 1586364061
transform 1 0 8924 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_90
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10948 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_109
timestamp 1586364061
transform 1 0 11132 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_116
timestamp 1586364061
transform 1 0 11776 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_36_124
timestamp 1586364061
transform 1 0 12512 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_128
timestamp 1586364061
transform 1 0 12880 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_4  FILLER_36_139
timestamp 1586364061
transform 1 0 13892 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_6  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 22304
box -38 -48 866 592
use scs8hd_fill_1  FILLER_36_160
timestamp 1586364061
transform 1 0 15824 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_170
timestamp 1586364061
transform 1 0 16744 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_182
timestamp 1586364061
transform 1 0 17848 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_194
timestamp 1586364061
transform 1 0 18952 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_206
timestamp 1586364061
transform 1 0 20056 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_buf_2  _254_
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__254__A
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_11
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_23
timestamp 1586364061
transform 1 0 3220 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_35
timestamp 1586364061
transform 1 0 4324 0 1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_47
timestamp 1586364061
transform 1 0 5428 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7084 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_76
timestamp 1586364061
transform 1 0 8096 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_80
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_83
timestamp 1586364061
transform 1 0 8740 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_97
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_101
timestamp 1586364061
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_108
timestamp 1586364061
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_112
timestamp 1586364061
transform 1 0 11408 0 1 22304
box -38 -48 222 592
use scs8hd_buf_1  _153_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_116
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_37_126
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_137
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_141
timestamp 1586364061
transform 1 0 14076 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14444 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14904 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_148
timestamp 1586364061
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_152
timestamp 1586364061
transform 1 0 15088 0 1 22304
box -38 -48 406 592
use scs8hd_conb_1  _247_
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_161
timestamp 1586364061
transform 1 0 15916 0 1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_169
timestamp 1586364061
transform 1 0 16652 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_175
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__261__A
timestamp 1586364061
transform 1 0 18216 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_188
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_200
timestamp 1586364061
transform 1 0 19504 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_212
timestamp 1586364061
transform 1 0 20608 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_224
timestamp 1586364061
transform 1 0 21712 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_236
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__263__A
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_buf_2  _252_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_64
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_70
timestamp 1586364061
transform 1 0 7544 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_74
timestamp 1586364061
transform 1 0 7912 0 -1 23392
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_113
timestamp 1586364061
transform 1 0 11500 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_124
timestamp 1586364061
transform 1 0 12512 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_132
timestamp 1586364061
transform 1 0 13248 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_138
timestamp 1586364061
transform 1 0 13800 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_150
timestamp 1586364061
transform 1 0 14904 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_159
timestamp 1586364061
transform 1 0 15732 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_167
timestamp 1586364061
transform 1 0 16468 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_173
timestamp 1586364061
transform 1 0 17020 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_2  _261_
timestamp 1586364061
transform 1 0 18032 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_38_181
timestamp 1586364061
transform 1 0 17756 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_188
timestamp 1586364061
transform 1 0 18400 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_200
timestamp 1586364061
transform 1 0 19504 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_212
timestamp 1586364061
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _263_
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_buf_2  _253_
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__253__A
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_23
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_35
timestamp 1586364061
transform 1 0 4324 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_47
timestamp 1586364061
transform 1 0 5428 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_1  _233_
timestamp 1586364061
transform 1 0 8924 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_82
timestamp 1586364061
transform 1 0 8648 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_88
timestamp 1586364061
transform 1 0 9200 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_conb_1  _244_
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_92
timestamp 1586364061
transform 1 0 9568 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_99
timestamp 1586364061
transform 1 0 10212 0 1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_101
timestamp 1586364061
transform 1 0 10396 0 -1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10580 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11592 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_105
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_106
timestamp 1586364061
transform 1 0 10856 0 -1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_116
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_126
timestamp 1586364061
transform 1 0 12696 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_130
timestamp 1586364061
transform 1 0 13064 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _287_
timestamp 1586364061
transform 1 0 14352 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__287__A
timestamp 1586364061
transform 1 0 14904 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_142
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_148
timestamp 1586364061
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_152
timestamp 1586364061
transform 1 0 15088 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _286_
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_160
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_166
timestamp 1586364061
transform 1 0 16376 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 590 592
use scs8hd_buf_2  _285_
timestamp 1586364061
transform 1 0 16928 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__286__A
timestamp 1586364061
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__285__A
timestamp 1586364061
transform 1 0 16928 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_170
timestamp 1586364061
transform 1 0 16744 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_174
timestamp 1586364061
transform 1 0 17112 0 1 23392
box -38 -48 590 592
use scs8hd_decap_8  FILLER_40_176
timestamp 1586364061
transform 1 0 17296 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _280_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _284_
timestamp 1586364061
transform 1 0 18032 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__284__A
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__280__A
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_180
timestamp 1586364061
transform 1 0 17664 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_192
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_188
timestamp 1586364061
transform 1 0 18400 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_39_204
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_200
timestamp 1586364061
transform 1 0 19504 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _283_
timestamp 1586364061
transform 1 0 20148 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__283__A
timestamp 1586364061
transform 1 0 20700 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_211
timestamp 1586364061
transform 1 0 20516 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_215
timestamp 1586364061
transform 1 0 20884 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_212
timestamp 1586364061
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _281_
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _282_
timestamp 1586364061
transform 1 0 21252 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__282__A
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_223
timestamp 1586364061
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__281__A
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_235
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_239
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _262_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__262__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 3330 0 3386 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 4250 0 4306 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 5262 0 5318 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 6182 0 6238 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 7194 0 7250 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 8114 0 8170 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 9126 0 9182 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 478 0 534 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal3 s 0 2048 480 2168 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal3 s 0 3408 480 3528 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal3 s 0 16056 480 16176 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal3 s 0 21632 480 21752 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal3 s 0 24488 480 24608 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal3 s 0 27208 480 27328 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal3 s 27520 2048 28000 2168 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal3 s 27520 3408 28000 3528 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal3 s 27520 4768 28000 4888 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal3 s 27520 6264 28000 6384 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal3 s 27520 8984 28000 9104 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal3 s 27520 13200 28000 13320 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal3 s 27520 16056 28000 16176 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal3 s 27520 17416 28000 17536 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal3 s 27520 18776 28000 18896 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 27520 21632 28000 21752 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal3 s 27520 22992 28000 23112 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal3 s 27520 24488 28000 24608 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 27520 25848 28000 25968 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal3 s 27520 27208 28000 27328 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 11058 0 11114 480 6 chany_bottom_in[0]
port 45 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[1]
port 46 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[2]
port 47 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[3]
port 48 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[4]
port 49 nsew default input
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_in[5]
port 50 nsew default input
rlabel metal2 s 16854 0 16910 480 6 chany_bottom_in[6]
port 51 nsew default input
rlabel metal2 s 17774 0 17830 480 6 chany_bottom_in[7]
port 52 nsew default input
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_in[8]
port 53 nsew default input
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[0]
port 54 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[1]
port 55 nsew default tristate
rlabel metal2 s 21638 0 21694 480 6 chany_bottom_out[2]
port 56 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[3]
port 57 nsew default tristate
rlabel metal2 s 23570 0 23626 480 6 chany_bottom_out[4]
port 58 nsew default tristate
rlabel metal2 s 24582 0 24638 480 6 chany_bottom_out[5]
port 59 nsew default tristate
rlabel metal2 s 25502 0 25558 480 6 chany_bottom_out[6]
port 60 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[7]
port 61 nsew default tristate
rlabel metal2 s 27434 0 27490 480 6 chany_bottom_out[8]
port 62 nsew default tristate
rlabel metal2 s 662 27520 718 28000 6 chany_top_in[0]
port 63 nsew default input
rlabel metal2 s 2042 27520 2098 28000 6 chany_top_in[1]
port 64 nsew default input
rlabel metal2 s 3422 27520 3478 28000 6 chany_top_in[2]
port 65 nsew default input
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[3]
port 66 nsew default input
rlabel metal2 s 6182 27520 6238 28000 6 chany_top_in[4]
port 67 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[5]
port 68 nsew default input
rlabel metal2 s 9034 27520 9090 28000 6 chany_top_in[6]
port 69 nsew default input
rlabel metal2 s 10414 27520 10470 28000 6 chany_top_in[7]
port 70 nsew default input
rlabel metal2 s 11794 27520 11850 28000 6 chany_top_in[8]
port 71 nsew default input
rlabel metal2 s 16026 27520 16082 28000 6 chany_top_out[0]
port 72 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 18786 27520 18842 28000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 20166 27520 20222 28000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 21638 27520 21694 28000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 23018 27520 23074 28000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 24398 27520 24454 28000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 25778 27520 25834 28000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 27158 27520 27214 28000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 10046 0 10102 480 6 data_in
port 81 nsew default input
rlabel metal2 s 2318 0 2374 480 6 enable
port 82 nsew default input
rlabel metal3 s 0 14696 480 14816 6 left_bottom_grid_pin_12_
port 83 nsew default input
rlabel metal3 s 0 688 480 808 6 left_top_grid_pin_10_
port 84 nsew default input
rlabel metal3 s 27520 14696 28000 14816 6 right_bottom_grid_pin_12_
port 85 nsew default input
rlabel metal3 s 27520 688 28000 808 6 right_top_grid_pin_10_
port 86 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 top_left_grid_pin_13_
port 87 nsew default input
rlabel metal2 s 14646 27520 14702 28000 6 top_right_grid_pin_11_
port 88 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 89 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 90 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
