VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga_core
  CLASS BLOCK ;
  FOREIGN fpga_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 1058.520 BY 1146.320 ;
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 96.520 51.880 97.120 ;
    END
  END Test_en
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1007.080 102.640 1009.480 103.240 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 944.480 51.880 945.080 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 201.920 51.880 202.520 ;
    END
  END clk
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.150 1101.720 129.430 1104.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 542.230 44.120 542.510 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[10]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 568.910 44.120 569.190 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[11]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 595.590 44.120 595.870 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[12]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 622.270 44.120 622.550 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[13]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 648.950 44.120 649.230 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[14]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 675.630 44.120 675.910 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[15]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 308.000 51.880 308.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[16]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 626.240 51.880 626.840 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[17]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 288.770 1101.720 289.050 1104.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1007.080 455.560 1009.480 456.160 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1007.080 573.200 1009.480 573.800 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.450 44.120 62.730 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.670 44.120 88.950 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.350 44.120 115.630 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[6]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 142.030 44.120 142.310 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[7]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 168.710 44.120 168.990 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[8]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 195.390 44.120 195.670 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[9]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 448.850 1101.720 449.130 1104.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 702.310 44.120 702.590 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[10]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 728.990 44.120 729.270 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[11]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 755.670 44.120 755.950 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[12]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 782.350 44.120 782.630 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[13]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 809.030 44.120 809.310 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[14]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 835.710 44.120 835.990 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[15]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 414.080 51.880 414.680 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[16]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 732.320 51.880 732.920 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[17]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 608.930 1101.720 609.210 1104.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1007.080 691.520 1009.480 692.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1007.080 809.160 1009.480 809.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.070 44.120 222.350 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 248.750 44.120 249.030 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.430 44.120 275.710 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[6]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.110 44.120 302.390 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[7]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 328.790 44.120 329.070 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[8]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 355.470 44.120 355.750 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[9]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 769.010 1101.720 769.290 1104.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 862.390 44.120 862.670 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[10]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 889.070 44.120 889.350 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[11]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 915.750 44.120 916.030 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[12]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.430 44.120 942.710 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[13]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 969.110 44.120 969.390 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[14]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.790 44.120 996.070 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[15]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 520.160 51.880 520.760 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[16]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 838.400 51.880 839.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[17]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 929.090 1101.720 929.370 1104.120 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1007.080 926.800 1009.480 927.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1007.080 1044.440 1009.480 1045.040 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 382.150 44.120 382.430 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 408.830 44.120 409.110 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 435.510 44.120 435.790 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[6]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 462.190 44.120 462.470 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[7]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 488.870 44.120 489.150 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[8]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 515.550 44.120 515.830 46.520 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1007.080 337.920 1009.480 338.520 ;
    END
  END prog_clk
  PIN sc_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1007.080 220.280 1009.480 220.880 ;
    END
  END sc_head
  PIN sc_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 49.480 1050.560 51.880 1051.160 ;
    END
  END sc_tail
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 1033.520 45.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 1058.520 20.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 103.555 88.065 953.800 1044.995 ;
      LAYER met1 ;
        RECT 62.430 58.440 996.090 1082.780 ;
      LAYER met2 ;
        RECT 62.460 1101.440 128.870 1101.720 ;
        RECT 129.710 1101.440 288.490 1101.720 ;
        RECT 289.330 1101.440 448.570 1101.720 ;
        RECT 449.410 1101.440 608.650 1101.720 ;
        RECT 609.490 1101.440 768.730 1101.720 ;
        RECT 769.570 1101.440 928.810 1101.720 ;
        RECT 929.650 1101.440 1006.650 1101.720 ;
        RECT 62.460 46.800 1006.650 1101.440 ;
        RECT 63.010 46.520 88.390 46.800 ;
        RECT 89.230 46.520 115.070 46.800 ;
        RECT 115.910 46.520 141.750 46.800 ;
        RECT 142.590 46.520 168.430 46.800 ;
        RECT 169.270 46.520 195.110 46.800 ;
        RECT 195.950 46.520 221.790 46.800 ;
        RECT 222.630 46.520 248.470 46.800 ;
        RECT 249.310 46.520 275.150 46.800 ;
        RECT 275.990 46.520 301.830 46.800 ;
        RECT 302.670 46.520 328.510 46.800 ;
        RECT 329.350 46.520 355.190 46.800 ;
        RECT 356.030 46.520 381.870 46.800 ;
        RECT 382.710 46.520 408.550 46.800 ;
        RECT 409.390 46.520 435.230 46.800 ;
        RECT 436.070 46.520 461.910 46.800 ;
        RECT 462.750 46.520 488.590 46.800 ;
        RECT 489.430 46.520 515.270 46.800 ;
        RECT 516.110 46.520 541.950 46.800 ;
        RECT 542.790 46.520 568.630 46.800 ;
        RECT 569.470 46.520 595.310 46.800 ;
        RECT 596.150 46.520 621.990 46.800 ;
        RECT 622.830 46.520 648.670 46.800 ;
        RECT 649.510 46.520 675.350 46.800 ;
        RECT 676.190 46.520 702.030 46.800 ;
        RECT 702.870 46.520 728.710 46.800 ;
        RECT 729.550 46.520 755.390 46.800 ;
        RECT 756.230 46.520 782.070 46.800 ;
        RECT 782.910 46.520 808.750 46.800 ;
        RECT 809.590 46.520 835.430 46.800 ;
        RECT 836.270 46.520 862.110 46.800 ;
        RECT 862.950 46.520 888.790 46.800 ;
        RECT 889.630 46.520 915.470 46.800 ;
        RECT 916.310 46.520 942.150 46.800 ;
        RECT 942.990 46.520 968.830 46.800 ;
        RECT 969.670 46.520 995.510 46.800 ;
        RECT 996.350 46.520 1006.650 46.800 ;
      LAYER met3 ;
        RECT 51.880 1051.560 1007.080 1065.985 ;
        RECT 52.280 1050.160 1007.080 1051.560 ;
        RECT 51.880 1045.440 1007.080 1050.160 ;
        RECT 51.880 1044.040 1006.680 1045.440 ;
        RECT 51.880 945.480 1007.080 1044.040 ;
        RECT 52.280 944.080 1007.080 945.480 ;
        RECT 51.880 927.800 1007.080 944.080 ;
        RECT 51.880 926.400 1006.680 927.800 ;
        RECT 51.880 839.400 1007.080 926.400 ;
        RECT 52.280 838.000 1007.080 839.400 ;
        RECT 51.880 810.160 1007.080 838.000 ;
        RECT 51.880 808.760 1006.680 810.160 ;
        RECT 51.880 733.320 1007.080 808.760 ;
        RECT 52.280 731.920 1007.080 733.320 ;
        RECT 51.880 692.520 1007.080 731.920 ;
        RECT 51.880 691.120 1006.680 692.520 ;
        RECT 51.880 627.240 1007.080 691.120 ;
        RECT 52.280 625.840 1007.080 627.240 ;
        RECT 51.880 574.200 1007.080 625.840 ;
        RECT 51.880 572.800 1006.680 574.200 ;
        RECT 51.880 521.160 1007.080 572.800 ;
        RECT 52.280 519.760 1007.080 521.160 ;
        RECT 51.880 456.560 1007.080 519.760 ;
        RECT 51.880 455.160 1006.680 456.560 ;
        RECT 51.880 415.080 1007.080 455.160 ;
        RECT 52.280 413.680 1007.080 415.080 ;
        RECT 51.880 338.920 1007.080 413.680 ;
        RECT 51.880 337.520 1006.680 338.920 ;
        RECT 51.880 309.000 1007.080 337.520 ;
        RECT 52.280 307.600 1007.080 309.000 ;
        RECT 51.880 221.280 1007.080 307.600 ;
        RECT 51.880 219.880 1006.680 221.280 ;
        RECT 51.880 202.920 1007.080 219.880 ;
        RECT 52.280 201.520 1007.080 202.920 ;
        RECT 51.880 103.640 1007.080 201.520 ;
        RECT 51.880 102.240 1006.680 103.640 ;
        RECT 51.880 97.520 1007.080 102.240 ;
        RECT 52.280 96.120 1007.080 97.520 ;
        RECT 51.880 85.095 1007.080 96.120 ;
      LAYER met4 ;
        RECT 0.000 0.000 1058.520 1146.320 ;
      LAYER met5 ;
        RECT 0.000 79.200 1058.520 1146.320 ;
  END
END fpga_core
END LIBRARY

