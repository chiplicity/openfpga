VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_io_bottom
  CLASS BLOCK ;
  FOREIGN grid_io_bottom ;
  ORIGIN 0.000 0.000 ;
  SIZE 2120.000 BY 50.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 2.400 9.480 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 2.400 15.600 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 2.400 ;
    END
  END address[3]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 12.280 2120.000 12.880 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 4.120 2120.000 4.720 ;
    END
  END enable
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 20.440 2120.000 21.040 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 2.400 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 29.280 2120.000 29.880 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 2.400 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 741.610 0.000 741.890 2.400 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 953.670 0.000 953.950 2.400 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 176.730 47.600 177.010 50.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 45.600 2120.000 46.200 ;
    END
  END top_width_0_height_0__pin_10_
  PIN top_width_0_height_0__pin_11_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 2.400 34.640 ;
    END
  END top_width_0_height_0__pin_11_
  PIN top_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 2.400 40.760 ;
    END
  END top_width_0_height_0__pin_12_
  PIN top_width_0_height_0__pin_13_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2013.970 0.000 2014.250 2.400 ;
    END
  END top_width_0_height_0__pin_13_
  PIN top_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1943.130 47.600 1943.410 50.000 ;
    END
  END top_width_0_height_0__pin_14_
  PIN top_width_0_height_0__pin_15_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 2.400 46.880 ;
    END
  END top_width_0_height_0__pin_15_
  PIN top_width_0_height_0__pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 530.010 47.600 530.290 50.000 ;
    END
  END top_width_0_height_0__pin_1_
  PIN top_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1165.730 0.000 1166.010 2.400 ;
    END
  END top_width_0_height_0__pin_2_
  PIN top_width_0_height_0__pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 883.290 47.600 883.570 50.000 ;
    END
  END top_width_0_height_0__pin_3_
  PIN top_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2117.600 37.440 2120.000 38.040 ;
    END
  END top_width_0_height_0__pin_4_
  PIN top_width_0_height_0__pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1377.790 0.000 1378.070 2.400 ;
    END
  END top_width_0_height_0__pin_5_
  PIN top_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1589.850 0.000 1590.130 2.400 ;
    END
  END top_width_0_height_0__pin_6_
  PIN top_width_0_height_0__pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1801.910 0.000 1802.190 2.400 ;
    END
  END top_width_0_height_0__pin_7_
  PIN top_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1236.570 47.600 1236.850 50.000 ;
    END
  END top_width_0_height_0__pin_8_
  PIN top_width_0_height_0__pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1589.850 47.600 1590.130 50.000 ;
    END
  END top_width_0_height_0__pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 358.055 10.640 359.655 38.320 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 711.385 10.640 712.985 38.320 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2114.160 38.165 ;
      LAYER met1 ;
        RECT 0.530 10.640 2118.230 41.100 ;
      LAYER met2 ;
        RECT 0.090 47.320 176.450 48.010 ;
        RECT 177.290 47.320 529.730 48.010 ;
        RECT 530.570 47.320 883.010 48.010 ;
        RECT 883.850 47.320 1236.290 48.010 ;
        RECT 1237.130 47.320 1589.570 48.010 ;
        RECT 1590.410 47.320 1942.850 48.010 ;
        RECT 1943.690 47.320 2118.670 48.010 ;
        RECT 0.090 2.680 2118.670 47.320 ;
        RECT 0.090 0.155 105.610 2.680 ;
        RECT 106.450 0.155 317.210 2.680 ;
        RECT 318.050 0.155 529.270 2.680 ;
        RECT 530.110 0.155 741.330 2.680 ;
        RECT 742.170 0.155 953.390 2.680 ;
        RECT 954.230 0.155 1165.450 2.680 ;
        RECT 1166.290 0.155 1377.510 2.680 ;
        RECT 1378.350 0.155 1589.570 2.680 ;
        RECT 1590.410 0.155 1801.630 2.680 ;
        RECT 1802.470 0.155 2013.690 2.680 ;
        RECT 2014.530 0.155 2118.670 2.680 ;
      LAYER met3 ;
        RECT 0.065 37.040 2117.200 38.245 ;
        RECT 0.065 35.040 2118.695 37.040 ;
        RECT 2.800 33.640 2118.695 35.040 ;
        RECT 0.065 30.280 2118.695 33.640 ;
        RECT 0.065 28.920 2117.200 30.280 ;
        RECT 2.800 28.880 2117.200 28.920 ;
        RECT 2.800 27.520 2118.695 28.880 ;
        RECT 0.065 22.120 2118.695 27.520 ;
        RECT 2.800 21.440 2118.695 22.120 ;
        RECT 2.800 20.720 2117.200 21.440 ;
        RECT 0.065 20.040 2117.200 20.720 ;
        RECT 0.065 16.000 2118.695 20.040 ;
        RECT 2.800 14.600 2118.695 16.000 ;
        RECT 0.065 13.280 2118.695 14.600 ;
        RECT 0.065 11.880 2117.200 13.280 ;
        RECT 0.065 9.880 2118.695 11.880 ;
        RECT 2.800 8.480 2118.695 9.880 ;
        RECT 0.065 5.120 2118.695 8.480 ;
        RECT 0.065 3.760 2117.200 5.120 ;
        RECT 2.800 3.720 2117.200 3.760 ;
        RECT 2.800 2.360 2118.695 3.720 ;
        RECT 0.065 0.175 2118.695 2.360 ;
      LAYER met4 ;
        RECT 0.295 10.240 357.655 38.320 ;
        RECT 360.055 10.240 710.985 38.320 ;
        RECT 713.385 10.240 2118.465 38.320 ;
        RECT 0.295 9.015 2118.465 10.240 ;
  END
END grid_io_bottom
END LIBRARY

