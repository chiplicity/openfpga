magic
tech sky130A
magscale 1 2
timestamp 1605003126
<< locali >>
rect 9873 19159 9907 19329
rect 24501 7191 24535 7361
<< viali >>
rect 16589 25449 16623 25483
rect 20177 25449 20211 25483
rect 21649 25449 21683 25483
rect 22845 25449 22879 25483
rect 24777 25449 24811 25483
rect 16405 25313 16439 25347
rect 18889 25313 18923 25347
rect 19993 25313 20027 25347
rect 21465 25313 21499 25347
rect 22661 25313 22695 25347
rect 24593 25313 24627 25347
rect 19073 25177 19107 25211
rect 19441 25109 19475 25143
rect 17049 24905 17083 24939
rect 23397 24837 23431 24871
rect 15945 24769 15979 24803
rect 14197 24701 14231 24735
rect 15301 24701 15335 24735
rect 16865 24701 16899 24735
rect 17417 24701 17451 24735
rect 18061 24701 18095 24735
rect 19165 24701 19199 24735
rect 20269 24701 20303 24735
rect 20821 24701 20855 24735
rect 21373 24701 21407 24735
rect 22477 24701 22511 24735
rect 23029 24701 23063 24735
rect 24593 24701 24627 24735
rect 25145 24701 25179 24735
rect 14381 24565 14415 24599
rect 14749 24565 14783 24599
rect 15485 24565 15519 24599
rect 16405 24565 16439 24599
rect 17785 24565 17819 24599
rect 18245 24565 18279 24599
rect 18981 24565 19015 24599
rect 19349 24565 19383 24599
rect 19993 24565 20027 24599
rect 20453 24565 20487 24599
rect 21557 24565 21591 24599
rect 21925 24565 21959 24599
rect 22385 24565 22419 24599
rect 22661 24565 22695 24599
rect 24409 24565 24443 24599
rect 24777 24565 24811 24599
rect 13093 24361 13127 24395
rect 14289 24361 14323 24395
rect 17969 24361 18003 24395
rect 19349 24361 19383 24395
rect 21097 24361 21131 24395
rect 22569 24361 22603 24395
rect 23673 24361 23707 24395
rect 15669 24293 15703 24327
rect 14105 24225 14139 24259
rect 15761 24225 15795 24259
rect 18061 24225 18095 24259
rect 19165 24225 19199 24259
rect 20913 24225 20947 24259
rect 22385 24225 22419 24259
rect 23489 24225 23523 24259
rect 24593 24225 24627 24259
rect 15945 24157 15979 24191
rect 18153 24157 18187 24191
rect 18613 24089 18647 24123
rect 15301 24021 15335 24055
rect 16681 24021 16715 24055
rect 17417 24021 17451 24055
rect 17601 24021 17635 24055
rect 24777 24021 24811 24055
rect 12817 23817 12851 23851
rect 16037 23817 16071 23851
rect 16405 23817 16439 23851
rect 17693 23817 17727 23851
rect 20729 23817 20763 23851
rect 22661 23817 22695 23851
rect 16865 23681 16899 23715
rect 12633 23613 12667 23647
rect 14105 23613 14139 23647
rect 16589 23613 16623 23647
rect 18061 23613 18095 23647
rect 18328 23613 18362 23647
rect 20545 23613 20579 23647
rect 21097 23613 21131 23647
rect 22477 23613 22511 23647
rect 24593 23613 24627 23647
rect 25145 23613 25179 23647
rect 13277 23545 13311 23579
rect 14350 23545 14384 23579
rect 19993 23545 20027 23579
rect 22385 23545 22419 23579
rect 13553 23477 13587 23511
rect 14013 23477 14047 23511
rect 15485 23477 15519 23511
rect 19441 23477 19475 23511
rect 21557 23477 21591 23511
rect 23029 23477 23063 23511
rect 23857 23477 23891 23511
rect 24409 23477 24443 23511
rect 24777 23477 24811 23511
rect 12449 23273 12483 23307
rect 14657 23273 14691 23307
rect 17693 23273 17727 23307
rect 18981 23273 19015 23307
rect 18337 23205 18371 23239
rect 22753 23205 22787 23239
rect 24041 23205 24075 23239
rect 10692 23137 10726 23171
rect 13277 23137 13311 23171
rect 15117 23137 15151 23171
rect 15752 23137 15786 23171
rect 19533 23137 19567 23171
rect 21281 23137 21315 23171
rect 22477 23137 22511 23171
rect 23765 23137 23799 23171
rect 25053 23137 25087 23171
rect 10425 23069 10459 23103
rect 13369 23069 13403 23103
rect 13553 23069 13587 23103
rect 15485 23069 15519 23103
rect 18429 23069 18463 23103
rect 18613 23069 18647 23103
rect 19809 23069 19843 23103
rect 21373 23069 21407 23103
rect 21465 23069 21499 23103
rect 22293 23069 22327 23103
rect 17969 23001 18003 23035
rect 10241 22933 10275 22967
rect 11805 22933 11839 22967
rect 12725 22933 12759 22967
rect 12909 22933 12943 22967
rect 14105 22933 14139 22967
rect 16865 22933 16899 22967
rect 20913 22933 20947 22967
rect 21925 22933 21959 22967
rect 25237 22933 25271 22967
rect 10609 22729 10643 22763
rect 10793 22729 10827 22763
rect 11897 22729 11931 22763
rect 12265 22729 12299 22763
rect 16865 22729 16899 22763
rect 17509 22729 17543 22763
rect 17877 22729 17911 22763
rect 21005 22729 21039 22763
rect 23489 22729 23523 22763
rect 25881 22729 25915 22763
rect 11253 22593 11287 22627
rect 11437 22593 11471 22627
rect 14933 22593 14967 22627
rect 18613 22593 18647 22627
rect 18981 22593 19015 22627
rect 21373 22593 21407 22627
rect 22017 22593 22051 22627
rect 22109 22593 22143 22627
rect 23949 22593 23983 22627
rect 10333 22525 10367 22559
rect 11161 22525 11195 22559
rect 12449 22525 12483 22559
rect 12716 22525 12750 22559
rect 19073 22525 19107 22559
rect 19340 22525 19374 22559
rect 21925 22525 21959 22559
rect 22569 22525 22603 22559
rect 23673 22525 23707 22559
rect 24409 22525 24443 22559
rect 24961 22525 24995 22559
rect 25513 22525 25547 22559
rect 9689 22457 9723 22491
rect 15178 22457 15212 22491
rect 9781 22389 9815 22423
rect 13829 22389 13863 22423
rect 14381 22389 14415 22423
rect 14749 22389 14783 22423
rect 16313 22389 16347 22423
rect 18061 22389 18095 22423
rect 20453 22389 20487 22423
rect 21557 22389 21591 22423
rect 22937 22389 22971 22423
rect 25145 22389 25179 22423
rect 11069 22185 11103 22219
rect 12265 22185 12299 22219
rect 13001 22185 13035 22219
rect 16037 22185 16071 22219
rect 17325 22185 17359 22219
rect 19625 22185 19659 22219
rect 8585 22117 8619 22151
rect 13737 22117 13771 22151
rect 20269 22117 20303 22151
rect 9956 22049 9990 22083
rect 13645 22049 13679 22083
rect 15301 22049 15335 22083
rect 17233 22049 17267 22083
rect 19717 22049 19751 22083
rect 21169 22049 21203 22083
rect 23765 22049 23799 22083
rect 24041 22049 24075 22083
rect 25053 22049 25087 22083
rect 9689 21981 9723 22015
rect 13921 21981 13955 22015
rect 15577 21981 15611 22015
rect 17417 21981 17451 22015
rect 19901 21981 19935 22015
rect 20913 21981 20947 22015
rect 13277 21913 13311 21947
rect 16865 21913 16899 21947
rect 8217 21845 8251 21879
rect 9413 21845 9447 21879
rect 14473 21845 14507 21879
rect 14841 21845 14875 21879
rect 16497 21845 16531 21879
rect 18153 21845 18187 21879
rect 19073 21845 19107 21879
rect 19257 21845 19291 21879
rect 20637 21845 20671 21879
rect 22293 21845 22327 21879
rect 25237 21845 25271 21879
rect 12725 21641 12759 21675
rect 13277 21641 13311 21675
rect 14289 21641 14323 21675
rect 16313 21641 16347 21675
rect 19717 21641 19751 21675
rect 20085 21641 20119 21675
rect 22477 21641 22511 21675
rect 25053 21641 25087 21675
rect 12265 21573 12299 21607
rect 10609 21505 10643 21539
rect 11161 21505 11195 21539
rect 11253 21505 11287 21539
rect 13829 21505 13863 21539
rect 15485 21505 15519 21539
rect 16957 21505 16991 21539
rect 18705 21505 18739 21539
rect 19349 21505 19383 21539
rect 20453 21505 20487 21539
rect 24225 21505 24259 21539
rect 25513 21505 25547 21539
rect 8217 21437 8251 21471
rect 10241 21437 10275 21471
rect 13645 21437 13679 21471
rect 15209 21437 15243 21471
rect 15945 21437 15979 21471
rect 18429 21437 18463 21471
rect 20545 21437 20579 21471
rect 20812 21437 20846 21471
rect 23949 21437 23983 21471
rect 24685 21437 24719 21471
rect 25237 21437 25271 21471
rect 25973 21437 26007 21471
rect 8125 21369 8159 21403
rect 8484 21369 8518 21403
rect 14657 21369 14691 21403
rect 15301 21369 15335 21403
rect 17785 21369 17819 21403
rect 18521 21369 18555 21403
rect 9597 21301 9631 21335
rect 10701 21301 10735 21335
rect 11069 21301 11103 21335
rect 13093 21301 13127 21335
rect 13737 21301 13771 21335
rect 14841 21301 14875 21335
rect 16405 21301 16439 21335
rect 16773 21301 16807 21335
rect 16865 21301 16899 21335
rect 17417 21301 17451 21335
rect 18061 21301 18095 21335
rect 21925 21301 21959 21335
rect 23489 21301 23523 21335
rect 8217 21097 8251 21131
rect 10701 21097 10735 21131
rect 12909 21097 12943 21131
rect 14105 21097 14139 21131
rect 15945 21097 15979 21131
rect 17509 21097 17543 21131
rect 18061 21097 18095 21131
rect 18521 21097 18555 21131
rect 19625 21097 19659 21131
rect 20361 21097 20395 21131
rect 22661 21097 22695 21131
rect 23581 21097 23615 21131
rect 9505 21029 9539 21063
rect 15485 21029 15519 21063
rect 10057 20961 10091 20995
rect 11253 20961 11287 20995
rect 13461 20961 13495 20995
rect 14841 20961 14875 20995
rect 16396 20961 16430 20995
rect 18981 20961 19015 20995
rect 19073 20961 19107 20995
rect 21281 20961 21315 20995
rect 22477 20961 22511 20995
rect 23949 20961 23983 20995
rect 25145 20961 25179 20995
rect 8309 20893 8343 20927
rect 8493 20893 8527 20927
rect 10149 20893 10183 20927
rect 10241 20893 10275 20927
rect 11529 20893 11563 20927
rect 13553 20893 13587 20927
rect 13737 20893 13771 20927
rect 16129 20893 16163 20927
rect 19165 20893 19199 20927
rect 21373 20893 21407 20927
rect 21465 20893 21499 20927
rect 23121 20893 23155 20927
rect 24041 20893 24075 20927
rect 24225 20893 24259 20927
rect 7849 20825 7883 20859
rect 20729 20825 20763 20859
rect 9689 20757 9723 20791
rect 12541 20757 12575 20791
rect 13093 20757 13127 20791
rect 14565 20757 14599 20791
rect 14657 20757 14691 20791
rect 18613 20757 18647 20791
rect 20913 20757 20947 20791
rect 23489 20757 23523 20791
rect 25329 20757 25363 20791
rect 7941 20553 7975 20587
rect 9689 20553 9723 20587
rect 11069 20553 11103 20587
rect 17417 20553 17451 20587
rect 20913 20553 20947 20587
rect 21925 20553 21959 20587
rect 22661 20553 22695 20587
rect 23673 20553 23707 20587
rect 25053 20553 25087 20587
rect 25973 20553 26007 20587
rect 11437 20485 11471 20519
rect 20085 20485 20119 20519
rect 22385 20485 22419 20519
rect 10149 20417 10183 20451
rect 10241 20417 10275 20451
rect 10793 20417 10827 20451
rect 21557 20417 21591 20451
rect 24225 20417 24259 20451
rect 25421 20417 25455 20451
rect 9597 20349 9631 20383
rect 10057 20349 10091 20383
rect 12449 20349 12483 20383
rect 12705 20349 12739 20383
rect 14381 20349 14415 20383
rect 14933 20349 14967 20383
rect 18061 20349 18095 20383
rect 18317 20349 18351 20383
rect 20361 20349 20395 20383
rect 21281 20349 21315 20383
rect 22477 20349 22511 20383
rect 23029 20349 23063 20383
rect 24133 20349 24167 20383
rect 25237 20349 25271 20383
rect 9229 20281 9263 20315
rect 11897 20281 11931 20315
rect 14841 20281 14875 20315
rect 15178 20281 15212 20315
rect 16957 20281 16991 20315
rect 20821 20281 20855 20315
rect 21373 20281 21407 20315
rect 24685 20281 24719 20315
rect 8309 20213 8343 20247
rect 8677 20213 8711 20247
rect 12173 20213 12207 20247
rect 13829 20213 13863 20247
rect 16313 20213 16347 20247
rect 17877 20213 17911 20247
rect 19441 20213 19475 20247
rect 23489 20213 23523 20247
rect 24041 20213 24075 20247
rect 9873 20009 9907 20043
rect 10241 20009 10275 20043
rect 13185 20009 13219 20043
rect 16681 20009 16715 20043
rect 17233 20009 17267 20043
rect 17785 20009 17819 20043
rect 20729 20009 20763 20043
rect 22293 20009 22327 20043
rect 22937 20009 22971 20043
rect 24777 20009 24811 20043
rect 25329 20009 25363 20043
rect 10876 19941 10910 19975
rect 13829 19941 13863 19975
rect 17601 19941 17635 19975
rect 18245 19941 18279 19975
rect 19165 19941 19199 19975
rect 21180 19941 21214 19975
rect 23305 19941 23339 19975
rect 13737 19873 13771 19907
rect 15557 19873 15591 19907
rect 18153 19873 18187 19907
rect 19349 19873 19383 19907
rect 20913 19873 20947 19907
rect 23653 19873 23687 19907
rect 10609 19805 10643 19839
rect 14013 19805 14047 19839
rect 15301 19805 15335 19839
rect 18337 19805 18371 19839
rect 19625 19805 19659 19839
rect 23404 19805 23438 19839
rect 15025 19737 15059 19771
rect 11989 19669 12023 19703
rect 12817 19669 12851 19703
rect 13369 19669 13403 19703
rect 14749 19669 14783 19703
rect 18797 19669 18831 19703
rect 9045 19465 9079 19499
rect 11161 19465 11195 19499
rect 12909 19465 12943 19499
rect 14749 19465 14783 19499
rect 15393 19465 15427 19499
rect 16405 19465 16439 19499
rect 17417 19465 17451 19499
rect 20821 19465 20855 19499
rect 21833 19465 21867 19499
rect 23397 19465 23431 19499
rect 25053 19465 25087 19499
rect 9873 19329 9907 19363
rect 10701 19329 10735 19363
rect 15945 19329 15979 19363
rect 17049 19329 17083 19363
rect 18613 19329 18647 19363
rect 21465 19329 21499 19363
rect 7665 19261 7699 19295
rect 7573 19193 7607 19227
rect 7910 19193 7944 19227
rect 9689 19193 9723 19227
rect 13369 19261 13403 19295
rect 17785 19261 17819 19295
rect 18521 19261 18555 19295
rect 19073 19261 19107 19295
rect 19809 19261 19843 19295
rect 20729 19261 20763 19295
rect 22477 19261 22511 19295
rect 23029 19261 23063 19295
rect 23673 19261 23707 19295
rect 10517 19193 10551 19227
rect 11529 19193 11563 19227
rect 13277 19193 13311 19227
rect 13636 19193 13670 19227
rect 16773 19193 16807 19227
rect 18429 19193 18463 19227
rect 19441 19193 19475 19227
rect 20361 19193 20395 19227
rect 23918 19193 23952 19227
rect 9873 19125 9907 19159
rect 9965 19125 9999 19159
rect 10149 19125 10183 19159
rect 10609 19125 10643 19159
rect 11989 19125 12023 19159
rect 16313 19125 16347 19159
rect 16865 19125 16899 19159
rect 18061 19125 18095 19159
rect 21189 19125 21223 19159
rect 21281 19125 21315 19159
rect 22201 19125 22235 19159
rect 22661 19125 22695 19159
rect 12173 18921 12207 18955
rect 13461 18921 13495 18955
rect 15761 18921 15795 18955
rect 16865 18921 16899 18955
rect 19901 18921 19935 18955
rect 21649 18921 21683 18955
rect 22753 18921 22787 18955
rect 23489 18921 23523 18955
rect 23673 18921 23707 18955
rect 21189 18853 21223 18887
rect 9505 18785 9539 18819
rect 9956 18785 9990 18819
rect 12541 18785 12575 18819
rect 15669 18785 15703 18819
rect 17141 18785 17175 18819
rect 17601 18785 17635 18819
rect 19257 18785 19291 18819
rect 19349 18785 19383 18819
rect 21465 18785 21499 18819
rect 22569 18785 22603 18819
rect 23121 18785 23155 18819
rect 24041 18785 24075 18819
rect 25237 18785 25271 18819
rect 9689 18717 9723 18751
rect 12633 18717 12667 18751
rect 12725 18717 12759 18751
rect 14197 18717 14231 18751
rect 15853 18717 15887 18751
rect 17693 18717 17727 18751
rect 17877 18717 17911 18751
rect 18797 18717 18831 18751
rect 19533 18717 19567 18751
rect 24133 18717 24167 18751
rect 24225 18717 24259 18751
rect 7757 18649 7791 18683
rect 9321 18649 9355 18683
rect 11069 18649 11103 18683
rect 15301 18649 15335 18683
rect 16957 18649 16991 18683
rect 11989 18581 12023 18615
rect 13829 18581 13863 18615
rect 14657 18581 14691 18615
rect 15025 18581 15059 18615
rect 16405 18581 16439 18615
rect 17233 18581 17267 18615
rect 18429 18581 18463 18615
rect 18889 18581 18923 18615
rect 20269 18581 20303 18615
rect 20637 18581 20671 18615
rect 24777 18581 24811 18615
rect 25053 18581 25087 18615
rect 25421 18581 25455 18615
rect 10333 18377 10367 18411
rect 11437 18377 11471 18411
rect 11897 18377 11931 18411
rect 12265 18377 12299 18411
rect 13645 18377 13679 18411
rect 13829 18377 13863 18411
rect 15301 18377 15335 18411
rect 16405 18377 16439 18411
rect 19717 18377 19751 18411
rect 20729 18377 20763 18411
rect 22109 18377 22143 18411
rect 25605 18377 25639 18411
rect 14933 18309 14967 18343
rect 21373 18309 21407 18343
rect 9229 18241 9263 18275
rect 10977 18241 11011 18275
rect 14381 18241 14415 18275
rect 15853 18241 15887 18275
rect 15945 18241 15979 18275
rect 18337 18241 18371 18275
rect 23029 18241 23063 18275
rect 12449 18173 12483 18207
rect 13369 18173 13403 18207
rect 14289 18173 14323 18207
rect 15761 18173 15795 18207
rect 17785 18173 17819 18207
rect 21189 18173 21223 18207
rect 22293 18173 22327 18207
rect 23673 18173 23707 18207
rect 23940 18173 23974 18207
rect 9321 18105 9355 18139
rect 9873 18105 9907 18139
rect 10701 18105 10735 18139
rect 12725 18105 12759 18139
rect 16865 18105 16899 18139
rect 17509 18105 17543 18139
rect 18604 18105 18638 18139
rect 20361 18105 20395 18139
rect 22569 18105 22603 18139
rect 10241 18037 10275 18071
rect 10793 18037 10827 18071
rect 14197 18037 14231 18071
rect 15393 18037 15427 18071
rect 16957 18037 16991 18071
rect 21097 18037 21131 18071
rect 21833 18037 21867 18071
rect 23489 18037 23523 18071
rect 25053 18037 25087 18071
rect 9413 17833 9447 17867
rect 10425 17833 10459 17867
rect 12081 17833 12115 17867
rect 13093 17833 13127 17867
rect 13645 17833 13679 17867
rect 14657 17833 14691 17867
rect 15025 17833 15059 17867
rect 18153 17833 18187 17867
rect 19625 17833 19659 17867
rect 24501 17833 24535 17867
rect 25237 17833 25271 17867
rect 10885 17765 10919 17799
rect 14105 17765 14139 17799
rect 20177 17765 20211 17799
rect 10793 17697 10827 17731
rect 11989 17697 12023 17731
rect 12449 17697 12483 17731
rect 14013 17697 14047 17731
rect 15761 17697 15795 17731
rect 16017 17697 16051 17731
rect 18501 17697 18535 17731
rect 21180 17697 21214 17731
rect 23857 17697 23891 17731
rect 25053 17697 25087 17731
rect 10977 17629 11011 17663
rect 12541 17629 12575 17663
rect 12725 17629 12759 17663
rect 14197 17629 14231 17663
rect 18245 17629 18279 17663
rect 20913 17629 20947 17663
rect 23949 17629 23983 17663
rect 24133 17629 24167 17663
rect 11621 17561 11655 17595
rect 13461 17561 13495 17595
rect 17693 17561 17727 17595
rect 23029 17561 23063 17595
rect 23489 17561 23523 17595
rect 9965 17493 9999 17527
rect 15577 17493 15611 17527
rect 17141 17493 17175 17527
rect 20545 17493 20579 17527
rect 22293 17493 22327 17527
rect 23397 17493 23431 17527
rect 24961 17493 24995 17527
rect 10149 17289 10183 17323
rect 12173 17289 12207 17323
rect 14749 17289 14783 17323
rect 16037 17289 16071 17323
rect 20177 17289 20211 17323
rect 21649 17289 21683 17323
rect 22661 17289 22695 17323
rect 23489 17289 23523 17323
rect 25145 17289 25179 17323
rect 10793 17221 10827 17255
rect 17049 17221 17083 17255
rect 10425 17153 10459 17187
rect 11345 17153 11379 17187
rect 12449 17153 12483 17187
rect 16497 17153 16531 17187
rect 16589 17153 16623 17187
rect 17509 17153 17543 17187
rect 18889 17153 18923 17187
rect 24133 17153 24167 17187
rect 24225 17153 24259 17187
rect 24685 17153 24719 17187
rect 11069 17085 11103 17119
rect 15485 17085 15519 17119
rect 18613 17085 18647 17119
rect 20269 17085 20303 17119
rect 22293 17085 22327 17119
rect 22937 17085 22971 17119
rect 24041 17085 24075 17119
rect 25237 17085 25271 17119
rect 25973 17085 26007 17119
rect 12716 17017 12750 17051
rect 17877 17017 17911 17051
rect 19625 17017 19659 17051
rect 20514 17017 20548 17051
rect 25513 17017 25547 17051
rect 13829 16949 13863 16983
rect 14381 16949 14415 16983
rect 15853 16949 15887 16983
rect 16405 16949 16439 16983
rect 18245 16949 18279 16983
rect 18705 16949 18739 16983
rect 19257 16949 19291 16983
rect 22753 16949 22787 16983
rect 23673 16949 23707 16983
rect 10517 16745 10551 16779
rect 13185 16745 13219 16779
rect 13553 16745 13587 16779
rect 15117 16745 15151 16779
rect 15669 16745 15703 16779
rect 16681 16745 16715 16779
rect 17141 16745 17175 16779
rect 17233 16745 17267 16779
rect 18245 16745 18279 16779
rect 18613 16745 18647 16779
rect 19257 16745 19291 16779
rect 20361 16745 20395 16779
rect 20913 16745 20947 16779
rect 22293 16745 22327 16779
rect 24133 16745 24167 16779
rect 25053 16745 25087 16779
rect 25421 16745 25455 16779
rect 14105 16677 14139 16711
rect 16037 16677 16071 16711
rect 17601 16677 17635 16711
rect 19809 16677 19843 16711
rect 22017 16677 22051 16711
rect 11161 16609 11195 16643
rect 11428 16609 11462 16643
rect 14013 16609 14047 16643
rect 15485 16609 15519 16643
rect 19165 16609 19199 16643
rect 21281 16609 21315 16643
rect 22753 16609 22787 16643
rect 23020 16609 23054 16643
rect 25237 16609 25271 16643
rect 14197 16541 14231 16575
rect 16129 16541 16163 16575
rect 16313 16541 16347 16575
rect 17693 16541 17727 16575
rect 17877 16541 17911 16575
rect 19349 16541 19383 16575
rect 21373 16541 21407 16575
rect 21465 16541 21499 16575
rect 10885 16405 10919 16439
rect 12541 16405 12575 16439
rect 13645 16405 13679 16439
rect 14657 16405 14691 16439
rect 18797 16405 18831 16439
rect 20637 16405 20671 16439
rect 10793 16201 10827 16235
rect 11897 16201 11931 16235
rect 13737 16201 13771 16235
rect 17509 16201 17543 16235
rect 17785 16201 17819 16235
rect 21097 16201 21131 16235
rect 21649 16201 21683 16235
rect 23489 16201 23523 16235
rect 23673 16201 23707 16235
rect 25973 16201 26007 16235
rect 12265 16133 12299 16167
rect 18061 16133 18095 16167
rect 11253 16065 11287 16099
rect 11345 16065 11379 16099
rect 13001 16065 13035 16099
rect 16865 16065 16899 16099
rect 18521 16065 18555 16099
rect 18613 16065 18647 16099
rect 19073 16065 19107 16099
rect 22477 16065 22511 16099
rect 24133 16065 24167 16099
rect 24317 16065 24351 16099
rect 25421 16065 25455 16099
rect 14197 15997 14231 16031
rect 14464 15997 14498 16031
rect 16497 15997 16531 16031
rect 16681 15997 16715 16031
rect 18429 15997 18463 16031
rect 19717 15997 19751 16031
rect 22293 15997 22327 16031
rect 23121 15997 23155 16031
rect 25237 15997 25271 16031
rect 10333 15929 10367 15963
rect 11161 15929 11195 15963
rect 12909 15929 12943 15963
rect 19962 15929 19996 15963
rect 22201 15929 22235 15963
rect 24041 15929 24075 15963
rect 24777 15929 24811 15963
rect 10701 15861 10735 15895
rect 12449 15861 12483 15895
rect 12817 15861 12851 15895
rect 14013 15861 14047 15895
rect 15577 15861 15611 15895
rect 16129 15861 16163 15895
rect 19533 15861 19567 15895
rect 25053 15861 25087 15895
rect 12633 15657 12667 15691
rect 13093 15657 13127 15691
rect 13553 15657 13587 15691
rect 14197 15657 14231 15691
rect 14473 15657 14507 15691
rect 15761 15657 15795 15691
rect 17693 15657 17727 15691
rect 18153 15657 18187 15691
rect 18797 15657 18831 15691
rect 19257 15657 19291 15691
rect 21189 15657 21223 15691
rect 22845 15657 22879 15691
rect 23765 15657 23799 15691
rect 23949 15657 23983 15691
rect 10876 15589 10910 15623
rect 17325 15589 17359 15623
rect 19625 15589 19659 15623
rect 20729 15589 20763 15623
rect 12909 15521 12943 15555
rect 13461 15521 13495 15555
rect 16497 15521 16531 15555
rect 18061 15521 18095 15555
rect 19717 15521 19751 15555
rect 21465 15521 21499 15555
rect 21732 15521 21766 15555
rect 24317 15521 24351 15555
rect 24409 15521 24443 15555
rect 10609 15453 10643 15487
rect 13645 15453 13679 15487
rect 16589 15453 16623 15487
rect 16773 15453 16807 15487
rect 18245 15453 18279 15487
rect 19165 15453 19199 15487
rect 19901 15453 19935 15487
rect 20361 15453 20395 15487
rect 24501 15453 24535 15487
rect 14841 15385 14875 15419
rect 11989 15317 12023 15351
rect 16129 15317 16163 15351
rect 24961 15317 24995 15351
rect 10701 15113 10735 15147
rect 12265 15113 12299 15147
rect 15393 15113 15427 15147
rect 19901 15113 19935 15147
rect 23121 15113 23155 15147
rect 23857 15113 23891 15147
rect 25421 15113 25455 15147
rect 11897 15045 11931 15079
rect 16865 15045 16899 15079
rect 21465 15045 21499 15079
rect 12449 14977 12483 15011
rect 14381 14977 14415 15011
rect 14473 14977 14507 15011
rect 15485 14977 15519 15011
rect 18613 14977 18647 15011
rect 20361 14977 20395 15011
rect 20453 14977 20487 15011
rect 22109 14977 22143 15011
rect 22569 14977 22603 15011
rect 14933 14909 14967 14943
rect 19533 14909 19567 14943
rect 24041 14909 24075 14943
rect 11345 14841 11379 14875
rect 13829 14841 13863 14875
rect 14289 14841 14323 14875
rect 15730 14841 15764 14875
rect 18429 14841 18463 14875
rect 21005 14841 21039 14875
rect 21833 14841 21867 14875
rect 23489 14841 23523 14875
rect 24308 14841 24342 14875
rect 10241 14773 10275 14807
rect 11161 14773 11195 14807
rect 13185 14773 13219 14807
rect 13921 14773 13955 14807
rect 17417 14773 17451 14807
rect 17785 14773 17819 14807
rect 18061 14773 18095 14807
rect 18521 14773 18555 14807
rect 19073 14773 19107 14807
rect 20269 14773 20303 14807
rect 21281 14773 21315 14807
rect 21925 14773 21959 14807
rect 10609 14569 10643 14603
rect 11621 14569 11655 14603
rect 11989 14569 12023 14603
rect 12449 14569 12483 14603
rect 14105 14569 14139 14603
rect 15301 14569 15335 14603
rect 16773 14569 16807 14603
rect 17049 14569 17083 14603
rect 17693 14569 17727 14603
rect 19165 14569 19199 14603
rect 20269 14569 20303 14603
rect 20913 14569 20947 14603
rect 21925 14569 21959 14603
rect 23765 14569 23799 14603
rect 23857 14569 23891 14603
rect 25421 14569 25455 14603
rect 12541 14501 12575 14535
rect 18052 14501 18086 14535
rect 21281 14501 21315 14535
rect 22753 14501 22787 14535
rect 24961 14501 24995 14535
rect 10793 14433 10827 14467
rect 13093 14433 13127 14467
rect 14013 14433 14047 14467
rect 15669 14433 15703 14467
rect 15761 14433 15795 14467
rect 17785 14433 17819 14467
rect 20729 14433 20763 14467
rect 22477 14433 22511 14467
rect 23213 14433 23247 14467
rect 24225 14433 24259 14467
rect 11069 14365 11103 14399
rect 12633 14365 12667 14399
rect 13553 14365 13587 14399
rect 14197 14365 14231 14399
rect 15853 14365 15887 14399
rect 19993 14365 20027 14399
rect 21373 14365 21407 14399
rect 21557 14365 21591 14399
rect 24317 14365 24351 14399
rect 24501 14365 24535 14399
rect 12081 14297 12115 14331
rect 13645 14297 13679 14331
rect 15117 14297 15151 14331
rect 14657 14229 14691 14263
rect 16313 14229 16347 14263
rect 22293 14229 22327 14263
rect 10609 14025 10643 14059
rect 11621 14025 11655 14059
rect 12173 14025 12207 14059
rect 14933 14025 14967 14059
rect 15485 14025 15519 14059
rect 16405 14025 16439 14059
rect 17509 14025 17543 14059
rect 18337 14025 18371 14059
rect 18889 14025 18923 14059
rect 21649 14025 21683 14059
rect 21833 14025 21867 14059
rect 23121 14025 23155 14059
rect 23857 14025 23891 14059
rect 13369 13957 13403 13991
rect 20361 13957 20395 13991
rect 11069 13889 11103 13923
rect 11161 13889 11195 13923
rect 13553 13889 13587 13923
rect 16221 13889 16255 13923
rect 16865 13889 16899 13923
rect 16957 13889 16991 13923
rect 22385 13889 22419 13923
rect 10149 13821 10183 13855
rect 15853 13821 15887 13855
rect 17785 13821 17819 13855
rect 18981 13821 19015 13855
rect 19237 13821 19271 13855
rect 20913 13821 20947 13855
rect 21373 13821 21407 13855
rect 22293 13821 22327 13855
rect 23489 13821 23523 13855
rect 24133 13821 24167 13855
rect 10517 13753 10551 13787
rect 10977 13753 11011 13787
rect 12541 13753 12575 13787
rect 13820 13753 13854 13787
rect 16773 13753 16807 13787
rect 24400 13753 24434 13787
rect 13093 13685 13127 13719
rect 22201 13685 22235 13719
rect 25513 13685 25547 13719
rect 11713 13481 11747 13515
rect 12357 13481 12391 13515
rect 12725 13481 12759 13515
rect 15025 13481 15059 13515
rect 15301 13481 15335 13515
rect 18245 13481 18279 13515
rect 19165 13481 19199 13515
rect 20913 13481 20947 13515
rect 21557 13481 21591 13515
rect 23489 13481 23523 13515
rect 24593 13481 24627 13515
rect 17110 13413 17144 13447
rect 18797 13413 18831 13447
rect 19625 13413 19659 13447
rect 21925 13413 21959 13447
rect 10589 13345 10623 13379
rect 12817 13345 12851 13379
rect 15669 13345 15703 13379
rect 15761 13345 15795 13379
rect 16865 13345 16899 13379
rect 19349 13345 19383 13379
rect 20085 13345 20119 13379
rect 22376 13345 22410 13379
rect 24961 13345 24995 13379
rect 9689 13277 9723 13311
rect 10333 13277 10367 13311
rect 14565 13277 14599 13311
rect 15853 13277 15887 13311
rect 22109 13277 22143 13311
rect 25053 13277 25087 13311
rect 25145 13277 25179 13311
rect 24225 13209 24259 13243
rect 10149 13141 10183 13175
rect 16405 13141 16439 13175
rect 10609 12937 10643 12971
rect 10793 12937 10827 12971
rect 15117 12937 15151 12971
rect 16037 12937 16071 12971
rect 17417 12937 17451 12971
rect 22017 12937 22051 12971
rect 23489 12937 23523 12971
rect 26341 12937 26375 12971
rect 10333 12869 10367 12903
rect 12173 12869 12207 12903
rect 16405 12869 16439 12903
rect 25697 12869 25731 12903
rect 25973 12869 26007 12903
rect 9781 12801 9815 12835
rect 11253 12801 11287 12835
rect 11437 12801 11471 12835
rect 11805 12801 11839 12835
rect 12725 12801 12759 12835
rect 16957 12801 16991 12835
rect 18337 12801 18371 12835
rect 19993 12801 20027 12835
rect 20453 12801 20487 12835
rect 21005 12801 21039 12835
rect 21557 12801 21591 12835
rect 22569 12801 22603 12835
rect 23029 12801 23063 12835
rect 9413 12733 9447 12767
rect 9505 12733 9539 12767
rect 11161 12733 11195 12767
rect 12449 12733 12483 12767
rect 13737 12733 13771 12767
rect 18061 12733 18095 12767
rect 19257 12733 19291 12767
rect 19901 12733 19935 12767
rect 21925 12733 21959 12767
rect 22477 12733 22511 12767
rect 23673 12733 23707 12767
rect 23929 12733 23963 12767
rect 13645 12665 13679 12699
rect 14004 12665 14038 12699
rect 16865 12665 16899 12699
rect 17785 12665 17819 12699
rect 18981 12665 19015 12699
rect 19809 12665 19843 12699
rect 13185 12597 13219 12631
rect 15669 12597 15703 12631
rect 16773 12597 16807 12631
rect 19441 12597 19475 12631
rect 20913 12597 20947 12631
rect 22385 12597 22419 12631
rect 25053 12597 25087 12631
rect 10333 12393 10367 12427
rect 12633 12393 12667 12427
rect 12817 12393 12851 12427
rect 13645 12393 13679 12427
rect 15301 12393 15335 12427
rect 16497 12393 16531 12427
rect 17233 12393 17267 12427
rect 17969 12393 18003 12427
rect 18245 12393 18279 12427
rect 19257 12393 19291 12427
rect 21189 12393 21223 12427
rect 22109 12393 22143 12427
rect 23581 12393 23615 12427
rect 24685 12393 24719 12427
rect 1654 12325 1688 12359
rect 10946 12325 10980 12359
rect 24501 12325 24535 12359
rect 1409 12257 1443 12291
rect 10057 12257 10091 12291
rect 10701 12257 10735 12291
rect 13185 12257 13219 12291
rect 14013 12257 14047 12291
rect 15669 12257 15703 12291
rect 19165 12257 19199 12291
rect 19625 12257 19659 12291
rect 20729 12257 20763 12291
rect 21741 12257 21775 12291
rect 22201 12257 22235 12291
rect 22468 12257 22502 12291
rect 25053 12257 25087 12291
rect 25145 12257 25179 12291
rect 13277 12189 13311 12223
rect 13369 12189 13403 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 14749 12189 14783 12223
rect 15761 12189 15795 12223
rect 15853 12189 15887 12223
rect 17325 12189 17359 12223
rect 17509 12189 17543 12223
rect 19717 12189 19751 12223
rect 19901 12189 19935 12223
rect 25237 12189 25271 12223
rect 18981 12121 19015 12155
rect 2789 12053 2823 12087
rect 9321 12053 9355 12087
rect 12081 12053 12115 12087
rect 15117 12053 15151 12087
rect 16865 12053 16899 12087
rect 18705 12053 18739 12087
rect 20269 12053 20303 12087
rect 24225 12053 24259 12087
rect 1593 11849 1627 11883
rect 10241 11849 10275 11883
rect 12265 11849 12299 11883
rect 13553 11849 13587 11883
rect 17141 11849 17175 11883
rect 17509 11849 17543 11883
rect 17601 11849 17635 11883
rect 22477 11849 22511 11883
rect 23029 11849 23063 11883
rect 9781 11713 9815 11747
rect 11345 11713 11379 11747
rect 12725 11713 12759 11747
rect 14013 11713 14047 11747
rect 14197 11713 14231 11747
rect 14933 11713 14967 11747
rect 15117 11713 15151 11747
rect 18613 11713 18647 11747
rect 21097 11713 21131 11747
rect 24593 11713 24627 11747
rect 25605 11713 25639 11747
rect 9689 11645 9723 11679
rect 13921 11645 13955 11679
rect 14565 11645 14599 11679
rect 15384 11645 15418 11679
rect 17785 11645 17819 11679
rect 20545 11645 20579 11679
rect 24501 11645 24535 11679
rect 25421 11645 25455 11679
rect 9045 11577 9079 11611
rect 10609 11577 10643 11611
rect 11161 11577 11195 11611
rect 13461 11577 13495 11611
rect 18880 11577 18914 11611
rect 20913 11577 20947 11611
rect 21342 11577 21376 11611
rect 23857 11577 23891 11611
rect 24409 11577 24443 11611
rect 2053 11509 2087 11543
rect 9229 11509 9263 11543
rect 9597 11509 9631 11543
rect 10793 11509 10827 11543
rect 11253 11509 11287 11543
rect 11805 11509 11839 11543
rect 13093 11509 13127 11543
rect 16497 11509 16531 11543
rect 18521 11509 18555 11543
rect 19993 11509 20027 11543
rect 23489 11509 23523 11543
rect 24041 11509 24075 11543
rect 25145 11509 25179 11543
rect 9229 11305 9263 11339
rect 9965 11305 9999 11339
rect 10517 11305 10551 11339
rect 11345 11305 11379 11339
rect 12081 11305 12115 11339
rect 14473 11305 14507 11339
rect 15117 11305 15151 11339
rect 15485 11305 15519 11339
rect 15945 11305 15979 11339
rect 16589 11305 16623 11339
rect 17417 11305 17451 11339
rect 17509 11305 17543 11339
rect 18613 11305 18647 11339
rect 19625 11305 19659 11339
rect 19993 11305 20027 11339
rect 20913 11305 20947 11339
rect 22109 11305 22143 11339
rect 23213 11305 23247 11339
rect 24777 11305 24811 11339
rect 25421 11305 25455 11339
rect 12357 11237 12391 11271
rect 18153 11237 18187 11271
rect 22477 11237 22511 11271
rect 12808 11169 12842 11203
rect 15853 11169 15887 11203
rect 18521 11169 18555 11203
rect 18981 11169 19015 11203
rect 20453 11169 20487 11203
rect 24041 11169 24075 11203
rect 25237 11169 25271 11203
rect 11437 11101 11471 11135
rect 11621 11101 11655 11135
rect 12548 11101 12582 11135
rect 16129 11101 16163 11135
rect 17601 11101 17635 11135
rect 19073 11101 19107 11135
rect 19165 11101 19199 11135
rect 22569 11101 22603 11135
rect 22661 11101 22695 11135
rect 23581 11101 23615 11135
rect 24133 11101 24167 11135
rect 24225 11101 24259 11135
rect 10977 11033 11011 11067
rect 17049 11033 17083 11067
rect 22017 11033 22051 11067
rect 10793 10965 10827 10999
rect 13921 10965 13955 10999
rect 16957 10965 16991 10999
rect 21465 10965 21499 10999
rect 23673 10965 23707 10999
rect 8953 10761 8987 10795
rect 12449 10761 12483 10795
rect 15853 10761 15887 10795
rect 16405 10761 16439 10795
rect 17877 10761 17911 10795
rect 18337 10761 18371 10795
rect 21373 10761 21407 10795
rect 22385 10761 22419 10795
rect 23121 10761 23155 10795
rect 25789 10761 25823 10795
rect 11529 10693 11563 10727
rect 12265 10693 12299 10727
rect 9321 10625 9355 10659
rect 13001 10625 13035 10659
rect 14381 10625 14415 10659
rect 16957 10625 16991 10659
rect 21925 10625 21959 10659
rect 9505 10557 9539 10591
rect 9761 10557 9795 10591
rect 14473 10557 14507 10591
rect 14740 10557 14774 10591
rect 16773 10557 16807 10591
rect 17417 10557 17451 10591
rect 18889 10557 18923 10591
rect 21281 10557 21315 10591
rect 21741 10557 21775 10591
rect 23864 10557 23898 10591
rect 24124 10557 24158 10591
rect 12817 10489 12851 10523
rect 19134 10489 19168 10523
rect 20821 10489 20855 10523
rect 23489 10489 23523 10523
rect 10885 10421 10919 10455
rect 11805 10421 11839 10455
rect 12909 10421 12943 10455
rect 13461 10421 13495 10455
rect 13829 10421 13863 10455
rect 18705 10421 18739 10455
rect 20269 10421 20303 10455
rect 21833 10421 21867 10455
rect 25237 10421 25271 10455
rect 10701 10217 10735 10251
rect 12173 10217 12207 10251
rect 12817 10217 12851 10251
rect 13277 10217 13311 10251
rect 17141 10217 17175 10251
rect 18613 10217 18647 10251
rect 18981 10217 19015 10251
rect 19717 10217 19751 10251
rect 20361 10217 20395 10251
rect 22477 10217 22511 10251
rect 23581 10217 23615 10251
rect 25145 10217 25179 10251
rect 15117 10149 15151 10183
rect 16129 10149 16163 10183
rect 17693 10149 17727 10183
rect 23489 10149 23523 10183
rect 11060 10081 11094 10115
rect 13645 10081 13679 10115
rect 16037 10081 16071 10115
rect 16681 10081 16715 10115
rect 17601 10081 17635 10115
rect 19625 10081 19659 10115
rect 21281 10081 21315 10115
rect 22109 10081 22143 10115
rect 23949 10081 23983 10115
rect 10793 10013 10827 10047
rect 13737 10013 13771 10047
rect 13829 10013 13863 10047
rect 16221 10013 16255 10047
rect 17785 10013 17819 10047
rect 19901 10013 19935 10047
rect 21373 10013 21407 10047
rect 21465 10013 21499 10047
rect 22569 10013 22603 10047
rect 24041 10013 24075 10047
rect 24133 10013 24167 10047
rect 17233 9945 17267 9979
rect 14473 9877 14507 9911
rect 15485 9877 15519 9911
rect 15669 9877 15703 9911
rect 19257 9877 19291 9911
rect 20913 9877 20947 9911
rect 23029 9877 23063 9911
rect 24593 9877 24627 9911
rect 9965 9673 9999 9707
rect 10241 9673 10275 9707
rect 12817 9673 12851 9707
rect 14381 9673 14415 9707
rect 17325 9673 17359 9707
rect 17601 9673 17635 9707
rect 10793 9605 10827 9639
rect 11805 9605 11839 9639
rect 13921 9605 13955 9639
rect 15853 9605 15887 9639
rect 18981 9605 19015 9639
rect 22017 9605 22051 9639
rect 11345 9537 11379 9571
rect 12173 9537 12207 9571
rect 13277 9537 13311 9571
rect 13461 9537 13495 9571
rect 15025 9537 15059 9571
rect 16405 9537 16439 9571
rect 16497 9537 16531 9571
rect 18429 9537 18463 9571
rect 19349 9537 19383 9571
rect 19441 9537 19475 9571
rect 22569 9537 22603 9571
rect 23765 9537 23799 9571
rect 11253 9469 11287 9503
rect 14289 9469 14323 9503
rect 14749 9469 14783 9503
rect 15393 9469 15427 9503
rect 21925 9469 21959 9503
rect 22385 9469 22419 9503
rect 12725 9401 12759 9435
rect 13185 9401 13219 9435
rect 19708 9401 19742 9435
rect 21373 9401 21407 9435
rect 22477 9401 22511 9435
rect 24010 9401 24044 9435
rect 10609 9333 10643 9367
rect 11161 9333 11195 9367
rect 14841 9333 14875 9367
rect 15945 9333 15979 9367
rect 16313 9333 16347 9367
rect 18337 9333 18371 9367
rect 20821 9333 20855 9367
rect 23029 9333 23063 9367
rect 23489 9333 23523 9367
rect 25145 9333 25179 9367
rect 11161 9129 11195 9163
rect 13369 9129 13403 9163
rect 13645 9129 13679 9163
rect 14105 9129 14139 9163
rect 15301 9129 15335 9163
rect 16037 9129 16071 9163
rect 17693 9129 17727 9163
rect 18797 9129 18831 9163
rect 20361 9129 20395 9163
rect 21465 9129 21499 9163
rect 24133 9129 24167 9163
rect 14381 9061 14415 9095
rect 16580 9061 16614 9095
rect 19165 9061 19199 9095
rect 21097 9061 21131 9095
rect 24961 9061 24995 9095
rect 11345 8993 11379 9027
rect 11601 8993 11635 9027
rect 16313 8993 16347 9027
rect 19625 8993 19659 9027
rect 22100 8993 22134 9027
rect 10793 8925 10827 8959
rect 19717 8925 19751 8959
rect 19901 8925 19935 8959
rect 21833 8925 21867 8959
rect 23857 8925 23891 8959
rect 25053 8925 25087 8959
rect 25145 8925 25179 8959
rect 12725 8789 12759 8823
rect 15025 8789 15059 8823
rect 19257 8789 19291 8823
rect 20637 8789 20671 8823
rect 23213 8789 23247 8823
rect 24593 8789 24627 8823
rect 11437 8585 11471 8619
rect 16221 8585 16255 8619
rect 17601 8585 17635 8619
rect 21833 8585 21867 8619
rect 22385 8585 22419 8619
rect 11713 8517 11747 8551
rect 15117 8517 15151 8551
rect 16129 8517 16163 8551
rect 18889 8517 18923 8551
rect 25053 8517 25087 8551
rect 15669 8449 15703 8483
rect 16681 8449 16715 8483
rect 16773 8449 16807 8483
rect 18797 8449 18831 8483
rect 19441 8449 19475 8483
rect 13737 8381 13771 8415
rect 16589 8381 16623 8415
rect 17233 8381 17267 8415
rect 19257 8381 19291 8415
rect 19993 8381 20027 8415
rect 20453 8381 20487 8415
rect 23121 8381 23155 8415
rect 23673 8381 23707 8415
rect 25973 8381 26007 8415
rect 13645 8313 13679 8347
rect 13982 8313 14016 8347
rect 18429 8313 18463 8347
rect 20361 8313 20395 8347
rect 20720 8313 20754 8347
rect 23489 8313 23523 8347
rect 23940 8313 23974 8347
rect 25697 8313 25731 8347
rect 13277 8245 13311 8279
rect 19349 8245 19383 8279
rect 13737 8041 13771 8075
rect 15301 8041 15335 8075
rect 15669 8041 15703 8075
rect 16681 8041 16715 8075
rect 18337 8041 18371 8075
rect 18981 8041 19015 8075
rect 20913 8041 20947 8075
rect 21281 8041 21315 8075
rect 25237 8041 25271 8075
rect 15761 7973 15795 8007
rect 23213 7973 23247 8007
rect 17224 7905 17258 7939
rect 22845 7905 22879 7939
rect 23305 7905 23339 7939
rect 23572 7905 23606 7939
rect 13829 7837 13863 7871
rect 13921 7837 13955 7871
rect 15945 7837 15979 7871
rect 16957 7837 16991 7871
rect 19441 7837 19475 7871
rect 21373 7837 21407 7871
rect 21557 7837 21591 7871
rect 19349 7769 19383 7803
rect 13369 7701 13403 7735
rect 14381 7701 14415 7735
rect 16405 7701 16439 7735
rect 20729 7701 20763 7735
rect 22017 7701 22051 7735
rect 24685 7701 24719 7735
rect 13093 7497 13127 7531
rect 15577 7497 15611 7531
rect 15945 7497 15979 7531
rect 17141 7497 17175 7531
rect 20085 7497 20119 7531
rect 22017 7497 22051 7531
rect 25421 7497 25455 7531
rect 16037 7429 16071 7463
rect 19533 7429 19567 7463
rect 21649 7429 21683 7463
rect 13461 7361 13495 7395
rect 16497 7361 16531 7395
rect 16589 7361 16623 7395
rect 21097 7361 21131 7395
rect 21281 7361 21315 7395
rect 24317 7361 24351 7395
rect 24501 7361 24535 7395
rect 13553 7293 13587 7327
rect 13820 7293 13854 7327
rect 18153 7293 18187 7327
rect 22201 7293 22235 7327
rect 22753 7293 22787 7327
rect 24041 7293 24075 7327
rect 17877 7225 17911 7259
rect 18420 7225 18454 7259
rect 21005 7225 21039 7259
rect 24133 7225 24167 7259
rect 25237 7293 25271 7327
rect 25789 7293 25823 7327
rect 25053 7225 25087 7259
rect 12541 7157 12575 7191
rect 14933 7157 14967 7191
rect 16405 7157 16439 7191
rect 17417 7157 17451 7191
rect 20453 7157 20487 7191
rect 20637 7157 20671 7191
rect 22385 7157 22419 7191
rect 23305 7157 23339 7191
rect 23673 7157 23707 7191
rect 24501 7157 24535 7191
rect 24777 7157 24811 7191
rect 13185 6953 13219 6987
rect 16221 6953 16255 6987
rect 18613 6953 18647 6987
rect 20729 6953 20763 6987
rect 23673 6953 23707 6987
rect 25145 6953 25179 6987
rect 15485 6885 15519 6919
rect 16497 6885 16531 6919
rect 21281 6885 21315 6919
rect 23581 6885 23615 6919
rect 12072 6817 12106 6851
rect 14197 6817 14231 6851
rect 15117 6817 15151 6851
rect 17049 6817 17083 6851
rect 17693 6817 17727 6851
rect 18705 6817 18739 6851
rect 20361 6817 20395 6851
rect 11805 6749 11839 6783
rect 15669 6749 15703 6783
rect 17141 6749 17175 6783
rect 17233 6749 17267 6783
rect 18797 6749 18831 6783
rect 19809 6749 19843 6783
rect 21373 6749 21407 6783
rect 21557 6749 21591 6783
rect 23765 6749 23799 6783
rect 25237 6749 25271 6783
rect 25421 6749 25455 6783
rect 13829 6681 13863 6715
rect 18245 6681 18279 6715
rect 23213 6681 23247 6715
rect 24225 6681 24259 6715
rect 14933 6613 14967 6647
rect 16681 6613 16715 6647
rect 18153 6613 18187 6647
rect 19349 6613 19383 6647
rect 19625 6613 19659 6647
rect 20913 6613 20947 6647
rect 23029 6613 23063 6647
rect 24777 6613 24811 6647
rect 11897 6409 11931 6443
rect 17509 6409 17543 6443
rect 21925 6409 21959 6443
rect 22661 6409 22695 6443
rect 23121 6409 23155 6443
rect 23673 6409 23707 6443
rect 24869 6409 24903 6443
rect 16313 6341 16347 6375
rect 19165 6341 19199 6375
rect 23489 6341 23523 6375
rect 14841 6273 14875 6307
rect 17049 6273 17083 6307
rect 18705 6273 18739 6307
rect 19441 6273 19475 6307
rect 24225 6273 24259 6307
rect 11529 6205 11563 6239
rect 12725 6205 12759 6239
rect 15301 6205 15335 6239
rect 16773 6205 16807 6239
rect 18521 6205 18555 6239
rect 19809 6205 19843 6239
rect 20545 6205 20579 6239
rect 24133 6205 24167 6239
rect 25237 6205 25271 6239
rect 25973 6205 26007 6239
rect 12265 6137 12299 6171
rect 12992 6137 13026 6171
rect 15209 6137 15243 6171
rect 18429 6137 18463 6171
rect 20453 6137 20487 6171
rect 20812 6137 20846 6171
rect 24041 6137 24075 6171
rect 25513 6137 25547 6171
rect 14105 6069 14139 6103
rect 15485 6069 15519 6103
rect 15945 6069 15979 6103
rect 16405 6069 16439 6103
rect 16865 6069 16899 6103
rect 17785 6069 17819 6103
rect 18061 6069 18095 6103
rect 19625 6069 19659 6103
rect 12909 5865 12943 5899
rect 14933 5865 14967 5899
rect 15669 5865 15703 5899
rect 17693 5865 17727 5899
rect 19625 5865 19659 5899
rect 20361 5865 20395 5899
rect 21373 5865 21407 5899
rect 23029 5865 23063 5899
rect 24501 5865 24535 5899
rect 25145 5865 25179 5899
rect 25421 5865 25455 5899
rect 13737 5797 13771 5831
rect 18490 5797 18524 5831
rect 21925 5797 21959 5831
rect 23388 5797 23422 5831
rect 16028 5729 16062 5763
rect 18245 5729 18279 5763
rect 21281 5729 21315 5763
rect 23121 5729 23155 5763
rect 11345 5661 11379 5695
rect 12357 5661 12391 5695
rect 13277 5661 13311 5695
rect 13829 5661 13863 5695
rect 13921 5661 13955 5695
rect 15761 5661 15795 5695
rect 21465 5661 21499 5695
rect 12265 5593 12299 5627
rect 20729 5593 20763 5627
rect 13369 5525 13403 5559
rect 14473 5525 14507 5559
rect 17141 5525 17175 5559
rect 18153 5525 18187 5559
rect 20913 5525 20947 5559
rect 13829 5321 13863 5355
rect 14197 5321 14231 5355
rect 15669 5321 15703 5355
rect 16221 5321 16255 5355
rect 16773 5321 16807 5355
rect 18061 5321 18095 5355
rect 19073 5321 19107 5355
rect 21281 5321 21315 5355
rect 21833 5321 21867 5355
rect 22201 5321 22235 5355
rect 23029 5321 23063 5355
rect 23489 5321 23523 5355
rect 23673 5321 23707 5355
rect 17417 5253 17451 5287
rect 25053 5253 25087 5287
rect 25421 5253 25455 5287
rect 12265 5185 12299 5219
rect 13277 5185 13311 5219
rect 18705 5185 18739 5219
rect 19809 5185 19843 5219
rect 24133 5185 24167 5219
rect 24317 5185 24351 5219
rect 24685 5185 24719 5219
rect 11897 5117 11931 5151
rect 13093 5117 13127 5151
rect 13185 5117 13219 5151
rect 14289 5117 14323 5151
rect 14545 5117 14579 5151
rect 16865 5117 16899 5151
rect 17877 5117 17911 5151
rect 18429 5117 18463 5151
rect 19901 5117 19935 5151
rect 20168 5117 20202 5151
rect 22477 5117 22511 5151
rect 25237 5117 25271 5151
rect 25789 5117 25823 5151
rect 24041 5049 24075 5083
rect 11345 4981 11379 5015
rect 12725 4981 12759 5015
rect 17049 4981 17083 5015
rect 18521 4981 18555 5015
rect 22661 4981 22695 5015
rect 13093 4777 13127 4811
rect 13461 4777 13495 4811
rect 13645 4777 13679 4811
rect 14105 4777 14139 4811
rect 16405 4777 16439 4811
rect 16773 4777 16807 4811
rect 17325 4777 17359 4811
rect 18061 4777 18095 4811
rect 19257 4777 19291 4811
rect 20729 4777 20763 4811
rect 20913 4777 20947 4811
rect 21373 4777 21407 4811
rect 22109 4777 22143 4811
rect 22845 4777 22879 4811
rect 24685 4777 24719 4811
rect 12541 4709 12575 4743
rect 17233 4709 17267 4743
rect 23213 4709 23247 4743
rect 12449 4641 12483 4675
rect 14013 4641 14047 4675
rect 15761 4641 15795 4675
rect 18429 4641 18463 4675
rect 19717 4641 19751 4675
rect 21281 4641 21315 4675
rect 23305 4641 23339 4675
rect 23561 4641 23595 4675
rect 12725 4573 12759 4607
rect 14289 4573 14323 4607
rect 17417 4573 17451 4607
rect 18613 4573 18647 4607
rect 21465 4573 21499 4607
rect 11989 4505 12023 4539
rect 15945 4505 15979 4539
rect 16865 4505 16899 4539
rect 20269 4505 20303 4539
rect 11345 4437 11379 4471
rect 12081 4437 12115 4471
rect 14749 4437 14783 4471
rect 15025 4437 15059 4471
rect 15577 4437 15611 4471
rect 19533 4437 19567 4471
rect 19901 4437 19935 4471
rect 22477 4437 22511 4471
rect 14749 4233 14783 4267
rect 16037 4233 16071 4267
rect 19717 4233 19751 4267
rect 20913 4233 20947 4267
rect 21281 4233 21315 4267
rect 23673 4233 23707 4267
rect 21833 4165 21867 4199
rect 23121 4165 23155 4199
rect 12909 4097 12943 4131
rect 13093 4097 13127 4131
rect 13645 4097 13679 4131
rect 14289 4097 14323 4131
rect 15301 4097 15335 4131
rect 16681 4097 16715 4131
rect 17785 4097 17819 4131
rect 18797 4097 18831 4131
rect 19349 4097 19383 4131
rect 20453 4097 20487 4131
rect 22661 4097 22695 4131
rect 24317 4097 24351 4131
rect 11253 4029 11287 4063
rect 14013 4029 14047 4063
rect 15393 4029 15427 4063
rect 16497 4029 16531 4063
rect 18613 4029 18647 4063
rect 20269 4029 20303 4063
rect 22477 4029 22511 4063
rect 23489 4029 23523 4063
rect 25053 4029 25087 4063
rect 25237 4029 25271 4063
rect 25789 4029 25823 4063
rect 12817 3961 12851 3995
rect 16313 3961 16347 3995
rect 17509 3961 17543 3995
rect 24133 3961 24167 3995
rect 24685 3961 24719 3995
rect 11161 3893 11195 3927
rect 11437 3893 11471 3927
rect 12081 3893 12115 3927
rect 12449 3893 12483 3927
rect 15577 3893 15611 3927
rect 18245 3893 18279 3927
rect 18705 3893 18739 3927
rect 19809 3893 19843 3927
rect 20177 3893 20211 3927
rect 22017 3893 22051 3927
rect 22385 3893 22419 3927
rect 24041 3893 24075 3927
rect 25421 3893 25455 3927
rect 11161 3689 11195 3723
rect 11621 3689 11655 3723
rect 13461 3689 13495 3723
rect 14013 3689 14047 3723
rect 14381 3689 14415 3723
rect 17233 3689 17267 3723
rect 19809 3689 19843 3723
rect 20269 3689 20303 3723
rect 21189 3689 21223 3723
rect 23305 3689 23339 3723
rect 23765 3689 23799 3723
rect 25237 3689 25271 3723
rect 12326 3621 12360 3655
rect 15546 3621 15580 3655
rect 9873 3553 9907 3587
rect 10977 3553 11011 3587
rect 12081 3553 12115 3587
rect 18041 3553 18075 3587
rect 21640 3553 21674 3587
rect 24113 3553 24147 3587
rect 15301 3485 15335 3519
rect 17785 3485 17819 3519
rect 21373 3485 21407 3519
rect 23857 3485 23891 3519
rect 10057 3417 10091 3451
rect 16681 3417 16715 3451
rect 20545 3417 20579 3451
rect 11989 3349 12023 3383
rect 15117 3349 15151 3383
rect 17693 3349 17727 3383
rect 19165 3349 19199 3383
rect 22753 3349 22787 3383
rect 10701 3145 10735 3179
rect 11437 3145 11471 3179
rect 11897 3145 11931 3179
rect 12265 3145 12299 3179
rect 13461 3145 13495 3179
rect 15945 3145 15979 3179
rect 17509 3145 17543 3179
rect 18337 3145 18371 3179
rect 23489 3145 23523 3179
rect 24409 3145 24443 3179
rect 24869 3145 24903 3179
rect 10333 3077 10367 3111
rect 11161 3077 11195 3111
rect 15025 3077 15059 3111
rect 22569 3077 22603 3111
rect 15669 3009 15703 3043
rect 16773 3009 16807 3043
rect 18797 3009 18831 3043
rect 18981 3009 19015 3043
rect 19349 3009 19383 3043
rect 19717 3009 19751 3043
rect 23857 3009 23891 3043
rect 10149 2941 10183 2975
rect 11253 2941 11287 2975
rect 12541 2941 12575 2975
rect 13645 2941 13679 2975
rect 13901 2941 13935 2975
rect 16589 2941 16623 2975
rect 19901 2941 19935 2975
rect 20157 2941 20191 2975
rect 22201 2941 22235 2975
rect 22385 2941 22419 2975
rect 22937 2941 22971 2975
rect 23673 2941 23707 2975
rect 24961 2941 24995 2975
rect 25697 2941 25731 2975
rect 13185 2873 13219 2907
rect 17877 2873 17911 2907
rect 18705 2873 18739 2907
rect 25237 2873 25271 2907
rect 9965 2805 9999 2839
rect 12725 2805 12759 2839
rect 16129 2805 16163 2839
rect 16497 2805 16531 2839
rect 21281 2805 21315 2839
rect 21925 2805 21959 2839
rect 10977 2601 11011 2635
rect 12081 2601 12115 2635
rect 12449 2601 12483 2635
rect 14013 2601 14047 2635
rect 18061 2601 18095 2635
rect 19809 2601 19843 2635
rect 20729 2601 20763 2635
rect 22017 2601 22051 2635
rect 23489 2601 23523 2635
rect 24501 2601 24535 2635
rect 25605 2601 25639 2635
rect 18674 2533 18708 2567
rect 20361 2533 20395 2567
rect 21557 2533 21591 2567
rect 8585 2465 8619 2499
rect 10333 2465 10367 2499
rect 11437 2465 11471 2499
rect 12817 2465 12851 2499
rect 13553 2465 13587 2499
rect 14105 2465 14139 2499
rect 15853 2465 15887 2499
rect 15945 2465 15979 2499
rect 17141 2465 17175 2499
rect 17785 2465 17819 2499
rect 18429 2465 18463 2499
rect 21833 2465 21867 2499
rect 22385 2465 22419 2499
rect 24409 2465 24443 2499
rect 13001 2397 13035 2431
rect 14289 2397 14323 2431
rect 14933 2397 14967 2431
rect 16129 2397 16163 2431
rect 16497 2397 16531 2431
rect 22477 2397 22511 2431
rect 22661 2397 22695 2431
rect 24593 2397 24627 2431
rect 25053 2397 25087 2431
rect 9229 2329 9263 2363
rect 15485 2329 15519 2363
rect 16865 2329 16899 2363
rect 23121 2329 23155 2363
rect 24041 2329 24075 2363
rect 8769 2261 8803 2295
rect 10517 2261 10551 2295
rect 11621 2261 11655 2295
rect 15301 2261 15335 2295
rect 17325 2261 17359 2295
rect 23765 2261 23799 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 16577 25483 16635 25489
rect 16577 25449 16589 25483
rect 16623 25480 16635 25483
rect 17310 25480 17316 25492
rect 16623 25452 17316 25480
rect 16623 25449 16635 25452
rect 16577 25443 16635 25449
rect 17310 25440 17316 25452
rect 17368 25440 17374 25492
rect 20165 25483 20223 25489
rect 20165 25449 20177 25483
rect 20211 25449 20223 25483
rect 20165 25443 20223 25449
rect 21637 25483 21695 25489
rect 21637 25449 21649 25483
rect 21683 25480 21695 25483
rect 22738 25480 22744 25492
rect 21683 25452 22744 25480
rect 21683 25449 21695 25452
rect 21637 25443 21695 25449
rect 20180 25412 20208 25443
rect 22738 25440 22744 25452
rect 22796 25440 22802 25492
rect 22833 25483 22891 25489
rect 22833 25449 22845 25483
rect 22879 25480 22891 25483
rect 24578 25480 24584 25492
rect 22879 25452 24584 25480
rect 22879 25449 22891 25452
rect 22833 25443 22891 25449
rect 24578 25440 24584 25452
rect 24636 25440 24642 25492
rect 24762 25480 24768 25492
rect 24723 25452 24768 25480
rect 24762 25440 24768 25452
rect 24820 25440 24826 25492
rect 24118 25412 24124 25424
rect 20180 25384 24124 25412
rect 24118 25372 24124 25384
rect 24176 25372 24182 25424
rect 16298 25304 16304 25356
rect 16356 25344 16362 25356
rect 16393 25347 16451 25353
rect 16393 25344 16405 25347
rect 16356 25316 16405 25344
rect 16356 25304 16362 25316
rect 16393 25313 16405 25316
rect 16439 25313 16451 25347
rect 16393 25307 16451 25313
rect 18877 25347 18935 25353
rect 18877 25313 18889 25347
rect 18923 25344 18935 25347
rect 18966 25344 18972 25356
rect 18923 25316 18972 25344
rect 18923 25313 18935 25316
rect 18877 25307 18935 25313
rect 18966 25304 18972 25316
rect 19024 25304 19030 25356
rect 19981 25347 20039 25353
rect 19981 25313 19993 25347
rect 20027 25344 20039 25347
rect 20162 25344 20168 25356
rect 20027 25316 20168 25344
rect 20027 25313 20039 25316
rect 19981 25307 20039 25313
rect 20162 25304 20168 25316
rect 20220 25304 20226 25356
rect 21453 25347 21511 25353
rect 21453 25313 21465 25347
rect 21499 25344 21511 25347
rect 22370 25344 22376 25356
rect 21499 25316 22376 25344
rect 21499 25313 21511 25316
rect 21453 25307 21511 25313
rect 22370 25304 22376 25316
rect 22428 25304 22434 25356
rect 22554 25304 22560 25356
rect 22612 25344 22618 25356
rect 22649 25347 22707 25353
rect 22649 25344 22661 25347
rect 22612 25316 22661 25344
rect 22612 25304 22618 25316
rect 22649 25313 22661 25316
rect 22695 25313 22707 25347
rect 22649 25307 22707 25313
rect 23934 25304 23940 25356
rect 23992 25344 23998 25356
rect 24581 25347 24639 25353
rect 24581 25344 24593 25347
rect 23992 25316 24593 25344
rect 23992 25304 23998 25316
rect 24581 25313 24593 25316
rect 24627 25313 24639 25347
rect 24581 25307 24639 25313
rect 19061 25211 19119 25217
rect 19061 25177 19073 25211
rect 19107 25208 19119 25211
rect 26878 25208 26884 25220
rect 19107 25180 26884 25208
rect 19107 25177 19119 25180
rect 19061 25171 19119 25177
rect 26878 25168 26884 25180
rect 26936 25168 26942 25220
rect 19426 25140 19432 25152
rect 19387 25112 19432 25140
rect 19426 25100 19432 25112
rect 19484 25100 19490 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 17037 24939 17095 24945
rect 17037 24905 17049 24939
rect 17083 24936 17095 24939
rect 24762 24936 24768 24948
rect 17083 24908 24768 24936
rect 17083 24905 17095 24908
rect 17037 24899 17095 24905
rect 24762 24896 24768 24908
rect 24820 24896 24826 24948
rect 22554 24828 22560 24880
rect 22612 24868 22618 24880
rect 23385 24871 23443 24877
rect 23385 24868 23397 24871
rect 22612 24840 23397 24868
rect 22612 24828 22618 24840
rect 23385 24837 23397 24840
rect 23431 24837 23443 24871
rect 23385 24831 23443 24837
rect 15933 24803 15991 24809
rect 15933 24800 15945 24803
rect 15304 24772 15945 24800
rect 15304 24741 15332 24772
rect 15933 24769 15945 24772
rect 15979 24800 15991 24803
rect 17034 24800 17040 24812
rect 15979 24772 17040 24800
rect 15979 24769 15991 24772
rect 15933 24763 15991 24769
rect 17034 24760 17040 24772
rect 17092 24760 17098 24812
rect 14185 24735 14243 24741
rect 14185 24701 14197 24735
rect 14231 24732 14243 24735
rect 15289 24735 15347 24741
rect 14231 24704 14596 24732
rect 14231 24701 14243 24704
rect 14185 24695 14243 24701
rect 14568 24608 14596 24704
rect 15289 24701 15301 24735
rect 15335 24701 15347 24735
rect 16850 24732 16856 24744
rect 16763 24704 16856 24732
rect 15289 24695 15347 24701
rect 16850 24692 16856 24704
rect 16908 24732 16914 24744
rect 17405 24735 17463 24741
rect 17405 24732 17417 24735
rect 16908 24704 17417 24732
rect 16908 24692 16914 24704
rect 17405 24701 17417 24704
rect 17451 24701 17463 24735
rect 18049 24735 18107 24741
rect 18049 24732 18061 24735
rect 17405 24695 17463 24701
rect 17788 24704 18061 24732
rect 16482 24664 16488 24676
rect 15488 24636 16488 24664
rect 14366 24596 14372 24608
rect 14327 24568 14372 24596
rect 14366 24556 14372 24568
rect 14424 24556 14430 24608
rect 14550 24556 14556 24608
rect 14608 24596 14614 24608
rect 15488 24605 15516 24636
rect 16482 24624 16488 24636
rect 16540 24624 16546 24676
rect 17788 24608 17816 24704
rect 18049 24701 18061 24704
rect 18095 24701 18107 24735
rect 18049 24695 18107 24701
rect 19153 24735 19211 24741
rect 19153 24701 19165 24735
rect 19199 24732 19211 24735
rect 19242 24732 19248 24744
rect 19199 24704 19248 24732
rect 19199 24701 19211 24704
rect 19153 24695 19211 24701
rect 19242 24692 19248 24704
rect 19300 24692 19306 24744
rect 20254 24732 20260 24744
rect 20215 24704 20260 24732
rect 20254 24692 20260 24704
rect 20312 24732 20318 24744
rect 20809 24735 20867 24741
rect 20809 24732 20821 24735
rect 20312 24704 20821 24732
rect 20312 24692 20318 24704
rect 20809 24701 20821 24704
rect 20855 24701 20867 24735
rect 20809 24695 20867 24701
rect 21361 24735 21419 24741
rect 21361 24701 21373 24735
rect 21407 24732 21419 24735
rect 21910 24732 21916 24744
rect 21407 24704 21916 24732
rect 21407 24701 21419 24704
rect 21361 24695 21419 24701
rect 21910 24692 21916 24704
rect 21968 24692 21974 24744
rect 22462 24732 22468 24744
rect 22423 24704 22468 24732
rect 22462 24692 22468 24704
rect 22520 24732 22526 24744
rect 23017 24735 23075 24741
rect 23017 24732 23029 24735
rect 22520 24704 23029 24732
rect 22520 24692 22526 24704
rect 23017 24701 23029 24704
rect 23063 24701 23075 24735
rect 23017 24695 23075 24701
rect 23842 24692 23848 24744
rect 23900 24732 23906 24744
rect 24581 24735 24639 24741
rect 24581 24732 24593 24735
rect 23900 24704 24593 24732
rect 23900 24692 23906 24704
rect 24581 24701 24593 24704
rect 24627 24732 24639 24735
rect 25133 24735 25191 24741
rect 25133 24732 25145 24735
rect 24627 24704 25145 24732
rect 24627 24701 24639 24704
rect 24581 24695 24639 24701
rect 25133 24701 25145 24704
rect 25179 24701 25191 24735
rect 25133 24695 25191 24701
rect 20070 24664 20076 24676
rect 19352 24636 20076 24664
rect 14737 24599 14795 24605
rect 14737 24596 14749 24599
rect 14608 24568 14749 24596
rect 14608 24556 14614 24568
rect 14737 24565 14749 24568
rect 14783 24565 14795 24599
rect 14737 24559 14795 24565
rect 15473 24599 15531 24605
rect 15473 24565 15485 24599
rect 15519 24565 15531 24599
rect 15473 24559 15531 24565
rect 16298 24556 16304 24608
rect 16356 24596 16362 24608
rect 16393 24599 16451 24605
rect 16393 24596 16405 24599
rect 16356 24568 16405 24596
rect 16356 24556 16362 24568
rect 16393 24565 16405 24568
rect 16439 24565 16451 24599
rect 17770 24596 17776 24608
rect 17731 24568 17776 24596
rect 16393 24559 16451 24565
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 17954 24556 17960 24608
rect 18012 24596 18018 24608
rect 18233 24599 18291 24605
rect 18233 24596 18245 24599
rect 18012 24568 18245 24596
rect 18012 24556 18018 24568
rect 18233 24565 18245 24568
rect 18279 24565 18291 24599
rect 18966 24596 18972 24608
rect 18927 24568 18972 24596
rect 18233 24559 18291 24565
rect 18966 24556 18972 24568
rect 19024 24556 19030 24608
rect 19352 24605 19380 24636
rect 20070 24624 20076 24636
rect 20128 24624 20134 24676
rect 22002 24664 22008 24676
rect 21560 24636 22008 24664
rect 19337 24599 19395 24605
rect 19337 24565 19349 24599
rect 19383 24565 19395 24599
rect 19337 24559 19395 24565
rect 19981 24599 20039 24605
rect 19981 24565 19993 24599
rect 20027 24596 20039 24599
rect 20162 24596 20168 24608
rect 20027 24568 20168 24596
rect 20027 24565 20039 24568
rect 19981 24559 20039 24565
rect 20162 24556 20168 24568
rect 20220 24556 20226 24608
rect 20441 24599 20499 24605
rect 20441 24565 20453 24599
rect 20487 24596 20499 24599
rect 20622 24596 20628 24608
rect 20487 24568 20628 24596
rect 20487 24565 20499 24568
rect 20441 24559 20499 24565
rect 20622 24556 20628 24568
rect 20680 24556 20686 24608
rect 21560 24605 21588 24636
rect 22002 24624 22008 24636
rect 22060 24624 22066 24676
rect 21545 24599 21603 24605
rect 21545 24565 21557 24599
rect 21591 24565 21603 24599
rect 21910 24596 21916 24608
rect 21871 24568 21916 24596
rect 21545 24559 21603 24565
rect 21910 24556 21916 24568
rect 21968 24556 21974 24608
rect 22370 24596 22376 24608
rect 22331 24568 22376 24596
rect 22370 24556 22376 24568
rect 22428 24556 22434 24608
rect 22649 24599 22707 24605
rect 22649 24565 22661 24599
rect 22695 24596 22707 24599
rect 23290 24596 23296 24608
rect 22695 24568 23296 24596
rect 22695 24565 22707 24568
rect 22649 24559 22707 24565
rect 23290 24556 23296 24568
rect 23348 24556 23354 24608
rect 23934 24556 23940 24608
rect 23992 24596 23998 24608
rect 24397 24599 24455 24605
rect 24397 24596 24409 24599
rect 23992 24568 24409 24596
rect 23992 24556 23998 24568
rect 24397 24565 24409 24568
rect 24443 24565 24455 24599
rect 24762 24596 24768 24608
rect 24723 24568 24768 24596
rect 24397 24559 24455 24565
rect 24762 24556 24768 24568
rect 24820 24556 24826 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 13081 24395 13139 24401
rect 13081 24361 13093 24395
rect 13127 24392 13139 24395
rect 13722 24392 13728 24404
rect 13127 24364 13728 24392
rect 13127 24361 13139 24364
rect 13081 24355 13139 24361
rect 13722 24352 13728 24364
rect 13780 24352 13786 24404
rect 14277 24395 14335 24401
rect 14277 24361 14289 24395
rect 14323 24392 14335 24395
rect 15102 24392 15108 24404
rect 14323 24364 15108 24392
rect 14323 24361 14335 24364
rect 14277 24355 14335 24361
rect 15102 24352 15108 24364
rect 15160 24352 15166 24404
rect 17954 24392 17960 24404
rect 17915 24364 17960 24392
rect 17954 24352 17960 24364
rect 18012 24352 18018 24404
rect 18690 24352 18696 24404
rect 18748 24392 18754 24404
rect 19337 24395 19395 24401
rect 19337 24392 19349 24395
rect 18748 24364 19349 24392
rect 18748 24352 18754 24364
rect 19337 24361 19349 24364
rect 19383 24361 19395 24395
rect 19337 24355 19395 24361
rect 21085 24395 21143 24401
rect 21085 24361 21097 24395
rect 21131 24392 21143 24395
rect 21358 24392 21364 24404
rect 21131 24364 21364 24392
rect 21131 24361 21143 24364
rect 21085 24355 21143 24361
rect 21358 24352 21364 24364
rect 21416 24352 21422 24404
rect 22557 24395 22615 24401
rect 22557 24361 22569 24395
rect 22603 24392 22615 24395
rect 23106 24392 23112 24404
rect 22603 24364 23112 24392
rect 22603 24361 22615 24364
rect 22557 24355 22615 24361
rect 23106 24352 23112 24364
rect 23164 24352 23170 24404
rect 23658 24392 23664 24404
rect 23619 24364 23664 24392
rect 23658 24352 23664 24364
rect 23716 24352 23722 24404
rect 13906 24284 13912 24336
rect 13964 24324 13970 24336
rect 15657 24327 15715 24333
rect 15657 24324 15669 24327
rect 13964 24296 15669 24324
rect 13964 24284 13970 24296
rect 15657 24293 15669 24296
rect 15703 24324 15715 24327
rect 16390 24324 16396 24336
rect 15703 24296 16396 24324
rect 15703 24293 15715 24296
rect 15657 24287 15715 24293
rect 16390 24284 16396 24296
rect 16448 24284 16454 24336
rect 20070 24324 20076 24336
rect 18708 24296 20076 24324
rect 14090 24256 14096 24268
rect 14051 24228 14096 24256
rect 14090 24216 14096 24228
rect 14148 24216 14154 24268
rect 14182 24216 14188 24268
rect 14240 24256 14246 24268
rect 15746 24256 15752 24268
rect 14240 24228 15752 24256
rect 14240 24216 14246 24228
rect 15746 24216 15752 24228
rect 15804 24216 15810 24268
rect 17678 24216 17684 24268
rect 17736 24256 17742 24268
rect 18049 24259 18107 24265
rect 18049 24256 18061 24259
rect 17736 24228 18061 24256
rect 17736 24216 17742 24228
rect 18049 24225 18061 24228
rect 18095 24256 18107 24259
rect 18708 24256 18736 24296
rect 20070 24284 20076 24296
rect 20128 24284 20134 24336
rect 19150 24256 19156 24268
rect 18095 24228 18736 24256
rect 19111 24228 19156 24256
rect 18095 24225 18107 24228
rect 18049 24219 18107 24225
rect 19150 24216 19156 24228
rect 19208 24216 19214 24268
rect 20901 24259 20959 24265
rect 20901 24225 20913 24259
rect 20947 24256 20959 24259
rect 21726 24256 21732 24268
rect 20947 24228 21732 24256
rect 20947 24225 20959 24228
rect 20901 24219 20959 24225
rect 21726 24216 21732 24228
rect 21784 24216 21790 24268
rect 22373 24259 22431 24265
rect 22373 24225 22385 24259
rect 22419 24256 22431 24259
rect 23014 24256 23020 24268
rect 22419 24228 23020 24256
rect 22419 24225 22431 24228
rect 22373 24219 22431 24225
rect 23014 24216 23020 24228
rect 23072 24216 23078 24268
rect 23474 24256 23480 24268
rect 23435 24228 23480 24256
rect 23474 24216 23480 24228
rect 23532 24216 23538 24268
rect 24026 24216 24032 24268
rect 24084 24256 24090 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 24084 24228 24593 24256
rect 24084 24216 24090 24228
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24188 15991 24191
rect 16022 24188 16028 24200
rect 15979 24160 16028 24188
rect 15979 24157 15991 24160
rect 15933 24151 15991 24157
rect 16022 24148 16028 24160
rect 16080 24148 16086 24200
rect 18141 24191 18199 24197
rect 18141 24157 18153 24191
rect 18187 24157 18199 24191
rect 18141 24151 18199 24157
rect 18156 24120 18184 24151
rect 18322 24120 18328 24132
rect 17420 24092 18328 24120
rect 17420 24064 17448 24092
rect 18322 24080 18328 24092
rect 18380 24120 18386 24132
rect 18601 24123 18659 24129
rect 18601 24120 18613 24123
rect 18380 24092 18613 24120
rect 18380 24080 18386 24092
rect 18601 24089 18613 24092
rect 18647 24089 18659 24123
rect 18601 24083 18659 24089
rect 15289 24055 15347 24061
rect 15289 24021 15301 24055
rect 15335 24052 15347 24055
rect 16482 24052 16488 24064
rect 15335 24024 16488 24052
rect 15335 24021 15347 24024
rect 15289 24015 15347 24021
rect 16482 24012 16488 24024
rect 16540 24012 16546 24064
rect 16666 24052 16672 24064
rect 16627 24024 16672 24052
rect 16666 24012 16672 24024
rect 16724 24012 16730 24064
rect 17402 24052 17408 24064
rect 17363 24024 17408 24052
rect 17402 24012 17408 24024
rect 17460 24012 17466 24064
rect 17586 24052 17592 24064
rect 17547 24024 17592 24052
rect 17586 24012 17592 24024
rect 17644 24012 17650 24064
rect 24670 24012 24676 24064
rect 24728 24052 24734 24064
rect 24765 24055 24823 24061
rect 24765 24052 24777 24055
rect 24728 24024 24777 24052
rect 24728 24012 24734 24024
rect 24765 24021 24777 24024
rect 24811 24021 24823 24055
rect 24765 24015 24823 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 12802 23848 12808 23860
rect 12763 23820 12808 23848
rect 12802 23808 12808 23820
rect 12860 23808 12866 23860
rect 15746 23808 15752 23860
rect 15804 23848 15810 23860
rect 16025 23851 16083 23857
rect 16025 23848 16037 23851
rect 15804 23820 16037 23848
rect 15804 23808 15810 23820
rect 16025 23817 16037 23820
rect 16071 23817 16083 23851
rect 16390 23848 16396 23860
rect 16351 23820 16396 23848
rect 16025 23811 16083 23817
rect 16390 23808 16396 23820
rect 16448 23808 16454 23860
rect 17126 23808 17132 23860
rect 17184 23848 17190 23860
rect 17678 23848 17684 23860
rect 17184 23820 17684 23848
rect 17184 23808 17190 23820
rect 17678 23808 17684 23820
rect 17736 23808 17742 23860
rect 19518 23808 19524 23860
rect 19576 23848 19582 23860
rect 20717 23851 20775 23857
rect 20717 23848 20729 23851
rect 19576 23820 20729 23848
rect 19576 23808 19582 23820
rect 20717 23817 20729 23820
rect 20763 23817 20775 23851
rect 20717 23811 20775 23817
rect 22649 23851 22707 23857
rect 22649 23817 22661 23851
rect 22695 23848 22707 23851
rect 23198 23848 23204 23860
rect 22695 23820 23204 23848
rect 22695 23817 22707 23820
rect 22649 23811 22707 23817
rect 23198 23808 23204 23820
rect 23256 23808 23262 23860
rect 16850 23712 16856 23724
rect 16811 23684 16856 23712
rect 16850 23672 16856 23684
rect 16908 23672 16914 23724
rect 12621 23647 12679 23653
rect 12621 23613 12633 23647
rect 12667 23644 12679 23647
rect 14093 23647 14151 23653
rect 14093 23644 14105 23647
rect 12667 23616 13308 23644
rect 12667 23613 12679 23616
rect 12621 23607 12679 23613
rect 13280 23585 13308 23616
rect 13556 23616 14105 23644
rect 13265 23579 13323 23585
rect 13265 23545 13277 23579
rect 13311 23576 13323 23579
rect 13446 23576 13452 23588
rect 13311 23548 13452 23576
rect 13311 23545 13323 23548
rect 13265 23539 13323 23545
rect 13446 23536 13452 23548
rect 13504 23536 13510 23588
rect 13556 23520 13584 23616
rect 14093 23613 14105 23616
rect 14139 23613 14151 23647
rect 14093 23607 14151 23613
rect 16577 23647 16635 23653
rect 16577 23613 16589 23647
rect 16623 23644 16635 23647
rect 16666 23644 16672 23656
rect 16623 23616 16672 23644
rect 16623 23613 16635 23616
rect 16577 23607 16635 23613
rect 16666 23604 16672 23616
rect 16724 23644 16730 23656
rect 17494 23644 17500 23656
rect 16724 23616 17500 23644
rect 16724 23604 16730 23616
rect 17494 23604 17500 23616
rect 17552 23604 17558 23656
rect 18046 23644 18052 23656
rect 18007 23616 18052 23644
rect 18046 23604 18052 23616
rect 18104 23604 18110 23656
rect 18322 23653 18328 23656
rect 18316 23644 18328 23653
rect 18283 23616 18328 23644
rect 18316 23607 18328 23616
rect 18322 23604 18328 23607
rect 18380 23604 18386 23656
rect 20070 23604 20076 23656
rect 20128 23644 20134 23656
rect 20533 23647 20591 23653
rect 20533 23644 20545 23647
rect 20128 23616 20545 23644
rect 20128 23604 20134 23616
rect 20533 23613 20545 23616
rect 20579 23644 20591 23647
rect 21085 23647 21143 23653
rect 21085 23644 21097 23647
rect 20579 23616 21097 23644
rect 20579 23613 20591 23616
rect 20533 23607 20591 23613
rect 21085 23613 21097 23616
rect 21131 23613 21143 23647
rect 21085 23607 21143 23613
rect 22465 23647 22523 23653
rect 22465 23613 22477 23647
rect 22511 23644 22523 23647
rect 22511 23616 22545 23644
rect 22511 23613 22523 23616
rect 22465 23607 22523 23613
rect 14338 23579 14396 23585
rect 14338 23576 14350 23579
rect 14016 23548 14350 23576
rect 14016 23520 14044 23548
rect 14338 23545 14350 23548
rect 14384 23545 14396 23579
rect 14338 23539 14396 23545
rect 19150 23536 19156 23588
rect 19208 23576 19214 23588
rect 19981 23579 20039 23585
rect 19981 23576 19993 23579
rect 19208 23548 19993 23576
rect 19208 23536 19214 23548
rect 19981 23545 19993 23548
rect 20027 23545 20039 23579
rect 19981 23539 20039 23545
rect 22373 23579 22431 23585
rect 22373 23545 22385 23579
rect 22419 23576 22431 23579
rect 22480 23576 22508 23607
rect 24210 23604 24216 23656
rect 24268 23644 24274 23656
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 24268 23616 24593 23644
rect 24268 23604 24274 23616
rect 24581 23613 24593 23616
rect 24627 23644 24639 23647
rect 25133 23647 25191 23653
rect 25133 23644 25145 23647
rect 24627 23616 25145 23644
rect 24627 23613 24639 23616
rect 24581 23607 24639 23613
rect 25133 23613 25145 23616
rect 25179 23613 25191 23647
rect 25133 23607 25191 23613
rect 23566 23576 23572 23588
rect 22419 23548 23572 23576
rect 22419 23545 22431 23548
rect 22373 23539 22431 23545
rect 23566 23536 23572 23548
rect 23624 23536 23630 23588
rect 13538 23508 13544 23520
rect 13499 23480 13544 23508
rect 13538 23468 13544 23480
rect 13596 23468 13602 23520
rect 13998 23508 14004 23520
rect 13959 23480 14004 23508
rect 13998 23468 14004 23480
rect 14056 23468 14062 23520
rect 15378 23468 15384 23520
rect 15436 23508 15442 23520
rect 15473 23511 15531 23517
rect 15473 23508 15485 23511
rect 15436 23480 15485 23508
rect 15436 23468 15442 23480
rect 15473 23477 15485 23480
rect 15519 23477 15531 23511
rect 15473 23471 15531 23477
rect 19334 23468 19340 23520
rect 19392 23508 19398 23520
rect 19429 23511 19487 23517
rect 19429 23508 19441 23511
rect 19392 23480 19441 23508
rect 19392 23468 19398 23480
rect 19429 23477 19441 23480
rect 19475 23477 19487 23511
rect 19429 23471 19487 23477
rect 21545 23511 21603 23517
rect 21545 23477 21557 23511
rect 21591 23508 21603 23511
rect 21726 23508 21732 23520
rect 21591 23480 21732 23508
rect 21591 23477 21603 23480
rect 21545 23471 21603 23477
rect 21726 23468 21732 23480
rect 21784 23468 21790 23520
rect 23014 23508 23020 23520
rect 22975 23480 23020 23508
rect 23014 23468 23020 23480
rect 23072 23468 23078 23520
rect 23474 23468 23480 23520
rect 23532 23508 23538 23520
rect 23845 23511 23903 23517
rect 23845 23508 23857 23511
rect 23532 23480 23857 23508
rect 23532 23468 23538 23480
rect 23845 23477 23857 23480
rect 23891 23477 23903 23511
rect 23845 23471 23903 23477
rect 24026 23468 24032 23520
rect 24084 23508 24090 23520
rect 24397 23511 24455 23517
rect 24397 23508 24409 23511
rect 24084 23480 24409 23508
rect 24084 23468 24090 23480
rect 24397 23477 24409 23480
rect 24443 23477 24455 23511
rect 24762 23508 24768 23520
rect 24723 23480 24768 23508
rect 24397 23471 24455 23477
rect 24762 23468 24768 23480
rect 24820 23468 24826 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 12437 23307 12495 23313
rect 12437 23273 12449 23307
rect 12483 23304 12495 23307
rect 12618 23304 12624 23316
rect 12483 23276 12624 23304
rect 12483 23273 12495 23276
rect 12437 23267 12495 23273
rect 12618 23264 12624 23276
rect 12676 23304 12682 23316
rect 13538 23304 13544 23316
rect 12676 23276 13544 23304
rect 12676 23264 12682 23276
rect 13538 23264 13544 23276
rect 13596 23304 13602 23316
rect 14642 23304 14648 23316
rect 13596 23276 14648 23304
rect 13596 23264 13602 23276
rect 14642 23264 14648 23276
rect 14700 23264 14706 23316
rect 17681 23307 17739 23313
rect 17681 23273 17693 23307
rect 17727 23304 17739 23307
rect 17862 23304 17868 23316
rect 17727 23276 17868 23304
rect 17727 23273 17739 23276
rect 17681 23267 17739 23273
rect 17862 23264 17868 23276
rect 17920 23264 17926 23316
rect 18046 23264 18052 23316
rect 18104 23304 18110 23316
rect 18969 23307 19027 23313
rect 18969 23304 18981 23307
rect 18104 23276 18981 23304
rect 18104 23264 18110 23276
rect 18969 23273 18981 23276
rect 19015 23304 19027 23307
rect 19058 23304 19064 23316
rect 19015 23276 19064 23304
rect 19015 23273 19027 23276
rect 18969 23267 19027 23273
rect 19058 23264 19064 23276
rect 19116 23264 19122 23316
rect 17586 23196 17592 23248
rect 17644 23236 17650 23248
rect 18325 23239 18383 23245
rect 18325 23236 18337 23239
rect 17644 23208 18337 23236
rect 17644 23196 17650 23208
rect 18325 23205 18337 23208
rect 18371 23205 18383 23239
rect 18325 23199 18383 23205
rect 22741 23239 22799 23245
rect 22741 23205 22753 23239
rect 22787 23236 22799 23239
rect 23474 23236 23480 23248
rect 22787 23208 23480 23236
rect 22787 23205 22799 23208
rect 22741 23199 22799 23205
rect 23474 23196 23480 23208
rect 23532 23196 23538 23248
rect 23566 23196 23572 23248
rect 23624 23236 23630 23248
rect 24029 23239 24087 23245
rect 24029 23236 24041 23239
rect 23624 23208 24041 23236
rect 23624 23196 23630 23208
rect 24029 23205 24041 23208
rect 24075 23205 24087 23239
rect 24029 23199 24087 23205
rect 10686 23177 10692 23180
rect 10680 23131 10692 23177
rect 10744 23168 10750 23180
rect 13262 23168 13268 23180
rect 10744 23140 10780 23168
rect 13223 23140 13268 23168
rect 10686 23128 10692 23131
rect 10744 23128 10750 23140
rect 13262 23128 13268 23140
rect 13320 23128 13326 23180
rect 15105 23171 15163 23177
rect 15105 23137 15117 23171
rect 15151 23168 15163 23171
rect 15378 23168 15384 23180
rect 15151 23140 15384 23168
rect 15151 23137 15163 23140
rect 15105 23131 15163 23137
rect 15378 23128 15384 23140
rect 15436 23168 15442 23180
rect 15740 23171 15798 23177
rect 15740 23168 15752 23171
rect 15436 23140 15752 23168
rect 15436 23128 15442 23140
rect 15740 23137 15752 23140
rect 15786 23168 15798 23171
rect 16022 23168 16028 23180
rect 15786 23140 16028 23168
rect 15786 23137 15798 23140
rect 15740 23131 15798 23137
rect 16022 23128 16028 23140
rect 16080 23128 16086 23180
rect 19521 23171 19579 23177
rect 19521 23168 19533 23171
rect 17972 23140 19533 23168
rect 10413 23103 10471 23109
rect 10413 23100 10425 23103
rect 10244 23072 10425 23100
rect 10042 22924 10048 22976
rect 10100 22964 10106 22976
rect 10244 22973 10272 23072
rect 10413 23069 10425 23072
rect 10459 23069 10471 23103
rect 13357 23103 13415 23109
rect 13357 23100 13369 23103
rect 10413 23063 10471 23069
rect 12728 23072 13369 23100
rect 12728 22976 12756 23072
rect 13357 23069 13369 23072
rect 13403 23069 13415 23103
rect 13538 23100 13544 23112
rect 13499 23072 13544 23100
rect 13357 23063 13415 23069
rect 13538 23060 13544 23072
rect 13596 23060 13602 23112
rect 14642 23060 14648 23112
rect 14700 23100 14706 23112
rect 15473 23103 15531 23109
rect 15473 23100 15485 23103
rect 14700 23072 15485 23100
rect 14700 23060 14706 23072
rect 15473 23069 15485 23072
rect 15519 23069 15531 23103
rect 15473 23063 15531 23069
rect 17972 23041 18000 23140
rect 19521 23137 19533 23140
rect 19567 23168 19579 23171
rect 20254 23168 20260 23180
rect 19567 23140 20260 23168
rect 19567 23137 19579 23140
rect 19521 23131 19579 23137
rect 20254 23128 20260 23140
rect 20312 23128 20318 23180
rect 20806 23128 20812 23180
rect 20864 23168 20870 23180
rect 21269 23171 21327 23177
rect 21269 23168 21281 23171
rect 20864 23140 21281 23168
rect 20864 23128 20870 23140
rect 21269 23137 21281 23140
rect 21315 23137 21327 23171
rect 21269 23131 21327 23137
rect 22465 23171 22523 23177
rect 22465 23137 22477 23171
rect 22511 23168 22523 23171
rect 22922 23168 22928 23180
rect 22511 23140 22928 23168
rect 22511 23137 22523 23140
rect 22465 23131 22523 23137
rect 22922 23128 22928 23140
rect 22980 23128 22986 23180
rect 23750 23168 23756 23180
rect 23711 23140 23756 23168
rect 23750 23128 23756 23140
rect 23808 23128 23814 23180
rect 25038 23168 25044 23180
rect 24999 23140 25044 23168
rect 25038 23128 25044 23140
rect 25096 23128 25102 23180
rect 18414 23100 18420 23112
rect 18375 23072 18420 23100
rect 18414 23060 18420 23072
rect 18472 23060 18478 23112
rect 18601 23103 18659 23109
rect 18601 23069 18613 23103
rect 18647 23100 18659 23103
rect 19334 23100 19340 23112
rect 18647 23072 19340 23100
rect 18647 23069 18659 23072
rect 18601 23063 18659 23069
rect 19334 23060 19340 23072
rect 19392 23060 19398 23112
rect 19794 23100 19800 23112
rect 19755 23072 19800 23100
rect 19794 23060 19800 23072
rect 19852 23060 19858 23112
rect 20990 23060 20996 23112
rect 21048 23100 21054 23112
rect 21361 23103 21419 23109
rect 21361 23100 21373 23103
rect 21048 23072 21373 23100
rect 21048 23060 21054 23072
rect 21361 23069 21373 23072
rect 21407 23069 21419 23103
rect 21361 23063 21419 23069
rect 21450 23060 21456 23112
rect 21508 23100 21514 23112
rect 22094 23100 22100 23112
rect 21508 23072 22100 23100
rect 21508 23060 21514 23072
rect 22094 23060 22100 23072
rect 22152 23100 22158 23112
rect 22281 23103 22339 23109
rect 22281 23100 22293 23103
rect 22152 23072 22293 23100
rect 22152 23060 22158 23072
rect 22281 23069 22293 23072
rect 22327 23069 22339 23103
rect 22281 23063 22339 23069
rect 17957 23035 18015 23041
rect 17957 23001 17969 23035
rect 18003 23001 18015 23035
rect 17957 22995 18015 23001
rect 10229 22967 10287 22973
rect 10229 22964 10241 22967
rect 10100 22936 10241 22964
rect 10100 22924 10106 22936
rect 10229 22933 10241 22936
rect 10275 22933 10287 22967
rect 11790 22964 11796 22976
rect 11751 22936 11796 22964
rect 10229 22927 10287 22933
rect 11790 22924 11796 22936
rect 11848 22924 11854 22976
rect 12710 22964 12716 22976
rect 12671 22936 12716 22964
rect 12710 22924 12716 22936
rect 12768 22924 12774 22976
rect 12894 22964 12900 22976
rect 12855 22936 12900 22964
rect 12894 22924 12900 22936
rect 12952 22924 12958 22976
rect 14090 22964 14096 22976
rect 14051 22936 14096 22964
rect 14090 22924 14096 22936
rect 14148 22924 14154 22976
rect 16853 22967 16911 22973
rect 16853 22933 16865 22967
rect 16899 22964 16911 22967
rect 17402 22964 17408 22976
rect 16899 22936 17408 22964
rect 16899 22933 16911 22936
rect 16853 22927 16911 22933
rect 17402 22924 17408 22936
rect 17460 22924 17466 22976
rect 20898 22964 20904 22976
rect 20859 22936 20904 22964
rect 20898 22924 20904 22936
rect 20956 22924 20962 22976
rect 21910 22964 21916 22976
rect 21871 22936 21916 22964
rect 21910 22924 21916 22936
rect 21968 22924 21974 22976
rect 25225 22967 25283 22973
rect 25225 22933 25237 22967
rect 25271 22964 25283 22967
rect 25314 22964 25320 22976
rect 25271 22936 25320 22964
rect 25271 22933 25283 22936
rect 25225 22927 25283 22933
rect 25314 22924 25320 22936
rect 25372 22924 25378 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 10594 22760 10600 22772
rect 10555 22732 10600 22760
rect 10594 22720 10600 22732
rect 10652 22720 10658 22772
rect 10778 22760 10784 22772
rect 10739 22732 10784 22760
rect 10778 22720 10784 22732
rect 10836 22720 10842 22772
rect 11790 22720 11796 22772
rect 11848 22760 11854 22772
rect 11885 22763 11943 22769
rect 11885 22760 11897 22763
rect 11848 22732 11897 22760
rect 11848 22720 11854 22732
rect 11885 22729 11897 22732
rect 11931 22760 11943 22763
rect 12253 22763 12311 22769
rect 12253 22760 12265 22763
rect 11931 22732 12265 22760
rect 11931 22729 11943 22732
rect 11885 22723 11943 22729
rect 12253 22729 12265 22732
rect 12299 22760 12311 22763
rect 12710 22760 12716 22772
rect 12299 22732 12716 22760
rect 12299 22729 12311 22732
rect 12253 22723 12311 22729
rect 12710 22720 12716 22732
rect 12768 22720 12774 22772
rect 16574 22720 16580 22772
rect 16632 22760 16638 22772
rect 16853 22763 16911 22769
rect 16853 22760 16865 22763
rect 16632 22732 16865 22760
rect 16632 22720 16638 22732
rect 16853 22729 16865 22732
rect 16899 22729 16911 22763
rect 16853 22723 16911 22729
rect 17497 22763 17555 22769
rect 17497 22729 17509 22763
rect 17543 22760 17555 22763
rect 17586 22760 17592 22772
rect 17543 22732 17592 22760
rect 17543 22729 17555 22732
rect 17497 22723 17555 22729
rect 17586 22720 17592 22732
rect 17644 22720 17650 22772
rect 17862 22760 17868 22772
rect 17775 22732 17868 22760
rect 17862 22720 17868 22732
rect 17920 22760 17926 22772
rect 18414 22760 18420 22772
rect 17920 22732 18420 22760
rect 17920 22720 17926 22732
rect 18414 22720 18420 22732
rect 18472 22720 18478 22772
rect 20990 22760 20996 22772
rect 20951 22732 20996 22760
rect 20990 22720 20996 22732
rect 21048 22720 21054 22772
rect 23477 22763 23535 22769
rect 23477 22729 23489 22763
rect 23523 22760 23535 22763
rect 23566 22760 23572 22772
rect 23523 22732 23572 22760
rect 23523 22729 23535 22732
rect 23477 22723 23535 22729
rect 23566 22720 23572 22732
rect 23624 22760 23630 22772
rect 23750 22760 23756 22772
rect 23624 22732 23756 22760
rect 23624 22720 23630 22732
rect 23750 22720 23756 22732
rect 23808 22720 23814 22772
rect 25038 22720 25044 22772
rect 25096 22760 25102 22772
rect 25498 22760 25504 22772
rect 25096 22732 25504 22760
rect 25096 22720 25102 22732
rect 25498 22720 25504 22732
rect 25556 22760 25562 22772
rect 25869 22763 25927 22769
rect 25869 22760 25881 22763
rect 25556 22732 25881 22760
rect 25556 22720 25562 22732
rect 25869 22729 25881 22732
rect 25915 22729 25927 22763
rect 25869 22723 25927 22729
rect 10612 22624 10640 22720
rect 11241 22627 11299 22633
rect 11241 22624 11253 22627
rect 10612 22596 11253 22624
rect 11241 22593 11253 22596
rect 11287 22593 11299 22627
rect 11241 22587 11299 22593
rect 11425 22627 11483 22633
rect 11425 22593 11437 22627
rect 11471 22624 11483 22627
rect 11808 22624 11836 22720
rect 11471 22596 11836 22624
rect 11471 22593 11483 22596
rect 11425 22587 11483 22593
rect 10321 22559 10379 22565
rect 10321 22525 10333 22559
rect 10367 22556 10379 22559
rect 11146 22556 11152 22568
rect 10367 22528 11152 22556
rect 10367 22525 10379 22528
rect 10321 22519 10379 22525
rect 11146 22516 11152 22528
rect 11204 22516 11210 22568
rect 11256 22556 11284 22587
rect 14642 22584 14648 22636
rect 14700 22624 14706 22636
rect 14921 22627 14979 22633
rect 14921 22624 14933 22627
rect 14700 22596 14933 22624
rect 14700 22584 14706 22596
rect 14921 22593 14933 22596
rect 14967 22593 14979 22627
rect 14921 22587 14979 22593
rect 18601 22627 18659 22633
rect 18601 22593 18613 22627
rect 18647 22624 18659 22627
rect 18969 22627 19027 22633
rect 18969 22624 18981 22627
rect 18647 22596 18981 22624
rect 18647 22593 18659 22596
rect 18601 22587 18659 22593
rect 18969 22593 18981 22596
rect 19015 22624 19027 22627
rect 21361 22627 21419 22633
rect 21361 22624 21373 22627
rect 19015 22596 19196 22624
rect 19015 22593 19027 22596
rect 18969 22587 19027 22593
rect 11882 22556 11888 22568
rect 11256 22528 11888 22556
rect 11882 22516 11888 22528
rect 11940 22516 11946 22568
rect 12710 22565 12716 22568
rect 12437 22559 12495 22565
rect 12437 22525 12449 22559
rect 12483 22556 12495 22559
rect 12483 22528 12572 22556
rect 12483 22525 12495 22528
rect 12437 22519 12495 22525
rect 9677 22491 9735 22497
rect 9677 22457 9689 22491
rect 9723 22488 9735 22491
rect 9858 22488 9864 22500
rect 9723 22460 9864 22488
rect 9723 22457 9735 22460
rect 9677 22451 9735 22457
rect 9858 22448 9864 22460
rect 9916 22448 9922 22500
rect 12544 22488 12572 22528
rect 12704 22519 12716 22565
rect 12768 22556 12774 22568
rect 19058 22556 19064 22568
rect 12768 22528 12804 22556
rect 19019 22528 19064 22556
rect 12710 22516 12716 22519
rect 12768 22516 12774 22528
rect 19058 22516 19064 22528
rect 19116 22516 19122 22568
rect 19168 22556 19196 22596
rect 20824 22596 21373 22624
rect 19334 22565 19340 22568
rect 19328 22556 19340 22565
rect 19168 22528 19340 22556
rect 19328 22519 19340 22528
rect 19334 22516 19340 22519
rect 19392 22516 19398 22568
rect 19886 22516 19892 22568
rect 19944 22556 19950 22568
rect 20162 22556 20168 22568
rect 19944 22528 20168 22556
rect 19944 22516 19950 22528
rect 20162 22516 20168 22528
rect 20220 22556 20226 22568
rect 20824 22556 20852 22596
rect 21361 22593 21373 22596
rect 21407 22624 21419 22627
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21407 22596 22017 22624
rect 21407 22593 21419 22596
rect 21361 22587 21419 22593
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 22094 22584 22100 22636
rect 22152 22624 22158 22636
rect 23934 22624 23940 22636
rect 22152 22596 22197 22624
rect 23895 22596 23940 22624
rect 22152 22584 22158 22596
rect 23934 22584 23940 22596
rect 23992 22584 23998 22636
rect 20220 22528 20852 22556
rect 20220 22516 20226 22528
rect 21082 22516 21088 22568
rect 21140 22556 21146 22568
rect 21910 22556 21916 22568
rect 21140 22528 21916 22556
rect 21140 22516 21146 22528
rect 21910 22516 21916 22528
rect 21968 22516 21974 22568
rect 22557 22559 22615 22565
rect 22557 22556 22569 22559
rect 22020 22528 22569 22556
rect 12618 22488 12624 22500
rect 12544 22460 12624 22488
rect 12618 22448 12624 22460
rect 12676 22448 12682 22500
rect 15166 22491 15224 22497
rect 15166 22488 15178 22491
rect 14752 22460 15178 22488
rect 9769 22423 9827 22429
rect 9769 22389 9781 22423
rect 9815 22420 9827 22423
rect 10134 22420 10140 22432
rect 9815 22392 10140 22420
rect 9815 22389 9827 22392
rect 9769 22383 9827 22389
rect 10134 22380 10140 22392
rect 10192 22380 10198 22432
rect 13538 22380 13544 22432
rect 13596 22420 13602 22432
rect 14752 22429 14780 22460
rect 15166 22457 15178 22460
rect 15212 22457 15224 22491
rect 15166 22451 15224 22457
rect 20806 22448 20812 22500
rect 20864 22488 20870 22500
rect 22020 22488 22048 22528
rect 22557 22525 22569 22528
rect 22603 22525 22615 22559
rect 23658 22556 23664 22568
rect 23619 22528 23664 22556
rect 22557 22519 22615 22525
rect 23658 22516 23664 22528
rect 23716 22556 23722 22568
rect 24397 22559 24455 22565
rect 24397 22556 24409 22559
rect 23716 22528 24409 22556
rect 23716 22516 23722 22528
rect 24397 22525 24409 22528
rect 24443 22525 24455 22559
rect 24946 22556 24952 22568
rect 24907 22528 24952 22556
rect 24397 22519 24455 22525
rect 24946 22516 24952 22528
rect 25004 22556 25010 22568
rect 25501 22559 25559 22565
rect 25501 22556 25513 22559
rect 25004 22528 25513 22556
rect 25004 22516 25010 22528
rect 25501 22525 25513 22528
rect 25547 22525 25559 22559
rect 25501 22519 25559 22525
rect 20864 22460 22048 22488
rect 20864 22448 20870 22460
rect 13817 22423 13875 22429
rect 13817 22420 13829 22423
rect 13596 22392 13829 22420
rect 13596 22380 13602 22392
rect 13817 22389 13829 22392
rect 13863 22420 13875 22423
rect 14369 22423 14427 22429
rect 14369 22420 14381 22423
rect 13863 22392 14381 22420
rect 13863 22389 13875 22392
rect 13817 22383 13875 22389
rect 14369 22389 14381 22392
rect 14415 22420 14427 22423
rect 14737 22423 14795 22429
rect 14737 22420 14749 22423
rect 14415 22392 14749 22420
rect 14415 22389 14427 22392
rect 14369 22383 14427 22389
rect 14737 22389 14749 22392
rect 14783 22389 14795 22423
rect 14737 22383 14795 22389
rect 14826 22380 14832 22432
rect 14884 22420 14890 22432
rect 16301 22423 16359 22429
rect 16301 22420 16313 22423
rect 14884 22392 16313 22420
rect 14884 22380 14890 22392
rect 16301 22389 16313 22392
rect 16347 22389 16359 22423
rect 18046 22420 18052 22432
rect 18007 22392 18052 22420
rect 16301 22383 16359 22389
rect 18046 22380 18052 22392
rect 18104 22380 18110 22432
rect 20441 22423 20499 22429
rect 20441 22389 20453 22423
rect 20487 22420 20499 22423
rect 20714 22420 20720 22432
rect 20487 22392 20720 22420
rect 20487 22389 20499 22392
rect 20441 22383 20499 22389
rect 20714 22380 20720 22392
rect 20772 22380 20778 22432
rect 21542 22420 21548 22432
rect 21503 22392 21548 22420
rect 21542 22380 21548 22392
rect 21600 22380 21606 22432
rect 22922 22420 22928 22432
rect 22883 22392 22928 22420
rect 22922 22380 22928 22392
rect 22980 22380 22986 22432
rect 24670 22380 24676 22432
rect 24728 22420 24734 22432
rect 25133 22423 25191 22429
rect 25133 22420 25145 22423
rect 24728 22392 25145 22420
rect 24728 22380 24734 22392
rect 25133 22389 25145 22392
rect 25179 22389 25191 22423
rect 25133 22383 25191 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 9858 22176 9864 22228
rect 9916 22216 9922 22228
rect 10686 22216 10692 22228
rect 9916 22188 10692 22216
rect 9916 22176 9922 22188
rect 10686 22176 10692 22188
rect 10744 22216 10750 22228
rect 11057 22219 11115 22225
rect 11057 22216 11069 22219
rect 10744 22188 11069 22216
rect 10744 22176 10750 22188
rect 11057 22185 11069 22188
rect 11103 22185 11115 22219
rect 12250 22216 12256 22228
rect 12211 22188 12256 22216
rect 11057 22179 11115 22185
rect 12250 22176 12256 22188
rect 12308 22176 12314 22228
rect 12986 22216 12992 22228
rect 12899 22188 12992 22216
rect 12986 22176 12992 22188
rect 13044 22216 13050 22228
rect 13262 22216 13268 22228
rect 13044 22188 13268 22216
rect 13044 22176 13050 22188
rect 13262 22176 13268 22188
rect 13320 22176 13326 22228
rect 16022 22216 16028 22228
rect 15983 22188 16028 22216
rect 16022 22176 16028 22188
rect 16080 22176 16086 22228
rect 16574 22176 16580 22228
rect 16632 22216 16638 22228
rect 17313 22219 17371 22225
rect 17313 22216 17325 22219
rect 16632 22188 17325 22216
rect 16632 22176 16638 22188
rect 17313 22185 17325 22188
rect 17359 22185 17371 22219
rect 17313 22179 17371 22185
rect 19518 22176 19524 22228
rect 19576 22216 19582 22228
rect 19613 22219 19671 22225
rect 19613 22216 19625 22219
rect 19576 22188 19625 22216
rect 19576 22176 19582 22188
rect 19613 22185 19625 22188
rect 19659 22216 19671 22219
rect 20898 22216 20904 22228
rect 19659 22188 20904 22216
rect 19659 22185 19671 22188
rect 19613 22179 19671 22185
rect 20898 22176 20904 22188
rect 20956 22176 20962 22228
rect 8573 22151 8631 22157
rect 8573 22117 8585 22151
rect 8619 22148 8631 22151
rect 8619 22120 9628 22148
rect 8619 22117 8631 22120
rect 8573 22111 8631 22117
rect 9600 22080 9628 22120
rect 12894 22108 12900 22160
rect 12952 22148 12958 22160
rect 13725 22151 13783 22157
rect 13725 22148 13737 22151
rect 12952 22120 13737 22148
rect 12952 22108 12958 22120
rect 13725 22117 13737 22120
rect 13771 22117 13783 22151
rect 20254 22148 20260 22160
rect 20215 22120 20260 22148
rect 13725 22111 13783 22117
rect 20254 22108 20260 22120
rect 20312 22108 20318 22160
rect 21542 22148 21548 22160
rect 20640 22120 21548 22148
rect 9766 22080 9772 22092
rect 9600 22052 9772 22080
rect 9766 22040 9772 22052
rect 9824 22040 9830 22092
rect 9944 22083 10002 22089
rect 9944 22049 9956 22083
rect 9990 22080 10002 22083
rect 10226 22080 10232 22092
rect 9990 22052 10232 22080
rect 9990 22049 10002 22052
rect 9944 22043 10002 22049
rect 10226 22040 10232 22052
rect 10284 22040 10290 22092
rect 13262 22040 13268 22092
rect 13320 22080 13326 22092
rect 13633 22083 13691 22089
rect 13633 22080 13645 22083
rect 13320 22052 13645 22080
rect 13320 22040 13326 22052
rect 13633 22049 13645 22052
rect 13679 22049 13691 22083
rect 13998 22080 14004 22092
rect 13633 22043 13691 22049
rect 13924 22052 14004 22080
rect 13924 22021 13952 22052
rect 13998 22040 14004 22052
rect 14056 22080 14062 22092
rect 14826 22080 14832 22092
rect 14056 22052 14832 22080
rect 14056 22040 14062 22052
rect 14826 22040 14832 22052
rect 14884 22040 14890 22092
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22049 15347 22083
rect 15289 22043 15347 22049
rect 17221 22083 17279 22089
rect 17221 22049 17233 22083
rect 17267 22080 17279 22083
rect 17310 22080 17316 22092
rect 17267 22052 17316 22080
rect 17267 22049 17279 22052
rect 17221 22043 17279 22049
rect 9677 22015 9735 22021
rect 9677 22012 9689 22015
rect 9416 21984 9689 22012
rect 8202 21876 8208 21888
rect 8163 21848 8208 21876
rect 8202 21836 8208 21848
rect 8260 21876 8266 21888
rect 9416 21885 9444 21984
rect 9677 21981 9689 21984
rect 9723 21981 9735 22015
rect 9677 21975 9735 21981
rect 13909 22015 13967 22021
rect 13909 21981 13921 22015
rect 13955 21981 13967 22015
rect 13909 21975 13967 21981
rect 13265 21947 13323 21953
rect 13265 21913 13277 21947
rect 13311 21944 13323 21947
rect 15304 21944 15332 22043
rect 17310 22040 17316 22052
rect 17368 22040 17374 22092
rect 19702 22080 19708 22092
rect 19615 22052 19708 22080
rect 19702 22040 19708 22052
rect 19760 22080 19766 22092
rect 20640 22080 20668 22120
rect 21542 22108 21548 22120
rect 21600 22108 21606 22160
rect 19760 22052 20668 22080
rect 19760 22040 19766 22052
rect 20714 22040 20720 22092
rect 20772 22080 20778 22092
rect 21157 22083 21215 22089
rect 21157 22080 21169 22083
rect 20772 22052 21169 22080
rect 20772 22040 20778 22052
rect 21157 22049 21169 22052
rect 21203 22080 21215 22083
rect 21450 22080 21456 22092
rect 21203 22052 21456 22080
rect 21203 22049 21215 22052
rect 21157 22043 21215 22049
rect 21450 22040 21456 22052
rect 21508 22040 21514 22092
rect 23750 22080 23756 22092
rect 23711 22052 23756 22080
rect 23750 22040 23756 22052
rect 23808 22040 23814 22092
rect 24026 22080 24032 22092
rect 23987 22052 24032 22080
rect 24026 22040 24032 22052
rect 24084 22040 24090 22092
rect 25038 22080 25044 22092
rect 24999 22052 25044 22080
rect 25038 22040 25044 22052
rect 25096 22040 25102 22092
rect 15562 22012 15568 22024
rect 15523 21984 15568 22012
rect 15562 21972 15568 21984
rect 15620 21972 15626 22024
rect 17402 22012 17408 22024
rect 17363 21984 17408 22012
rect 17402 21972 17408 21984
rect 17460 21972 17466 22024
rect 19886 22012 19892 22024
rect 19847 21984 19892 22012
rect 19886 21972 19892 21984
rect 19944 21972 19950 22024
rect 20070 21972 20076 22024
rect 20128 21972 20134 22024
rect 20898 22012 20904 22024
rect 20859 21984 20904 22012
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 15470 21944 15476 21956
rect 13311 21916 15476 21944
rect 13311 21913 13323 21916
rect 13265 21907 13323 21913
rect 15470 21904 15476 21916
rect 15528 21904 15534 21956
rect 16853 21947 16911 21953
rect 16853 21913 16865 21947
rect 16899 21944 16911 21947
rect 17862 21944 17868 21956
rect 16899 21916 17868 21944
rect 16899 21913 16911 21916
rect 16853 21907 16911 21913
rect 17862 21904 17868 21916
rect 17920 21904 17926 21956
rect 18506 21904 18512 21956
rect 18564 21944 18570 21956
rect 20088 21944 20116 21972
rect 18564 21916 20116 21944
rect 18564 21904 18570 21916
rect 9401 21879 9459 21885
rect 9401 21876 9413 21879
rect 8260 21848 9413 21876
rect 8260 21836 8266 21848
rect 9401 21845 9413 21848
rect 9447 21876 9459 21879
rect 10042 21876 10048 21888
rect 9447 21848 10048 21876
rect 9447 21845 9459 21848
rect 9401 21839 9459 21845
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 14458 21876 14464 21888
rect 14419 21848 14464 21876
rect 14458 21836 14464 21848
rect 14516 21876 14522 21888
rect 14642 21876 14648 21888
rect 14516 21848 14648 21876
rect 14516 21836 14522 21848
rect 14642 21836 14648 21848
rect 14700 21836 14706 21888
rect 14734 21836 14740 21888
rect 14792 21876 14798 21888
rect 14829 21879 14887 21885
rect 14829 21876 14841 21879
rect 14792 21848 14841 21876
rect 14792 21836 14798 21848
rect 14829 21845 14841 21848
rect 14875 21845 14887 21879
rect 14829 21839 14887 21845
rect 16485 21879 16543 21885
rect 16485 21845 16497 21879
rect 16531 21876 16543 21879
rect 16942 21876 16948 21888
rect 16531 21848 16948 21876
rect 16531 21845 16543 21848
rect 16485 21839 16543 21845
rect 16942 21836 16948 21848
rect 17000 21836 17006 21888
rect 18138 21876 18144 21888
rect 18099 21848 18144 21876
rect 18138 21836 18144 21848
rect 18196 21836 18202 21888
rect 19058 21876 19064 21888
rect 19019 21848 19064 21876
rect 19058 21836 19064 21848
rect 19116 21836 19122 21888
rect 19242 21876 19248 21888
rect 19203 21848 19248 21876
rect 19242 21836 19248 21848
rect 19300 21836 19306 21888
rect 20070 21836 20076 21888
rect 20128 21876 20134 21888
rect 20625 21879 20683 21885
rect 20625 21876 20637 21879
rect 20128 21848 20637 21876
rect 20128 21836 20134 21848
rect 20625 21845 20637 21848
rect 20671 21876 20683 21879
rect 20714 21876 20720 21888
rect 20671 21848 20720 21876
rect 20671 21845 20683 21848
rect 20625 21839 20683 21845
rect 20714 21836 20720 21848
rect 20772 21836 20778 21888
rect 22278 21876 22284 21888
rect 22239 21848 22284 21876
rect 22278 21836 22284 21848
rect 22336 21836 22342 21888
rect 24854 21836 24860 21888
rect 24912 21876 24918 21888
rect 25225 21879 25283 21885
rect 25225 21876 25237 21879
rect 24912 21848 25237 21876
rect 24912 21836 24918 21848
rect 25225 21845 25237 21848
rect 25271 21845 25283 21879
rect 25225 21839 25283 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 12710 21672 12716 21684
rect 12671 21644 12716 21672
rect 12710 21632 12716 21644
rect 12768 21632 12774 21684
rect 13262 21672 13268 21684
rect 13223 21644 13268 21672
rect 13262 21632 13268 21644
rect 13320 21632 13326 21684
rect 13998 21632 14004 21684
rect 14056 21672 14062 21684
rect 14277 21675 14335 21681
rect 14277 21672 14289 21675
rect 14056 21644 14289 21672
rect 14056 21632 14062 21644
rect 14277 21641 14289 21644
rect 14323 21641 14335 21675
rect 14277 21635 14335 21641
rect 16301 21675 16359 21681
rect 16301 21641 16313 21675
rect 16347 21672 16359 21675
rect 17402 21672 17408 21684
rect 16347 21644 17408 21672
rect 16347 21641 16359 21644
rect 16301 21635 16359 21641
rect 17402 21632 17408 21644
rect 17460 21632 17466 21684
rect 19702 21672 19708 21684
rect 19663 21644 19708 21672
rect 19702 21632 19708 21644
rect 19760 21632 19766 21684
rect 20070 21672 20076 21684
rect 20031 21644 20076 21672
rect 20070 21632 20076 21644
rect 20128 21632 20134 21684
rect 20898 21632 20904 21684
rect 20956 21672 20962 21684
rect 21266 21672 21272 21684
rect 20956 21644 21272 21672
rect 20956 21632 20962 21644
rect 21266 21632 21272 21644
rect 21324 21672 21330 21684
rect 22465 21675 22523 21681
rect 22465 21672 22477 21675
rect 21324 21644 22477 21672
rect 21324 21632 21330 21644
rect 22465 21641 22477 21644
rect 22511 21641 22523 21675
rect 25038 21672 25044 21684
rect 24999 21644 25044 21672
rect 22465 21635 22523 21641
rect 25038 21632 25044 21644
rect 25096 21632 25102 21684
rect 12253 21607 12311 21613
rect 12253 21573 12265 21607
rect 12299 21604 12311 21607
rect 13280 21604 13308 21632
rect 12299 21576 13308 21604
rect 12299 21573 12311 21576
rect 12253 21567 12311 21573
rect 10597 21539 10655 21545
rect 10597 21505 10609 21539
rect 10643 21536 10655 21539
rect 11146 21536 11152 21548
rect 10643 21508 11152 21536
rect 10643 21505 10655 21508
rect 10597 21499 10655 21505
rect 11146 21496 11152 21508
rect 11204 21496 11210 21548
rect 11241 21539 11299 21545
rect 11241 21505 11253 21539
rect 11287 21505 11299 21539
rect 11241 21499 11299 21505
rect 7650 21428 7656 21480
rect 7708 21468 7714 21480
rect 8202 21468 8208 21480
rect 7708 21440 8208 21468
rect 7708 21428 7714 21440
rect 8202 21428 8208 21440
rect 8260 21428 8266 21480
rect 10134 21428 10140 21480
rect 10192 21468 10198 21480
rect 10229 21471 10287 21477
rect 10229 21468 10241 21471
rect 10192 21440 10241 21468
rect 10192 21428 10198 21440
rect 10229 21437 10241 21440
rect 10275 21468 10287 21471
rect 11256 21468 11284 21499
rect 13078 21496 13084 21548
rect 13136 21536 13142 21548
rect 13262 21536 13268 21548
rect 13136 21508 13268 21536
rect 13136 21496 13142 21508
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 13538 21496 13544 21548
rect 13596 21536 13602 21548
rect 13817 21539 13875 21545
rect 13817 21536 13829 21539
rect 13596 21508 13829 21536
rect 13596 21496 13602 21508
rect 13817 21505 13829 21508
rect 13863 21505 13875 21539
rect 13817 21499 13875 21505
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21505 15531 21539
rect 16942 21536 16948 21548
rect 16903 21508 16948 21536
rect 15473 21499 15531 21505
rect 10275 21440 11284 21468
rect 10275 21437 10287 21440
rect 10229 21431 10287 21437
rect 12710 21428 12716 21480
rect 12768 21468 12774 21480
rect 13633 21471 13691 21477
rect 13633 21468 13645 21471
rect 12768 21440 13645 21468
rect 12768 21428 12774 21440
rect 13633 21437 13645 21440
rect 13679 21437 13691 21471
rect 13633 21431 13691 21437
rect 14734 21428 14740 21480
rect 14792 21468 14798 21480
rect 15197 21471 15255 21477
rect 15197 21468 15209 21471
rect 14792 21440 15209 21468
rect 14792 21428 14798 21440
rect 15197 21437 15209 21440
rect 15243 21437 15255 21471
rect 15488 21468 15516 21499
rect 16942 21496 16948 21508
rect 17000 21496 17006 21548
rect 18138 21496 18144 21548
rect 18196 21536 18202 21548
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 18196 21508 18705 21536
rect 18196 21496 18202 21508
rect 18693 21505 18705 21508
rect 18739 21536 18751 21539
rect 19150 21536 19156 21548
rect 18739 21508 19156 21536
rect 18739 21505 18751 21508
rect 18693 21499 18751 21505
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 19337 21539 19395 21545
rect 19337 21505 19349 21539
rect 19383 21536 19395 21539
rect 19886 21536 19892 21548
rect 19383 21508 19892 21536
rect 19383 21505 19395 21508
rect 19337 21499 19395 21505
rect 19886 21496 19892 21508
rect 19944 21536 19950 21548
rect 20441 21539 20499 21545
rect 20441 21536 20453 21539
rect 19944 21508 20453 21536
rect 19944 21496 19950 21508
rect 20441 21505 20453 21508
rect 20487 21536 20499 21539
rect 24210 21536 24216 21548
rect 20487 21508 20668 21536
rect 24171 21508 24216 21536
rect 20487 21505 20499 21508
rect 20441 21499 20499 21505
rect 15933 21471 15991 21477
rect 15933 21468 15945 21471
rect 15488 21440 15945 21468
rect 15197 21431 15255 21437
rect 15933 21437 15945 21440
rect 15979 21468 15991 21471
rect 16390 21468 16396 21480
rect 15979 21440 16396 21468
rect 15979 21437 15991 21440
rect 15933 21431 15991 21437
rect 16390 21428 16396 21440
rect 16448 21428 16454 21480
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 18417 21471 18475 21477
rect 18417 21468 18429 21471
rect 18104 21440 18429 21468
rect 18104 21428 18110 21440
rect 18417 21437 18429 21440
rect 18463 21437 18475 21471
rect 18417 21431 18475 21437
rect 19058 21428 19064 21480
rect 19116 21468 19122 21480
rect 20530 21468 20536 21480
rect 19116 21440 20536 21468
rect 19116 21428 19122 21440
rect 20530 21428 20536 21440
rect 20588 21428 20594 21480
rect 20640 21468 20668 21508
rect 24210 21496 24216 21508
rect 24268 21496 24274 21548
rect 25498 21536 25504 21548
rect 25459 21508 25504 21536
rect 25498 21496 25504 21508
rect 25556 21496 25562 21548
rect 20800 21471 20858 21477
rect 20800 21468 20812 21471
rect 20640 21440 20812 21468
rect 20800 21437 20812 21440
rect 20846 21468 20858 21471
rect 22278 21468 22284 21480
rect 20846 21440 22284 21468
rect 20846 21437 20858 21440
rect 20800 21431 20858 21437
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 23934 21468 23940 21480
rect 23847 21440 23940 21468
rect 23934 21428 23940 21440
rect 23992 21468 23998 21480
rect 24673 21471 24731 21477
rect 24673 21468 24685 21471
rect 23992 21440 24685 21468
rect 23992 21428 23998 21440
rect 24673 21437 24685 21440
rect 24719 21437 24731 21471
rect 25222 21468 25228 21480
rect 25183 21440 25228 21468
rect 24673 21431 24731 21437
rect 25222 21428 25228 21440
rect 25280 21468 25286 21480
rect 25961 21471 26019 21477
rect 25961 21468 25973 21471
rect 25280 21440 25973 21468
rect 25280 21428 25286 21440
rect 25961 21437 25973 21440
rect 26007 21437 26019 21471
rect 25961 21431 26019 21437
rect 8478 21409 8484 21412
rect 8113 21403 8171 21409
rect 8113 21369 8125 21403
rect 8159 21400 8171 21403
rect 8472 21400 8484 21409
rect 8159 21372 8484 21400
rect 8159 21369 8171 21372
rect 8113 21363 8171 21369
rect 8472 21363 8484 21372
rect 8478 21360 8484 21363
rect 8536 21360 8542 21412
rect 12802 21360 12808 21412
rect 12860 21400 12866 21412
rect 12986 21400 12992 21412
rect 12860 21372 12992 21400
rect 12860 21360 12866 21372
rect 12986 21360 12992 21372
rect 13044 21360 13050 21412
rect 14642 21400 14648 21412
rect 14603 21372 14648 21400
rect 14642 21360 14648 21372
rect 14700 21400 14706 21412
rect 15289 21403 15347 21409
rect 15289 21400 15301 21403
rect 14700 21372 15301 21400
rect 14700 21360 14706 21372
rect 15289 21369 15301 21372
rect 15335 21369 15347 21403
rect 15289 21363 15347 21369
rect 17218 21360 17224 21412
rect 17276 21400 17282 21412
rect 17773 21403 17831 21409
rect 17773 21400 17785 21403
rect 17276 21372 17785 21400
rect 17276 21360 17282 21372
rect 17773 21369 17785 21372
rect 17819 21400 17831 21403
rect 18506 21400 18512 21412
rect 17819 21372 18512 21400
rect 17819 21369 17831 21372
rect 17773 21363 17831 21369
rect 18506 21360 18512 21372
rect 18564 21360 18570 21412
rect 9585 21335 9643 21341
rect 9585 21301 9597 21335
rect 9631 21332 9643 21335
rect 10134 21332 10140 21344
rect 9631 21304 10140 21332
rect 9631 21301 9643 21304
rect 9585 21295 9643 21301
rect 10134 21292 10140 21304
rect 10192 21292 10198 21344
rect 10686 21332 10692 21344
rect 10647 21304 10692 21332
rect 10686 21292 10692 21304
rect 10744 21292 10750 21344
rect 11054 21332 11060 21344
rect 11015 21304 11060 21332
rect 11054 21292 11060 21304
rect 11112 21292 11118 21344
rect 12618 21292 12624 21344
rect 12676 21332 12682 21344
rect 13081 21335 13139 21341
rect 13081 21332 13093 21335
rect 12676 21304 13093 21332
rect 12676 21292 12682 21304
rect 13081 21301 13093 21304
rect 13127 21332 13139 21335
rect 13725 21335 13783 21341
rect 13725 21332 13737 21335
rect 13127 21304 13737 21332
rect 13127 21301 13139 21304
rect 13081 21295 13139 21301
rect 13725 21301 13737 21304
rect 13771 21301 13783 21335
rect 14826 21332 14832 21344
rect 14787 21304 14832 21332
rect 13725 21295 13783 21301
rect 14826 21292 14832 21304
rect 14884 21292 14890 21344
rect 16393 21335 16451 21341
rect 16393 21301 16405 21335
rect 16439 21332 16451 21335
rect 16482 21332 16488 21344
rect 16439 21304 16488 21332
rect 16439 21301 16451 21304
rect 16393 21295 16451 21301
rect 16482 21292 16488 21304
rect 16540 21292 16546 21344
rect 16758 21332 16764 21344
rect 16719 21304 16764 21332
rect 16758 21292 16764 21304
rect 16816 21292 16822 21344
rect 16850 21292 16856 21344
rect 16908 21332 16914 21344
rect 16908 21304 16953 21332
rect 16908 21292 16914 21304
rect 17310 21292 17316 21344
rect 17368 21332 17374 21344
rect 17405 21335 17463 21341
rect 17405 21332 17417 21335
rect 17368 21304 17417 21332
rect 17368 21292 17374 21304
rect 17405 21301 17417 21304
rect 17451 21301 17463 21335
rect 17405 21295 17463 21301
rect 18049 21335 18107 21341
rect 18049 21301 18061 21335
rect 18095 21332 18107 21335
rect 18414 21332 18420 21344
rect 18095 21304 18420 21332
rect 18095 21301 18107 21304
rect 18049 21295 18107 21301
rect 18414 21292 18420 21304
rect 18472 21292 18478 21344
rect 21910 21332 21916 21344
rect 21871 21304 21916 21332
rect 21910 21292 21916 21304
rect 21968 21292 21974 21344
rect 23477 21335 23535 21341
rect 23477 21301 23489 21335
rect 23523 21332 23535 21335
rect 23750 21332 23756 21344
rect 23523 21304 23756 21332
rect 23523 21301 23535 21304
rect 23477 21295 23535 21301
rect 23750 21292 23756 21304
rect 23808 21292 23814 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 8202 21128 8208 21140
rect 8163 21100 8208 21128
rect 8202 21088 8208 21100
rect 8260 21088 8266 21140
rect 9766 21088 9772 21140
rect 9824 21128 9830 21140
rect 10689 21131 10747 21137
rect 10689 21128 10701 21131
rect 9824 21100 10701 21128
rect 9824 21088 9830 21100
rect 10689 21097 10701 21100
rect 10735 21128 10747 21131
rect 11054 21128 11060 21140
rect 10735 21100 11060 21128
rect 10735 21097 10747 21100
rect 10689 21091 10747 21097
rect 11054 21088 11060 21100
rect 11112 21088 11118 21140
rect 12894 21128 12900 21140
rect 12855 21100 12900 21128
rect 12894 21088 12900 21100
rect 12952 21088 12958 21140
rect 12986 21088 12992 21140
rect 13044 21128 13050 21140
rect 13446 21128 13452 21140
rect 13044 21100 13452 21128
rect 13044 21088 13050 21100
rect 13446 21088 13452 21100
rect 13504 21088 13510 21140
rect 13538 21088 13544 21140
rect 13596 21128 13602 21140
rect 14093 21131 14151 21137
rect 14093 21128 14105 21131
rect 13596 21100 14105 21128
rect 13596 21088 13602 21100
rect 14093 21097 14105 21100
rect 14139 21097 14151 21131
rect 14093 21091 14151 21097
rect 14826 21088 14832 21140
rect 14884 21128 14890 21140
rect 15933 21131 15991 21137
rect 15933 21128 15945 21131
rect 14884 21100 15945 21128
rect 14884 21088 14890 21100
rect 15933 21097 15945 21100
rect 15979 21128 15991 21131
rect 16850 21128 16856 21140
rect 15979 21100 16856 21128
rect 15979 21097 15991 21100
rect 15933 21091 15991 21097
rect 16850 21088 16856 21100
rect 16908 21088 16914 21140
rect 16942 21088 16948 21140
rect 17000 21128 17006 21140
rect 17402 21128 17408 21140
rect 17000 21100 17408 21128
rect 17000 21088 17006 21100
rect 17402 21088 17408 21100
rect 17460 21128 17466 21140
rect 17497 21131 17555 21137
rect 17497 21128 17509 21131
rect 17460 21100 17509 21128
rect 17460 21088 17466 21100
rect 17497 21097 17509 21100
rect 17543 21097 17555 21131
rect 18046 21128 18052 21140
rect 18007 21100 18052 21128
rect 17497 21091 17555 21097
rect 18046 21088 18052 21100
rect 18104 21088 18110 21140
rect 18138 21088 18144 21140
rect 18196 21128 18202 21140
rect 18509 21131 18567 21137
rect 18509 21128 18521 21131
rect 18196 21100 18521 21128
rect 18196 21088 18202 21100
rect 18509 21097 18521 21100
rect 18555 21128 18567 21131
rect 19058 21128 19064 21140
rect 18555 21100 19064 21128
rect 18555 21097 18567 21100
rect 18509 21091 18567 21097
rect 19058 21088 19064 21100
rect 19116 21088 19122 21140
rect 19518 21088 19524 21140
rect 19576 21128 19582 21140
rect 19613 21131 19671 21137
rect 19613 21128 19625 21131
rect 19576 21100 19625 21128
rect 19576 21088 19582 21100
rect 19613 21097 19625 21100
rect 19659 21097 19671 21131
rect 19613 21091 19671 21097
rect 20349 21131 20407 21137
rect 20349 21097 20361 21131
rect 20395 21128 20407 21131
rect 20530 21128 20536 21140
rect 20395 21100 20536 21128
rect 20395 21097 20407 21100
rect 20349 21091 20407 21097
rect 20530 21088 20536 21100
rect 20588 21088 20594 21140
rect 22646 21128 22652 21140
rect 22607 21100 22652 21128
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 23569 21131 23627 21137
rect 23569 21097 23581 21131
rect 23615 21128 23627 21131
rect 23934 21128 23940 21140
rect 23615 21100 23940 21128
rect 23615 21097 23627 21100
rect 23569 21091 23627 21097
rect 23934 21088 23940 21100
rect 23992 21088 23998 21140
rect 9493 21063 9551 21069
rect 9493 21029 9505 21063
rect 9539 21060 9551 21063
rect 9858 21060 9864 21072
rect 9539 21032 9864 21060
rect 9539 21029 9551 21032
rect 9493 21023 9551 21029
rect 9858 21020 9864 21032
rect 9916 21060 9922 21072
rect 10134 21060 10140 21072
rect 9916 21032 10140 21060
rect 9916 21020 9922 21032
rect 10134 21020 10140 21032
rect 10192 21020 10198 21072
rect 15470 21060 15476 21072
rect 15431 21032 15476 21060
rect 15470 21020 15476 21032
rect 15528 21020 15534 21072
rect 9766 20952 9772 21004
rect 9824 20992 9830 21004
rect 10045 20995 10103 21001
rect 10045 20992 10057 20995
rect 9824 20964 10057 20992
rect 9824 20952 9830 20964
rect 10045 20961 10057 20964
rect 10091 20961 10103 20995
rect 10152 20992 10180 21020
rect 11238 20992 11244 21004
rect 10152 20964 10272 20992
rect 11199 20964 11244 20992
rect 10045 20955 10103 20961
rect 7098 20884 7104 20936
rect 7156 20924 7162 20936
rect 8294 20924 8300 20936
rect 7156 20896 8300 20924
rect 7156 20884 7162 20896
rect 8294 20884 8300 20896
rect 8352 20884 8358 20936
rect 8478 20924 8484 20936
rect 8439 20896 8484 20924
rect 8478 20884 8484 20896
rect 8536 20884 8542 20936
rect 10244 20933 10272 20964
rect 11238 20952 11244 20964
rect 11296 20952 11302 21004
rect 12250 20952 12256 21004
rect 12308 20992 12314 21004
rect 13449 20995 13507 21001
rect 13449 20992 13461 20995
rect 12308 20964 13461 20992
rect 12308 20952 12314 20964
rect 13449 20961 13461 20964
rect 13495 20961 13507 20995
rect 13449 20955 13507 20961
rect 14734 20952 14740 21004
rect 14792 20992 14798 21004
rect 16390 21001 16396 21004
rect 14829 20995 14887 21001
rect 14829 20992 14841 20995
rect 14792 20964 14841 20992
rect 14792 20952 14798 20964
rect 14829 20961 14841 20964
rect 14875 20961 14887 20995
rect 16384 20992 16396 21001
rect 16351 20964 16396 20992
rect 14829 20955 14887 20961
rect 16384 20955 16396 20964
rect 16390 20952 16396 20955
rect 16448 20952 16454 21004
rect 17954 20952 17960 21004
rect 18012 20992 18018 21004
rect 18969 20995 19027 21001
rect 18969 20992 18981 20995
rect 18012 20964 18981 20992
rect 18012 20952 18018 20964
rect 18969 20961 18981 20964
rect 19015 20961 19027 20995
rect 18969 20955 19027 20961
rect 19058 20952 19064 21004
rect 19116 20992 19122 21004
rect 21269 20995 21327 21001
rect 21269 20992 21281 20995
rect 19116 20964 19161 20992
rect 20824 20964 21281 20992
rect 19116 20952 19122 20964
rect 10137 20927 10195 20933
rect 10137 20893 10149 20927
rect 10183 20893 10195 20927
rect 10137 20887 10195 20893
rect 10229 20927 10287 20933
rect 10229 20893 10241 20927
rect 10275 20893 10287 20927
rect 11514 20924 11520 20936
rect 11475 20896 11520 20924
rect 10229 20887 10287 20893
rect 7837 20859 7895 20865
rect 7837 20825 7849 20859
rect 7883 20856 7895 20859
rect 10152 20856 10180 20887
rect 11514 20884 11520 20896
rect 11572 20884 11578 20936
rect 13170 20884 13176 20936
rect 13228 20924 13234 20936
rect 13354 20924 13360 20936
rect 13228 20896 13360 20924
rect 13228 20884 13234 20896
rect 13354 20884 13360 20896
rect 13412 20924 13418 20936
rect 13541 20927 13599 20933
rect 13541 20924 13553 20927
rect 13412 20896 13553 20924
rect 13412 20884 13418 20896
rect 13541 20893 13553 20896
rect 13587 20893 13599 20927
rect 13722 20924 13728 20936
rect 13683 20896 13728 20924
rect 13541 20887 13599 20893
rect 13722 20884 13728 20896
rect 13780 20884 13786 20936
rect 16117 20927 16175 20933
rect 16117 20924 16129 20927
rect 14844 20896 16129 20924
rect 10778 20856 10784 20868
rect 7883 20828 10784 20856
rect 7883 20825 7895 20828
rect 7837 20819 7895 20825
rect 10778 20816 10784 20828
rect 10836 20816 10842 20868
rect 14844 20800 14872 20896
rect 16117 20893 16129 20896
rect 16163 20893 16175 20927
rect 19150 20924 19156 20936
rect 19111 20896 19156 20924
rect 16117 20887 16175 20893
rect 19150 20884 19156 20896
rect 19208 20884 19214 20936
rect 20824 20868 20852 20964
rect 21269 20961 21281 20964
rect 21315 20961 21327 20995
rect 22462 20992 22468 21004
rect 22423 20964 22468 20992
rect 21269 20955 21327 20961
rect 22462 20952 22468 20964
rect 22520 20952 22526 21004
rect 23934 20992 23940 21004
rect 23895 20964 23940 20992
rect 23934 20952 23940 20964
rect 23992 20952 23998 21004
rect 25130 20992 25136 21004
rect 25091 20964 25136 20992
rect 25130 20952 25136 20964
rect 25188 20952 25194 21004
rect 21358 20924 21364 20936
rect 21319 20896 21364 20924
rect 21358 20884 21364 20896
rect 21416 20884 21422 20936
rect 21453 20927 21511 20933
rect 21453 20893 21465 20927
rect 21499 20924 21511 20927
rect 22002 20924 22008 20936
rect 21499 20896 22008 20924
rect 21499 20893 21511 20896
rect 21453 20887 21511 20893
rect 20717 20859 20775 20865
rect 20717 20825 20729 20859
rect 20763 20856 20775 20859
rect 20806 20856 20812 20868
rect 20763 20828 20812 20856
rect 20763 20825 20775 20828
rect 20717 20819 20775 20825
rect 20806 20816 20812 20828
rect 20864 20816 20870 20868
rect 20990 20816 20996 20868
rect 21048 20856 21054 20868
rect 21468 20856 21496 20887
rect 22002 20884 22008 20896
rect 22060 20884 22066 20936
rect 23109 20927 23167 20933
rect 23109 20893 23121 20927
rect 23155 20924 23167 20927
rect 23658 20924 23664 20936
rect 23155 20896 23664 20924
rect 23155 20893 23167 20896
rect 23109 20887 23167 20893
rect 23658 20884 23664 20896
rect 23716 20924 23722 20936
rect 24029 20927 24087 20933
rect 24029 20924 24041 20927
rect 23716 20896 24041 20924
rect 23716 20884 23722 20896
rect 24029 20893 24041 20896
rect 24075 20893 24087 20927
rect 24029 20887 24087 20893
rect 24213 20927 24271 20933
rect 24213 20893 24225 20927
rect 24259 20924 24271 20927
rect 24854 20924 24860 20936
rect 24259 20896 24860 20924
rect 24259 20893 24271 20896
rect 24213 20887 24271 20893
rect 24854 20884 24860 20896
rect 24912 20884 24918 20936
rect 21048 20828 21496 20856
rect 21048 20816 21054 20828
rect 9674 20788 9680 20800
rect 9635 20760 9680 20788
rect 9674 20748 9680 20760
rect 9732 20748 9738 20800
rect 12526 20788 12532 20800
rect 12487 20760 12532 20788
rect 12526 20748 12532 20760
rect 12584 20748 12590 20800
rect 13078 20788 13084 20800
rect 13039 20760 13084 20788
rect 13078 20748 13084 20760
rect 13136 20748 13142 20800
rect 14458 20748 14464 20800
rect 14516 20788 14522 20800
rect 14553 20791 14611 20797
rect 14553 20788 14565 20791
rect 14516 20760 14565 20788
rect 14516 20748 14522 20760
rect 14553 20757 14565 20760
rect 14599 20788 14611 20791
rect 14645 20791 14703 20797
rect 14645 20788 14657 20791
rect 14599 20760 14657 20788
rect 14599 20757 14611 20760
rect 14553 20751 14611 20757
rect 14645 20757 14657 20760
rect 14691 20788 14703 20791
rect 14826 20788 14832 20800
rect 14691 20760 14832 20788
rect 14691 20757 14703 20760
rect 14645 20751 14703 20757
rect 14826 20748 14832 20760
rect 14884 20748 14890 20800
rect 18506 20748 18512 20800
rect 18564 20788 18570 20800
rect 18601 20791 18659 20797
rect 18601 20788 18613 20791
rect 18564 20760 18613 20788
rect 18564 20748 18570 20760
rect 18601 20757 18613 20760
rect 18647 20757 18659 20791
rect 20898 20788 20904 20800
rect 20859 20760 20904 20788
rect 18601 20751 18659 20757
rect 20898 20748 20904 20760
rect 20956 20748 20962 20800
rect 23474 20788 23480 20800
rect 23435 20760 23480 20788
rect 23474 20748 23480 20760
rect 23532 20748 23538 20800
rect 25314 20788 25320 20800
rect 25275 20760 25320 20788
rect 25314 20748 25320 20760
rect 25372 20748 25378 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 7929 20587 7987 20593
rect 7929 20553 7941 20587
rect 7975 20584 7987 20587
rect 8202 20584 8208 20596
rect 7975 20556 8208 20584
rect 7975 20553 7987 20556
rect 7929 20547 7987 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 9677 20587 9735 20593
rect 9677 20553 9689 20587
rect 9723 20553 9735 20587
rect 9677 20547 9735 20553
rect 9692 20516 9720 20547
rect 10686 20544 10692 20596
rect 10744 20584 10750 20596
rect 11057 20587 11115 20593
rect 11057 20584 11069 20587
rect 10744 20556 11069 20584
rect 10744 20544 10750 20556
rect 11057 20553 11069 20556
rect 11103 20553 11115 20587
rect 17402 20584 17408 20596
rect 17363 20556 17408 20584
rect 11057 20547 11115 20553
rect 17402 20544 17408 20556
rect 17460 20544 17466 20596
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 20901 20587 20959 20593
rect 20901 20584 20913 20587
rect 20772 20556 20913 20584
rect 20772 20544 20778 20556
rect 20901 20553 20913 20556
rect 20947 20584 20959 20587
rect 21358 20584 21364 20596
rect 20947 20556 21364 20584
rect 20947 20553 20959 20556
rect 20901 20547 20959 20553
rect 21358 20544 21364 20556
rect 21416 20544 21422 20596
rect 21910 20584 21916 20596
rect 21871 20556 21916 20584
rect 21910 20544 21916 20556
rect 21968 20544 21974 20596
rect 22646 20584 22652 20596
rect 22607 20556 22652 20584
rect 22646 20544 22652 20556
rect 22704 20544 22710 20596
rect 23661 20587 23719 20593
rect 23661 20553 23673 20587
rect 23707 20584 23719 20587
rect 23934 20584 23940 20596
rect 23707 20556 23940 20584
rect 23707 20553 23719 20556
rect 23661 20547 23719 20553
rect 23934 20544 23940 20556
rect 23992 20544 23998 20596
rect 24854 20544 24860 20596
rect 24912 20584 24918 20596
rect 25041 20587 25099 20593
rect 25041 20584 25053 20587
rect 24912 20556 25053 20584
rect 24912 20544 24918 20556
rect 25041 20553 25053 20556
rect 25087 20553 25099 20587
rect 25041 20547 25099 20553
rect 25130 20544 25136 20596
rect 25188 20584 25194 20596
rect 25961 20587 26019 20593
rect 25961 20584 25973 20587
rect 25188 20556 25973 20584
rect 25188 20544 25194 20556
rect 25961 20553 25973 20556
rect 26007 20553 26019 20587
rect 25961 20547 26019 20553
rect 11238 20516 11244 20528
rect 9692 20488 11244 20516
rect 11238 20476 11244 20488
rect 11296 20516 11302 20528
rect 11425 20519 11483 20525
rect 11425 20516 11437 20519
rect 11296 20488 11437 20516
rect 11296 20476 11302 20488
rect 11425 20485 11437 20488
rect 11471 20485 11483 20519
rect 11425 20479 11483 20485
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 10134 20448 10140 20460
rect 9732 20420 10140 20448
rect 9732 20408 9738 20420
rect 10134 20408 10140 20420
rect 10192 20408 10198 20460
rect 10226 20408 10232 20460
rect 10284 20448 10290 20460
rect 10778 20448 10784 20460
rect 10284 20420 10329 20448
rect 10739 20420 10784 20448
rect 10284 20408 10290 20420
rect 10778 20408 10784 20420
rect 10836 20408 10842 20460
rect 17420 20448 17448 20544
rect 20073 20519 20131 20525
rect 20073 20485 20085 20519
rect 20119 20516 20131 20519
rect 20990 20516 20996 20528
rect 20119 20488 20996 20516
rect 20119 20485 20131 20488
rect 20073 20479 20131 20485
rect 20990 20476 20996 20488
rect 21048 20476 21054 20528
rect 21542 20448 21548 20460
rect 17420 20420 18184 20448
rect 21455 20420 21548 20448
rect 9582 20380 9588 20392
rect 9543 20352 9588 20380
rect 9582 20340 9588 20352
rect 9640 20340 9646 20392
rect 10045 20383 10103 20389
rect 10045 20349 10057 20383
rect 10091 20380 10103 20383
rect 10686 20380 10692 20392
rect 10091 20352 10692 20380
rect 10091 20349 10103 20352
rect 10045 20343 10103 20349
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 12437 20383 12495 20389
rect 12437 20380 12449 20383
rect 12360 20352 12449 20380
rect 9217 20315 9275 20321
rect 9217 20281 9229 20315
rect 9263 20312 9275 20315
rect 10226 20312 10232 20324
rect 9263 20284 10232 20312
rect 9263 20281 9275 20284
rect 9217 20275 9275 20281
rect 10226 20272 10232 20284
rect 10284 20272 10290 20324
rect 11885 20315 11943 20321
rect 11885 20281 11897 20315
rect 11931 20312 11943 20315
rect 12360 20312 12388 20352
rect 12437 20349 12449 20352
rect 12483 20349 12495 20383
rect 12437 20343 12495 20349
rect 12526 20340 12532 20392
rect 12584 20380 12590 20392
rect 12693 20383 12751 20389
rect 12693 20380 12705 20383
rect 12584 20352 12705 20380
rect 12584 20340 12590 20352
rect 12693 20349 12705 20352
rect 12739 20349 12751 20383
rect 12693 20343 12751 20349
rect 13814 20340 13820 20392
rect 13872 20380 13878 20392
rect 14369 20383 14427 20389
rect 14369 20380 14381 20383
rect 13872 20352 14381 20380
rect 13872 20340 13878 20352
rect 14369 20349 14381 20352
rect 14415 20349 14427 20383
rect 14918 20380 14924 20392
rect 14879 20352 14924 20380
rect 14369 20343 14427 20349
rect 14918 20340 14924 20352
rect 14976 20340 14982 20392
rect 18046 20380 18052 20392
rect 18007 20352 18052 20380
rect 18046 20340 18052 20352
rect 18104 20340 18110 20392
rect 18156 20380 18184 20420
rect 21542 20408 21548 20420
rect 21600 20448 21606 20460
rect 21928 20448 21956 20544
rect 22373 20519 22431 20525
rect 22373 20485 22385 20519
rect 22419 20516 22431 20519
rect 22462 20516 22468 20528
rect 22419 20488 22468 20516
rect 22419 20485 22431 20488
rect 22373 20479 22431 20485
rect 22462 20476 22468 20488
rect 22520 20516 22526 20528
rect 22520 20488 25452 20516
rect 22520 20476 22526 20488
rect 21600 20420 21956 20448
rect 21600 20408 21606 20420
rect 23474 20408 23480 20460
rect 23532 20448 23538 20460
rect 25424 20457 25452 20488
rect 24213 20451 24271 20457
rect 24213 20448 24225 20451
rect 23532 20420 24225 20448
rect 23532 20408 23538 20420
rect 24213 20417 24225 20420
rect 24259 20417 24271 20451
rect 24213 20411 24271 20417
rect 25409 20451 25467 20457
rect 25409 20417 25421 20451
rect 25455 20417 25467 20451
rect 25409 20411 25467 20417
rect 18305 20383 18363 20389
rect 18305 20380 18317 20383
rect 18156 20352 18317 20380
rect 18305 20349 18317 20352
rect 18351 20349 18363 20383
rect 18305 20343 18363 20349
rect 18690 20340 18696 20392
rect 18748 20380 18754 20392
rect 19058 20380 19064 20392
rect 18748 20352 19064 20380
rect 18748 20340 18754 20352
rect 19058 20340 19064 20352
rect 19116 20380 19122 20392
rect 20349 20383 20407 20389
rect 20349 20380 20361 20383
rect 19116 20352 20361 20380
rect 19116 20340 19122 20352
rect 20349 20349 20361 20352
rect 20395 20380 20407 20383
rect 21269 20383 21327 20389
rect 21269 20380 21281 20383
rect 20395 20352 21281 20380
rect 20395 20349 20407 20352
rect 20349 20343 20407 20349
rect 21269 20349 21281 20352
rect 21315 20349 21327 20383
rect 21269 20343 21327 20349
rect 22465 20383 22523 20389
rect 22465 20349 22477 20383
rect 22511 20380 22523 20383
rect 22830 20380 22836 20392
rect 22511 20352 22836 20380
rect 22511 20349 22523 20352
rect 22465 20343 22523 20349
rect 22830 20340 22836 20352
rect 22888 20380 22894 20392
rect 23017 20383 23075 20389
rect 23017 20380 23029 20383
rect 22888 20352 23029 20380
rect 22888 20340 22894 20352
rect 23017 20349 23029 20352
rect 23063 20349 23075 20383
rect 24121 20383 24179 20389
rect 24121 20380 24133 20383
rect 23017 20343 23075 20349
rect 23860 20352 24133 20380
rect 12802 20312 12808 20324
rect 11931 20284 12808 20312
rect 11931 20281 11943 20284
rect 11885 20275 11943 20281
rect 12802 20272 12808 20284
rect 12860 20272 12866 20324
rect 14829 20315 14887 20321
rect 14829 20281 14841 20315
rect 14875 20312 14887 20315
rect 15166 20315 15224 20321
rect 15166 20312 15178 20315
rect 14875 20284 15178 20312
rect 14875 20281 14887 20284
rect 14829 20275 14887 20281
rect 15166 20281 15178 20284
rect 15212 20312 15224 20315
rect 15838 20312 15844 20324
rect 15212 20284 15844 20312
rect 15212 20281 15224 20284
rect 15166 20275 15224 20281
rect 15838 20272 15844 20284
rect 15896 20312 15902 20324
rect 16666 20312 16672 20324
rect 15896 20284 16672 20312
rect 15896 20272 15902 20284
rect 16666 20272 16672 20284
rect 16724 20272 16730 20324
rect 16945 20315 17003 20321
rect 16945 20281 16957 20315
rect 16991 20312 17003 20315
rect 17034 20312 17040 20324
rect 16991 20284 17040 20312
rect 16991 20281 17003 20284
rect 16945 20275 17003 20281
rect 8294 20244 8300 20256
rect 8255 20216 8300 20244
rect 8294 20204 8300 20216
rect 8352 20204 8358 20256
rect 8478 20204 8484 20256
rect 8536 20244 8542 20256
rect 8665 20247 8723 20253
rect 8665 20244 8677 20247
rect 8536 20216 8677 20244
rect 8536 20204 8542 20216
rect 8665 20213 8677 20216
rect 8711 20244 8723 20247
rect 9030 20244 9036 20256
rect 8711 20216 9036 20244
rect 8711 20213 8723 20216
rect 8665 20207 8723 20213
rect 9030 20204 9036 20216
rect 9088 20204 9094 20256
rect 11422 20204 11428 20256
rect 11480 20244 11486 20256
rect 12161 20247 12219 20253
rect 12161 20244 12173 20247
rect 11480 20216 12173 20244
rect 11480 20204 11486 20216
rect 12161 20213 12173 20216
rect 12207 20244 12219 20247
rect 12250 20244 12256 20256
rect 12207 20216 12256 20244
rect 12207 20213 12219 20216
rect 12161 20207 12219 20213
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 13814 20244 13820 20256
rect 13775 20216 13820 20244
rect 13814 20204 13820 20216
rect 13872 20204 13878 20256
rect 16301 20247 16359 20253
rect 16301 20213 16313 20247
rect 16347 20244 16359 20247
rect 16390 20244 16396 20256
rect 16347 20216 16396 20244
rect 16347 20213 16359 20216
rect 16301 20207 16359 20213
rect 16390 20204 16396 20216
rect 16448 20244 16454 20256
rect 16960 20244 16988 20275
rect 17034 20272 17040 20284
rect 17092 20312 17098 20324
rect 19150 20312 19156 20324
rect 17092 20284 19156 20312
rect 17092 20272 17098 20284
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 20809 20315 20867 20321
rect 20809 20281 20821 20315
rect 20855 20312 20867 20315
rect 20898 20312 20904 20324
rect 20855 20284 20904 20312
rect 20855 20281 20867 20284
rect 20809 20275 20867 20281
rect 20898 20272 20904 20284
rect 20956 20312 20962 20324
rect 21361 20315 21419 20321
rect 21361 20312 21373 20315
rect 20956 20284 21373 20312
rect 20956 20272 20962 20284
rect 21361 20281 21373 20284
rect 21407 20281 21419 20315
rect 21361 20275 21419 20281
rect 23860 20256 23888 20352
rect 24121 20349 24133 20352
rect 24167 20349 24179 20383
rect 25222 20380 25228 20392
rect 25183 20352 25228 20380
rect 24121 20343 24179 20349
rect 25222 20340 25228 20352
rect 25280 20340 25286 20392
rect 24673 20315 24731 20321
rect 24673 20312 24685 20315
rect 24044 20284 24685 20312
rect 24044 20256 24072 20284
rect 24673 20281 24685 20284
rect 24719 20281 24731 20315
rect 24673 20275 24731 20281
rect 17862 20244 17868 20256
rect 16448 20216 16988 20244
rect 17823 20216 17868 20244
rect 16448 20204 16454 20216
rect 17862 20204 17868 20216
rect 17920 20204 17926 20256
rect 18322 20204 18328 20256
rect 18380 20244 18386 20256
rect 19429 20247 19487 20253
rect 19429 20244 19441 20247
rect 18380 20216 19441 20244
rect 18380 20204 18386 20216
rect 19429 20213 19441 20216
rect 19475 20213 19487 20247
rect 19429 20207 19487 20213
rect 23477 20247 23535 20253
rect 23477 20213 23489 20247
rect 23523 20244 23535 20247
rect 23842 20244 23848 20256
rect 23523 20216 23848 20244
rect 23523 20213 23535 20216
rect 23477 20207 23535 20213
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 24026 20244 24032 20256
rect 23987 20216 24032 20244
rect 24026 20204 24032 20216
rect 24084 20204 24090 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 9858 20040 9864 20052
rect 9819 20012 9864 20040
rect 9858 20000 9864 20012
rect 9916 20000 9922 20052
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 10229 20043 10287 20049
rect 10229 20040 10241 20043
rect 10192 20012 10241 20040
rect 10192 20000 10198 20012
rect 10229 20009 10241 20012
rect 10275 20009 10287 20043
rect 13170 20040 13176 20052
rect 13131 20012 13176 20040
rect 10229 20003 10287 20009
rect 13170 20000 13176 20012
rect 13228 20000 13234 20052
rect 16666 20040 16672 20052
rect 16627 20012 16672 20040
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 16758 20000 16764 20052
rect 16816 20040 16822 20052
rect 17221 20043 17279 20049
rect 17221 20040 17233 20043
rect 16816 20012 17233 20040
rect 16816 20000 16822 20012
rect 17221 20009 17233 20012
rect 17267 20009 17279 20043
rect 17221 20003 17279 20009
rect 17773 20043 17831 20049
rect 17773 20009 17785 20043
rect 17819 20040 17831 20043
rect 20714 20040 20720 20052
rect 17819 20012 19380 20040
rect 20675 20012 20720 20040
rect 17819 20009 17831 20012
rect 17773 20003 17831 20009
rect 10870 19981 10876 19984
rect 10864 19972 10876 19981
rect 10831 19944 10876 19972
rect 10864 19935 10876 19944
rect 10870 19932 10876 19935
rect 10928 19932 10934 19984
rect 13078 19932 13084 19984
rect 13136 19972 13142 19984
rect 13817 19975 13875 19981
rect 13817 19972 13829 19975
rect 13136 19944 13829 19972
rect 13136 19932 13142 19944
rect 13817 19941 13829 19944
rect 13863 19941 13875 19975
rect 13817 19935 13875 19941
rect 16574 19932 16580 19984
rect 16632 19972 16638 19984
rect 17589 19975 17647 19981
rect 17589 19972 17601 19975
rect 16632 19944 17601 19972
rect 16632 19932 16638 19944
rect 17589 19941 17601 19944
rect 17635 19972 17647 19975
rect 18233 19975 18291 19981
rect 18233 19972 18245 19975
rect 17635 19944 18245 19972
rect 17635 19941 17647 19944
rect 17589 19935 17647 19941
rect 18233 19941 18245 19944
rect 18279 19941 18291 19975
rect 19150 19972 19156 19984
rect 19111 19944 19156 19972
rect 18233 19935 18291 19941
rect 19150 19932 19156 19944
rect 19208 19932 19214 19984
rect 19352 19916 19380 20012
rect 20714 20000 20720 20012
rect 20772 20000 20778 20052
rect 20898 20000 20904 20052
rect 20956 20040 20962 20052
rect 21266 20040 21272 20052
rect 20956 20012 21272 20040
rect 20956 20000 20962 20012
rect 21266 20000 21272 20012
rect 21324 20040 21330 20052
rect 22002 20040 22008 20052
rect 21324 20012 22008 20040
rect 21324 20000 21330 20012
rect 22002 20000 22008 20012
rect 22060 20000 22066 20052
rect 22094 20000 22100 20052
rect 22152 20040 22158 20052
rect 22281 20043 22339 20049
rect 22281 20040 22293 20043
rect 22152 20012 22293 20040
rect 22152 20000 22158 20012
rect 22281 20009 22293 20012
rect 22327 20009 22339 20043
rect 22281 20003 22339 20009
rect 22925 20043 22983 20049
rect 22925 20009 22937 20043
rect 22971 20040 22983 20043
rect 23934 20040 23940 20052
rect 22971 20012 23940 20040
rect 22971 20009 22983 20012
rect 22925 20003 22983 20009
rect 21168 19975 21226 19981
rect 21168 19941 21180 19975
rect 21214 19972 21226 19975
rect 21542 19972 21548 19984
rect 21214 19944 21548 19972
rect 21214 19941 21226 19944
rect 21168 19935 21226 19941
rect 21542 19932 21548 19944
rect 21600 19932 21606 19984
rect 13722 19904 13728 19916
rect 13683 19876 13728 19904
rect 13722 19864 13728 19876
rect 13780 19864 13786 19916
rect 15378 19904 15384 19916
rect 15212 19876 15384 19904
rect 9674 19796 9680 19848
rect 9732 19836 9738 19848
rect 10597 19839 10655 19845
rect 10597 19836 10609 19839
rect 9732 19808 10609 19836
rect 9732 19796 9738 19808
rect 10597 19805 10609 19808
rect 10643 19805 10655 19839
rect 10597 19799 10655 19805
rect 13446 19796 13452 19848
rect 13504 19836 13510 19848
rect 14001 19839 14059 19845
rect 14001 19836 14013 19839
rect 13504 19808 14013 19836
rect 13504 19796 13510 19808
rect 14001 19805 14013 19808
rect 14047 19836 14059 19839
rect 15212 19836 15240 19876
rect 15378 19864 15384 19876
rect 15436 19904 15442 19916
rect 15545 19907 15603 19913
rect 15545 19904 15557 19907
rect 15436 19876 15557 19904
rect 15436 19864 15442 19876
rect 15545 19873 15557 19876
rect 15591 19873 15603 19907
rect 15545 19867 15603 19873
rect 18046 19864 18052 19916
rect 18104 19904 18110 19916
rect 18141 19907 18199 19913
rect 18141 19904 18153 19907
rect 18104 19876 18153 19904
rect 18104 19864 18110 19876
rect 18141 19873 18153 19876
rect 18187 19873 18199 19907
rect 19334 19904 19340 19916
rect 19247 19876 19340 19904
rect 18141 19867 18199 19873
rect 19334 19864 19340 19876
rect 19392 19864 19398 19916
rect 20530 19864 20536 19916
rect 20588 19904 20594 19916
rect 20898 19904 20904 19916
rect 20588 19876 20904 19904
rect 20588 19864 20594 19876
rect 20898 19864 20904 19876
rect 20956 19864 20962 19916
rect 22296 19904 22324 20003
rect 23934 20000 23940 20012
rect 23992 20000 23998 20052
rect 24765 20043 24823 20049
rect 24765 20009 24777 20043
rect 24811 20009 24823 20043
rect 24765 20003 24823 20009
rect 23293 19975 23351 19981
rect 23293 19941 23305 19975
rect 23339 19972 23351 19975
rect 23474 19972 23480 19984
rect 23339 19944 23480 19972
rect 23339 19941 23351 19944
rect 23293 19935 23351 19941
rect 23474 19932 23480 19944
rect 23532 19972 23538 19984
rect 24780 19972 24808 20003
rect 25222 20000 25228 20052
rect 25280 20040 25286 20052
rect 25317 20043 25375 20049
rect 25317 20040 25329 20043
rect 25280 20012 25329 20040
rect 25280 20000 25286 20012
rect 25317 20009 25329 20012
rect 25363 20009 25375 20043
rect 25317 20003 25375 20009
rect 23532 19944 24808 19972
rect 23532 19932 23538 19944
rect 23198 19904 23204 19916
rect 22296 19876 23204 19904
rect 23198 19864 23204 19876
rect 23256 19904 23262 19916
rect 23641 19907 23699 19913
rect 23641 19904 23653 19907
rect 23256 19876 23653 19904
rect 23256 19864 23262 19876
rect 23641 19873 23653 19876
rect 23687 19873 23699 19907
rect 23641 19867 23699 19873
rect 14047 19808 15240 19836
rect 15289 19839 15347 19845
rect 14047 19805 14059 19808
rect 14001 19799 14059 19805
rect 15289 19805 15301 19839
rect 15335 19805 15347 19839
rect 15289 19799 15347 19805
rect 13906 19728 13912 19780
rect 13964 19768 13970 19780
rect 14918 19768 14924 19780
rect 13964 19740 14924 19768
rect 13964 19728 13970 19740
rect 14918 19728 14924 19740
rect 14976 19768 14982 19780
rect 15013 19771 15071 19777
rect 15013 19768 15025 19771
rect 14976 19740 15025 19768
rect 14976 19728 14982 19740
rect 15013 19737 15025 19740
rect 15059 19768 15071 19771
rect 15304 19768 15332 19799
rect 17678 19796 17684 19848
rect 17736 19836 17742 19848
rect 18322 19836 18328 19848
rect 17736 19808 18328 19836
rect 17736 19796 17742 19808
rect 18322 19796 18328 19808
rect 18380 19796 18386 19848
rect 19610 19836 19616 19848
rect 19571 19808 19616 19836
rect 19610 19796 19616 19808
rect 19668 19796 19674 19848
rect 23392 19839 23450 19845
rect 23392 19805 23404 19839
rect 23438 19805 23450 19839
rect 23392 19799 23450 19805
rect 15059 19740 15332 19768
rect 15059 19737 15071 19740
rect 15013 19731 15071 19737
rect 23290 19728 23296 19780
rect 23348 19768 23354 19780
rect 23400 19768 23428 19799
rect 23348 19740 23428 19768
rect 23348 19728 23354 19740
rect 11882 19660 11888 19712
rect 11940 19700 11946 19712
rect 11977 19703 12035 19709
rect 11977 19700 11989 19703
rect 11940 19672 11989 19700
rect 11940 19660 11946 19672
rect 11977 19669 11989 19672
rect 12023 19669 12035 19703
rect 12802 19700 12808 19712
rect 12763 19672 12808 19700
rect 11977 19663 12035 19669
rect 12802 19660 12808 19672
rect 12860 19660 12866 19712
rect 13354 19700 13360 19712
rect 13315 19672 13360 19700
rect 13354 19660 13360 19672
rect 13412 19660 13418 19712
rect 14737 19703 14795 19709
rect 14737 19669 14749 19703
rect 14783 19700 14795 19703
rect 14826 19700 14832 19712
rect 14783 19672 14832 19700
rect 14783 19669 14795 19672
rect 14737 19663 14795 19669
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 18690 19660 18696 19712
rect 18748 19700 18754 19712
rect 18785 19703 18843 19709
rect 18785 19700 18797 19703
rect 18748 19672 18797 19700
rect 18748 19660 18754 19672
rect 18785 19669 18797 19672
rect 18831 19669 18843 19703
rect 18785 19663 18843 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 9030 19496 9036 19508
rect 8991 19468 9036 19496
rect 9030 19456 9036 19468
rect 9088 19456 9094 19508
rect 10870 19456 10876 19508
rect 10928 19496 10934 19508
rect 11149 19499 11207 19505
rect 11149 19496 11161 19499
rect 10928 19468 11161 19496
rect 10928 19456 10934 19468
rect 11149 19465 11161 19468
rect 11195 19465 11207 19499
rect 11149 19459 11207 19465
rect 12897 19499 12955 19505
rect 12897 19465 12909 19499
rect 12943 19496 12955 19499
rect 13078 19496 13084 19508
rect 12943 19468 13084 19496
rect 12943 19465 12955 19468
rect 12897 19459 12955 19465
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 14737 19499 14795 19505
rect 14737 19465 14749 19499
rect 14783 19496 14795 19499
rect 15378 19496 15384 19508
rect 14783 19468 15384 19496
rect 14783 19465 14795 19468
rect 14737 19459 14795 19465
rect 15378 19456 15384 19468
rect 15436 19456 15442 19508
rect 15746 19456 15752 19508
rect 15804 19496 15810 19508
rect 16206 19496 16212 19508
rect 15804 19468 16212 19496
rect 15804 19456 15810 19468
rect 16206 19456 16212 19468
rect 16264 19456 16270 19508
rect 16393 19499 16451 19505
rect 16393 19465 16405 19499
rect 16439 19496 16451 19499
rect 16758 19496 16764 19508
rect 16439 19468 16764 19496
rect 16439 19465 16451 19468
rect 16393 19459 16451 19465
rect 16758 19456 16764 19468
rect 16816 19456 16822 19508
rect 17402 19496 17408 19508
rect 17363 19468 17408 19496
rect 17402 19456 17408 19468
rect 17460 19456 17466 19508
rect 20806 19496 20812 19508
rect 20767 19468 20812 19496
rect 20806 19456 20812 19468
rect 20864 19456 20870 19508
rect 21542 19456 21548 19508
rect 21600 19496 21606 19508
rect 21821 19499 21879 19505
rect 21821 19496 21833 19499
rect 21600 19468 21833 19496
rect 21600 19456 21606 19468
rect 21821 19465 21833 19468
rect 21867 19465 21879 19499
rect 21821 19459 21879 19465
rect 23198 19456 23204 19508
rect 23256 19496 23262 19508
rect 23385 19499 23443 19505
rect 23385 19496 23397 19499
rect 23256 19468 23397 19496
rect 23256 19456 23262 19468
rect 23385 19465 23397 19468
rect 23431 19465 23443 19499
rect 23385 19459 23443 19465
rect 24854 19456 24860 19508
rect 24912 19496 24918 19508
rect 25041 19499 25099 19505
rect 25041 19496 25053 19499
rect 24912 19468 25053 19496
rect 24912 19456 24918 19468
rect 25041 19465 25053 19468
rect 25087 19465 25099 19499
rect 25041 19459 25099 19465
rect 9861 19363 9919 19369
rect 9861 19329 9873 19363
rect 9907 19360 9919 19363
rect 10689 19363 10747 19369
rect 10689 19360 10701 19363
rect 9907 19332 10701 19360
rect 9907 19329 9919 19332
rect 9861 19323 9919 19329
rect 10689 19329 10701 19332
rect 10735 19360 10747 19363
rect 10962 19360 10968 19372
rect 10735 19332 10968 19360
rect 10735 19329 10747 19332
rect 10689 19323 10747 19329
rect 10962 19320 10968 19332
rect 11020 19320 11026 19372
rect 15933 19363 15991 19369
rect 15933 19329 15945 19363
rect 15979 19360 15991 19363
rect 17034 19360 17040 19372
rect 15979 19332 17040 19360
rect 15979 19329 15991 19332
rect 15933 19323 15991 19329
rect 17034 19320 17040 19332
rect 17092 19320 17098 19372
rect 17420 19360 17448 19456
rect 18601 19363 18659 19369
rect 18601 19360 18613 19363
rect 17420 19332 18613 19360
rect 18601 19329 18613 19332
rect 18647 19329 18659 19363
rect 18601 19323 18659 19329
rect 21453 19363 21511 19369
rect 21453 19329 21465 19363
rect 21499 19360 21511 19363
rect 21560 19360 21588 19456
rect 22002 19388 22008 19440
rect 22060 19428 22066 19440
rect 23290 19428 23296 19440
rect 22060 19400 23296 19428
rect 22060 19388 22066 19400
rect 23290 19388 23296 19400
rect 23348 19388 23354 19440
rect 21499 19332 21588 19360
rect 21499 19329 21511 19332
rect 21453 19323 21511 19329
rect 21818 19320 21824 19372
rect 21876 19360 21882 19372
rect 22922 19360 22928 19372
rect 21876 19332 22928 19360
rect 21876 19320 21882 19332
rect 22922 19320 22928 19332
rect 22980 19320 22986 19372
rect 7650 19292 7656 19304
rect 7611 19264 7656 19292
rect 7650 19252 7656 19264
rect 7708 19252 7714 19304
rect 12802 19252 12808 19304
rect 12860 19292 12866 19304
rect 13357 19295 13415 19301
rect 13357 19292 13369 19295
rect 12860 19264 13369 19292
rect 12860 19252 12866 19264
rect 13357 19261 13369 19264
rect 13403 19292 13415 19295
rect 13906 19292 13912 19304
rect 13403 19264 13912 19292
rect 13403 19261 13415 19264
rect 13357 19255 13415 19261
rect 13906 19252 13912 19264
rect 13964 19252 13970 19304
rect 17310 19252 17316 19304
rect 17368 19252 17374 19304
rect 17678 19252 17684 19304
rect 17736 19292 17742 19304
rect 17773 19295 17831 19301
rect 17773 19292 17785 19295
rect 17736 19264 17785 19292
rect 17736 19252 17742 19264
rect 17773 19261 17785 19264
rect 17819 19261 17831 19295
rect 18506 19292 18512 19304
rect 18467 19264 18512 19292
rect 17773 19255 17831 19261
rect 18506 19252 18512 19264
rect 18564 19292 18570 19304
rect 19061 19295 19119 19301
rect 19061 19292 19073 19295
rect 18564 19264 19073 19292
rect 18564 19252 18570 19264
rect 19061 19261 19073 19264
rect 19107 19261 19119 19295
rect 19794 19292 19800 19304
rect 19755 19264 19800 19292
rect 19061 19255 19119 19261
rect 19794 19252 19800 19264
rect 19852 19252 19858 19304
rect 20717 19295 20775 19301
rect 20717 19261 20729 19295
rect 20763 19292 20775 19295
rect 20763 19264 21312 19292
rect 20763 19261 20775 19264
rect 20717 19255 20775 19261
rect 7561 19227 7619 19233
rect 7561 19193 7573 19227
rect 7607 19224 7619 19227
rect 7898 19227 7956 19233
rect 7898 19224 7910 19227
rect 7607 19196 7910 19224
rect 7607 19193 7619 19196
rect 7561 19187 7619 19193
rect 7898 19193 7910 19196
rect 7944 19224 7956 19227
rect 9677 19227 9735 19233
rect 7944 19196 8248 19224
rect 7944 19193 7956 19196
rect 7898 19187 7956 19193
rect 8220 19156 8248 19196
rect 9677 19193 9689 19227
rect 9723 19224 9735 19227
rect 10505 19227 10563 19233
rect 9723 19196 10456 19224
rect 9723 19193 9735 19196
rect 9677 19187 9735 19193
rect 9861 19159 9919 19165
rect 9861 19156 9873 19159
rect 8220 19128 9873 19156
rect 9861 19125 9873 19128
rect 9907 19156 9919 19159
rect 9953 19159 10011 19165
rect 9953 19156 9965 19159
rect 9907 19128 9965 19156
rect 9907 19125 9919 19128
rect 9861 19119 9919 19125
rect 9953 19125 9965 19128
rect 9999 19125 10011 19159
rect 10134 19156 10140 19168
rect 10095 19128 10140 19156
rect 9953 19119 10011 19125
rect 10134 19116 10140 19128
rect 10192 19116 10198 19168
rect 10428 19156 10456 19196
rect 10505 19193 10517 19227
rect 10551 19224 10563 19227
rect 10686 19224 10692 19236
rect 10551 19196 10692 19224
rect 10551 19193 10563 19196
rect 10505 19187 10563 19193
rect 10686 19184 10692 19196
rect 10744 19224 10750 19236
rect 13630 19233 13636 19236
rect 11517 19227 11575 19233
rect 11517 19224 11529 19227
rect 10744 19196 11529 19224
rect 10744 19184 10750 19196
rect 11517 19193 11529 19196
rect 11563 19193 11575 19227
rect 11517 19187 11575 19193
rect 13265 19227 13323 19233
rect 13265 19193 13277 19227
rect 13311 19224 13323 19227
rect 13624 19224 13636 19233
rect 13311 19196 13636 19224
rect 13311 19193 13323 19196
rect 13265 19187 13323 19193
rect 13624 19187 13636 19196
rect 13630 19184 13636 19187
rect 13688 19184 13694 19236
rect 16114 19184 16120 19236
rect 16172 19224 16178 19236
rect 16761 19227 16819 19233
rect 16761 19224 16773 19227
rect 16172 19196 16773 19224
rect 16172 19184 16178 19196
rect 16761 19193 16773 19196
rect 16807 19224 16819 19227
rect 17328 19224 17356 19252
rect 18414 19224 18420 19236
rect 16807 19196 17356 19224
rect 18375 19196 18420 19224
rect 16807 19193 16819 19196
rect 16761 19187 16819 19193
rect 18414 19184 18420 19196
rect 18472 19224 18478 19236
rect 19429 19227 19487 19233
rect 19429 19224 19441 19227
rect 18472 19196 19441 19224
rect 18472 19184 18478 19196
rect 19429 19193 19441 19196
rect 19475 19193 19487 19227
rect 19429 19187 19487 19193
rect 20349 19227 20407 19233
rect 20349 19193 20361 19227
rect 20395 19224 20407 19227
rect 20395 19196 20944 19224
rect 20395 19193 20407 19196
rect 20349 19187 20407 19193
rect 20916 19168 20944 19196
rect 10597 19159 10655 19165
rect 10597 19156 10609 19159
rect 10428 19128 10609 19156
rect 10597 19125 10609 19128
rect 10643 19156 10655 19159
rect 10778 19156 10784 19168
rect 10643 19128 10784 19156
rect 10643 19125 10655 19128
rect 10597 19119 10655 19125
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 11977 19159 12035 19165
rect 11977 19125 11989 19159
rect 12023 19156 12035 19159
rect 12158 19156 12164 19168
rect 12023 19128 12164 19156
rect 12023 19125 12035 19128
rect 11977 19119 12035 19125
rect 12158 19116 12164 19128
rect 12216 19116 12222 19168
rect 16301 19159 16359 19165
rect 16301 19125 16313 19159
rect 16347 19156 16359 19159
rect 16390 19156 16396 19168
rect 16347 19128 16396 19156
rect 16347 19125 16359 19128
rect 16301 19119 16359 19125
rect 16390 19116 16396 19128
rect 16448 19156 16454 19168
rect 16853 19159 16911 19165
rect 16853 19156 16865 19159
rect 16448 19128 16865 19156
rect 16448 19116 16454 19128
rect 16853 19125 16865 19128
rect 16899 19125 16911 19159
rect 18046 19156 18052 19168
rect 18007 19128 18052 19156
rect 16853 19119 16911 19125
rect 18046 19116 18052 19128
rect 18104 19116 18110 19168
rect 20898 19116 20904 19168
rect 20956 19156 20962 19168
rect 21284 19165 21312 19264
rect 22186 19252 22192 19304
rect 22244 19292 22250 19304
rect 22465 19295 22523 19301
rect 22465 19292 22477 19295
rect 22244 19264 22477 19292
rect 22244 19252 22250 19264
rect 22465 19261 22477 19264
rect 22511 19292 22523 19295
rect 23017 19295 23075 19301
rect 23017 19292 23029 19295
rect 22511 19264 23029 19292
rect 22511 19261 22523 19264
rect 22465 19255 22523 19261
rect 23017 19261 23029 19264
rect 23063 19292 23075 19295
rect 23198 19292 23204 19304
rect 23063 19264 23204 19292
rect 23063 19261 23075 19264
rect 23017 19255 23075 19261
rect 23198 19252 23204 19264
rect 23256 19252 23262 19304
rect 23290 19252 23296 19304
rect 23348 19292 23354 19304
rect 23661 19295 23719 19301
rect 23661 19292 23673 19295
rect 23348 19264 23673 19292
rect 23348 19252 23354 19264
rect 23661 19261 23673 19264
rect 23707 19292 23719 19295
rect 24946 19292 24952 19304
rect 23707 19264 24952 19292
rect 23707 19261 23719 19264
rect 23661 19255 23719 19261
rect 24946 19252 24952 19264
rect 25004 19252 25010 19304
rect 22554 19224 22560 19236
rect 21836 19196 22560 19224
rect 21836 19168 21864 19196
rect 22554 19184 22560 19196
rect 22612 19184 22618 19236
rect 23474 19184 23480 19236
rect 23532 19224 23538 19236
rect 23906 19227 23964 19233
rect 23906 19224 23918 19227
rect 23532 19196 23918 19224
rect 23532 19184 23538 19196
rect 23906 19193 23918 19196
rect 23952 19193 23964 19227
rect 23906 19187 23964 19193
rect 21177 19159 21235 19165
rect 21177 19156 21189 19159
rect 20956 19128 21189 19156
rect 20956 19116 20962 19128
rect 21177 19125 21189 19128
rect 21223 19125 21235 19159
rect 21177 19119 21235 19125
rect 21269 19159 21327 19165
rect 21269 19125 21281 19159
rect 21315 19156 21327 19159
rect 21818 19156 21824 19168
rect 21315 19128 21824 19156
rect 21315 19125 21327 19128
rect 21269 19119 21327 19125
rect 21818 19116 21824 19128
rect 21876 19116 21882 19168
rect 22002 19116 22008 19168
rect 22060 19156 22066 19168
rect 22189 19159 22247 19165
rect 22189 19156 22201 19159
rect 22060 19128 22201 19156
rect 22060 19116 22066 19128
rect 22189 19125 22201 19128
rect 22235 19125 22247 19159
rect 22646 19156 22652 19168
rect 22607 19128 22652 19156
rect 22189 19119 22247 19125
rect 22646 19116 22652 19128
rect 22704 19116 22710 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 10778 18912 10784 18964
rect 10836 18952 10842 18964
rect 12161 18955 12219 18961
rect 12161 18952 12173 18955
rect 10836 18924 12173 18952
rect 10836 18912 10842 18924
rect 12161 18921 12173 18924
rect 12207 18921 12219 18955
rect 13446 18952 13452 18964
rect 13407 18924 13452 18952
rect 12161 18915 12219 18921
rect 13446 18912 13452 18924
rect 13504 18912 13510 18964
rect 14458 18912 14464 18964
rect 14516 18952 14522 18964
rect 15286 18952 15292 18964
rect 14516 18924 15292 18952
rect 14516 18912 14522 18924
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 15746 18952 15752 18964
rect 15707 18924 15752 18952
rect 15746 18912 15752 18924
rect 15804 18912 15810 18964
rect 16853 18955 16911 18961
rect 16853 18921 16865 18955
rect 16899 18952 16911 18955
rect 18046 18952 18052 18964
rect 16899 18924 18052 18952
rect 16899 18921 16911 18924
rect 16853 18915 16911 18921
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 19889 18955 19947 18961
rect 19889 18952 19901 18955
rect 19392 18924 19901 18952
rect 19392 18912 19398 18924
rect 19889 18921 19901 18924
rect 19935 18921 19947 18955
rect 21634 18952 21640 18964
rect 21595 18924 21640 18952
rect 19889 18915 19947 18921
rect 21634 18912 21640 18924
rect 21692 18912 21698 18964
rect 22738 18952 22744 18964
rect 22699 18924 22744 18952
rect 22738 18912 22744 18924
rect 22796 18912 22802 18964
rect 23474 18952 23480 18964
rect 23435 18924 23480 18952
rect 23474 18912 23480 18924
rect 23532 18912 23538 18964
rect 23658 18952 23664 18964
rect 23619 18924 23664 18952
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 21177 18887 21235 18893
rect 21177 18853 21189 18887
rect 21223 18884 21235 18887
rect 21542 18884 21548 18896
rect 21223 18856 21548 18884
rect 21223 18853 21235 18856
rect 21177 18847 21235 18853
rect 21542 18844 21548 18856
rect 21600 18844 21606 18896
rect 23492 18884 23520 18912
rect 23492 18856 24256 18884
rect 9490 18816 9496 18828
rect 9451 18788 9496 18816
rect 9490 18776 9496 18788
rect 9548 18776 9554 18828
rect 9950 18825 9956 18828
rect 9944 18816 9956 18825
rect 9911 18788 9956 18816
rect 9944 18779 9956 18788
rect 9950 18776 9956 18779
rect 10008 18776 10014 18828
rect 12250 18776 12256 18828
rect 12308 18816 12314 18828
rect 12529 18819 12587 18825
rect 12529 18816 12541 18819
rect 12308 18788 12541 18816
rect 12308 18776 12314 18788
rect 12529 18785 12541 18788
rect 12575 18785 12587 18819
rect 15657 18819 15715 18825
rect 15657 18816 15669 18819
rect 12529 18779 12587 18785
rect 15028 18788 15669 18816
rect 9674 18748 9680 18760
rect 9324 18720 9680 18748
rect 7650 18640 7656 18692
rect 7708 18680 7714 18692
rect 9324 18689 9352 18720
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 12621 18751 12679 18757
rect 12621 18748 12633 18751
rect 11992 18720 12633 18748
rect 7745 18683 7803 18689
rect 7745 18680 7757 18683
rect 7708 18652 7757 18680
rect 7708 18640 7714 18652
rect 7745 18649 7757 18652
rect 7791 18680 7803 18683
rect 9309 18683 9367 18689
rect 9309 18680 9321 18683
rect 7791 18652 9321 18680
rect 7791 18649 7803 18652
rect 7745 18643 7803 18649
rect 9309 18649 9321 18652
rect 9355 18649 9367 18683
rect 9309 18643 9367 18649
rect 10962 18640 10968 18692
rect 11020 18680 11026 18692
rect 11057 18683 11115 18689
rect 11057 18680 11069 18683
rect 11020 18652 11069 18680
rect 11020 18640 11026 18652
rect 11057 18649 11069 18652
rect 11103 18649 11115 18683
rect 11057 18643 11115 18649
rect 11146 18572 11152 18624
rect 11204 18612 11210 18624
rect 11992 18621 12020 18720
rect 12621 18717 12633 18720
rect 12667 18717 12679 18751
rect 12621 18711 12679 18717
rect 12710 18708 12716 18760
rect 12768 18748 12774 18760
rect 14185 18751 14243 18757
rect 12768 18720 12813 18748
rect 12768 18708 12774 18720
rect 14185 18717 14197 18751
rect 14231 18748 14243 18751
rect 14274 18748 14280 18760
rect 14231 18720 14280 18748
rect 14231 18717 14243 18720
rect 14185 18711 14243 18717
rect 14274 18708 14280 18720
rect 14332 18708 14338 18760
rect 11977 18615 12035 18621
rect 11977 18612 11989 18615
rect 11204 18584 11989 18612
rect 11204 18572 11210 18584
rect 11977 18581 11989 18584
rect 12023 18581 12035 18615
rect 13814 18612 13820 18624
rect 13775 18584 13820 18612
rect 11977 18575 12035 18581
rect 13814 18572 13820 18584
rect 13872 18572 13878 18624
rect 13906 18572 13912 18624
rect 13964 18612 13970 18624
rect 14645 18615 14703 18621
rect 14645 18612 14657 18615
rect 13964 18584 14657 18612
rect 13964 18572 13970 18584
rect 14645 18581 14657 18584
rect 14691 18581 14703 18615
rect 14645 18575 14703 18581
rect 14826 18572 14832 18624
rect 14884 18612 14890 18624
rect 15028 18621 15056 18788
rect 15657 18785 15669 18788
rect 15703 18785 15715 18819
rect 15657 18779 15715 18785
rect 16758 18776 16764 18828
rect 16816 18816 16822 18828
rect 17129 18819 17187 18825
rect 17129 18816 17141 18819
rect 16816 18788 17141 18816
rect 16816 18776 16822 18788
rect 17129 18785 17141 18788
rect 17175 18785 17187 18819
rect 17586 18816 17592 18828
rect 17547 18788 17592 18816
rect 17129 18779 17187 18785
rect 17586 18776 17592 18788
rect 17644 18776 17650 18828
rect 18138 18776 18144 18828
rect 18196 18816 18202 18828
rect 19242 18816 19248 18828
rect 18196 18788 19248 18816
rect 18196 18776 18202 18788
rect 19242 18776 19248 18788
rect 19300 18776 19306 18828
rect 19337 18819 19395 18825
rect 19337 18785 19349 18819
rect 19383 18816 19395 18819
rect 19383 18788 20760 18816
rect 19383 18785 19395 18788
rect 19337 18779 19395 18785
rect 15838 18748 15844 18760
rect 15799 18720 15844 18748
rect 15838 18708 15844 18720
rect 15896 18708 15902 18760
rect 17678 18748 17684 18760
rect 17639 18720 17684 18748
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 17865 18751 17923 18757
rect 17865 18717 17877 18751
rect 17911 18748 17923 18751
rect 18782 18748 18788 18760
rect 17911 18720 18460 18748
rect 18695 18720 18788 18748
rect 17911 18717 17923 18720
rect 17865 18711 17923 18717
rect 15286 18680 15292 18692
rect 15247 18652 15292 18680
rect 15286 18640 15292 18652
rect 15344 18640 15350 18692
rect 16666 18640 16672 18692
rect 16724 18680 16730 18692
rect 16945 18683 17003 18689
rect 16945 18680 16957 18683
rect 16724 18652 16957 18680
rect 16724 18640 16730 18652
rect 16945 18649 16957 18652
rect 16991 18680 17003 18683
rect 18230 18680 18236 18692
rect 16991 18652 18236 18680
rect 16991 18649 17003 18652
rect 16945 18643 17003 18649
rect 18230 18640 18236 18652
rect 18288 18640 18294 18692
rect 18432 18624 18460 18720
rect 18782 18708 18788 18720
rect 18840 18748 18846 18760
rect 19518 18748 19524 18760
rect 18840 18720 19524 18748
rect 18840 18708 18846 18720
rect 19518 18708 19524 18720
rect 19576 18708 19582 18760
rect 20732 18748 20760 18788
rect 21082 18776 21088 18828
rect 21140 18816 21146 18828
rect 21453 18819 21511 18825
rect 21453 18816 21465 18819
rect 21140 18788 21465 18816
rect 21140 18776 21146 18788
rect 21453 18785 21465 18788
rect 21499 18785 21511 18819
rect 22554 18816 22560 18828
rect 22515 18788 22560 18816
rect 21453 18779 21511 18785
rect 22554 18776 22560 18788
rect 22612 18816 22618 18828
rect 23109 18819 23167 18825
rect 23109 18816 23121 18819
rect 22612 18788 23121 18816
rect 22612 18776 22618 18788
rect 23109 18785 23121 18788
rect 23155 18785 23167 18819
rect 23109 18779 23167 18785
rect 23290 18776 23296 18828
rect 23348 18816 23354 18828
rect 24029 18819 24087 18825
rect 24029 18816 24041 18819
rect 23348 18788 24041 18816
rect 23348 18776 23354 18788
rect 24029 18785 24041 18788
rect 24075 18785 24087 18819
rect 24029 18779 24087 18785
rect 21174 18748 21180 18760
rect 20732 18720 21180 18748
rect 21174 18708 21180 18720
rect 21232 18708 21238 18760
rect 23474 18708 23480 18760
rect 23532 18748 23538 18760
rect 24228 18757 24256 18856
rect 25222 18816 25228 18828
rect 25183 18788 25228 18816
rect 25222 18776 25228 18788
rect 25280 18776 25286 18828
rect 24121 18751 24179 18757
rect 24121 18748 24133 18751
rect 23532 18720 24133 18748
rect 23532 18708 23538 18720
rect 24121 18717 24133 18720
rect 24167 18717 24179 18751
rect 24121 18711 24179 18717
rect 24213 18751 24271 18757
rect 24213 18717 24225 18751
rect 24259 18717 24271 18751
rect 24213 18711 24271 18717
rect 15013 18615 15071 18621
rect 15013 18612 15025 18615
rect 14884 18584 15025 18612
rect 14884 18572 14890 18584
rect 15013 18581 15025 18584
rect 15059 18581 15071 18615
rect 15013 18575 15071 18581
rect 16114 18572 16120 18624
rect 16172 18612 16178 18624
rect 16393 18615 16451 18621
rect 16393 18612 16405 18615
rect 16172 18584 16405 18612
rect 16172 18572 16178 18584
rect 16393 18581 16405 18584
rect 16439 18581 16451 18615
rect 17218 18612 17224 18624
rect 17179 18584 17224 18612
rect 16393 18575 16451 18581
rect 17218 18572 17224 18584
rect 17276 18572 17282 18624
rect 18414 18612 18420 18624
rect 18375 18584 18420 18612
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 18874 18612 18880 18624
rect 18835 18584 18880 18612
rect 18874 18572 18880 18584
rect 18932 18572 18938 18624
rect 20070 18572 20076 18624
rect 20128 18612 20134 18624
rect 20257 18615 20315 18621
rect 20257 18612 20269 18615
rect 20128 18584 20269 18612
rect 20128 18572 20134 18584
rect 20257 18581 20269 18584
rect 20303 18612 20315 18615
rect 20530 18612 20536 18624
rect 20303 18584 20536 18612
rect 20303 18581 20315 18584
rect 20257 18575 20315 18581
rect 20530 18572 20536 18584
rect 20588 18612 20594 18624
rect 20625 18615 20683 18621
rect 20625 18612 20637 18615
rect 20588 18584 20637 18612
rect 20588 18572 20594 18584
rect 20625 18581 20637 18584
rect 20671 18581 20683 18615
rect 20625 18575 20683 18581
rect 24765 18615 24823 18621
rect 24765 18581 24777 18615
rect 24811 18612 24823 18615
rect 24946 18612 24952 18624
rect 24811 18584 24952 18612
rect 24811 18581 24823 18584
rect 24765 18575 24823 18581
rect 24946 18572 24952 18584
rect 25004 18612 25010 18624
rect 25041 18615 25099 18621
rect 25041 18612 25053 18615
rect 25004 18584 25053 18612
rect 25004 18572 25010 18584
rect 25041 18581 25053 18584
rect 25087 18581 25099 18615
rect 25406 18612 25412 18624
rect 25367 18584 25412 18612
rect 25041 18575 25099 18581
rect 25406 18572 25412 18584
rect 25464 18572 25470 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 10321 18411 10379 18417
rect 10321 18377 10333 18411
rect 10367 18408 10379 18411
rect 10686 18408 10692 18420
rect 10367 18380 10692 18408
rect 10367 18377 10379 18380
rect 10321 18371 10379 18377
rect 10686 18368 10692 18380
rect 10744 18368 10750 18420
rect 11425 18411 11483 18417
rect 11425 18377 11437 18411
rect 11471 18408 11483 18411
rect 11882 18408 11888 18420
rect 11471 18380 11888 18408
rect 11471 18377 11483 18380
rect 11425 18371 11483 18377
rect 9217 18275 9275 18281
rect 9217 18241 9229 18275
rect 9263 18272 9275 18275
rect 9950 18272 9956 18284
rect 9263 18244 9956 18272
rect 9263 18241 9275 18244
rect 9217 18235 9275 18241
rect 9950 18232 9956 18244
rect 10008 18272 10014 18284
rect 10965 18275 11023 18281
rect 10965 18272 10977 18275
rect 10008 18244 10977 18272
rect 10008 18232 10014 18244
rect 10965 18241 10977 18244
rect 11011 18272 11023 18275
rect 11440 18272 11468 18371
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 12250 18408 12256 18420
rect 12211 18380 12256 18408
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 13446 18368 13452 18420
rect 13504 18408 13510 18420
rect 13633 18411 13691 18417
rect 13633 18408 13645 18411
rect 13504 18380 13645 18408
rect 13504 18368 13510 18380
rect 13633 18377 13645 18380
rect 13679 18377 13691 18411
rect 13633 18371 13691 18377
rect 13817 18411 13875 18417
rect 13817 18377 13829 18411
rect 13863 18408 13875 18411
rect 14826 18408 14832 18420
rect 13863 18380 14832 18408
rect 13863 18377 13875 18380
rect 13817 18371 13875 18377
rect 11011 18244 11468 18272
rect 11900 18272 11928 18368
rect 12710 18272 12716 18284
rect 11900 18244 12716 18272
rect 11011 18241 11023 18244
rect 10965 18235 11023 18241
rect 12710 18232 12716 18244
rect 12768 18232 12774 18284
rect 13648 18272 13676 18371
rect 14826 18368 14832 18380
rect 14884 18368 14890 18420
rect 15289 18411 15347 18417
rect 15289 18377 15301 18411
rect 15335 18408 15347 18411
rect 15470 18408 15476 18420
rect 15335 18380 15476 18408
rect 15335 18377 15347 18380
rect 15289 18371 15347 18377
rect 15470 18368 15476 18380
rect 15528 18368 15534 18420
rect 15838 18368 15844 18420
rect 15896 18408 15902 18420
rect 16393 18411 16451 18417
rect 16393 18408 16405 18411
rect 15896 18380 16405 18408
rect 15896 18368 15902 18380
rect 16393 18377 16405 18380
rect 16439 18377 16451 18411
rect 16393 18371 16451 18377
rect 19518 18368 19524 18420
rect 19576 18408 19582 18420
rect 19705 18411 19763 18417
rect 19705 18408 19717 18411
rect 19576 18380 19717 18408
rect 19576 18368 19582 18380
rect 19705 18377 19717 18380
rect 19751 18377 19763 18411
rect 20714 18408 20720 18420
rect 20675 18380 20720 18408
rect 19705 18371 19763 18377
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 22094 18368 22100 18420
rect 22152 18408 22158 18420
rect 22152 18380 22197 18408
rect 22152 18368 22158 18380
rect 25222 18368 25228 18420
rect 25280 18408 25286 18420
rect 25593 18411 25651 18417
rect 25593 18408 25605 18411
rect 25280 18380 25605 18408
rect 25280 18368 25286 18380
rect 25593 18377 25605 18380
rect 25639 18377 25651 18411
rect 25593 18371 25651 18377
rect 13998 18300 14004 18352
rect 14056 18340 14062 18352
rect 14921 18343 14979 18349
rect 14921 18340 14933 18343
rect 14056 18312 14933 18340
rect 14056 18300 14062 18312
rect 14921 18309 14933 18312
rect 14967 18309 14979 18343
rect 14921 18303 14979 18309
rect 14369 18275 14427 18281
rect 14369 18272 14381 18275
rect 13648 18244 14381 18272
rect 14369 18241 14381 18244
rect 14415 18241 14427 18275
rect 14369 18235 14427 18241
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 13357 18207 13415 18213
rect 12492 18176 12537 18204
rect 12492 18164 12498 18176
rect 13357 18173 13369 18207
rect 13403 18204 13415 18207
rect 14277 18207 14335 18213
rect 14277 18204 14289 18207
rect 13403 18176 14289 18204
rect 13403 18173 13415 18176
rect 13357 18167 13415 18173
rect 14277 18173 14289 18176
rect 14323 18204 14335 18207
rect 14458 18204 14464 18216
rect 14323 18176 14464 18204
rect 14323 18173 14335 18176
rect 14277 18167 14335 18173
rect 14458 18164 14464 18176
rect 14516 18164 14522 18216
rect 14936 18204 14964 18303
rect 15488 18272 15516 18368
rect 15841 18275 15899 18281
rect 15841 18272 15853 18275
rect 15488 18244 15853 18272
rect 15841 18241 15853 18244
rect 15887 18241 15899 18275
rect 15841 18235 15899 18241
rect 15933 18275 15991 18281
rect 15933 18241 15945 18275
rect 15979 18241 15991 18275
rect 15933 18235 15991 18241
rect 15749 18207 15807 18213
rect 15749 18204 15761 18207
rect 14936 18176 15761 18204
rect 9309 18139 9367 18145
rect 9309 18105 9321 18139
rect 9355 18136 9367 18139
rect 9861 18139 9919 18145
rect 9861 18136 9873 18139
rect 9355 18108 9873 18136
rect 9355 18105 9367 18108
rect 9309 18099 9367 18105
rect 9861 18105 9873 18108
rect 9907 18136 9919 18139
rect 10689 18139 10747 18145
rect 10689 18136 10701 18139
rect 9907 18108 10701 18136
rect 9907 18105 9919 18108
rect 9861 18099 9919 18105
rect 10689 18105 10701 18108
rect 10735 18105 10747 18139
rect 12710 18136 12716 18148
rect 12671 18108 12716 18136
rect 10689 18099 10747 18105
rect 12710 18096 12716 18108
rect 12768 18096 12774 18148
rect 10229 18071 10287 18077
rect 10229 18037 10241 18071
rect 10275 18068 10287 18071
rect 10781 18071 10839 18077
rect 10781 18068 10793 18071
rect 10275 18040 10793 18068
rect 10275 18037 10287 18040
rect 10229 18031 10287 18037
rect 10781 18037 10793 18040
rect 10827 18068 10839 18071
rect 11330 18068 11336 18080
rect 10827 18040 11336 18068
rect 10827 18037 10839 18040
rect 10781 18031 10839 18037
rect 11330 18028 11336 18040
rect 11388 18068 11394 18080
rect 11514 18068 11520 18080
rect 11388 18040 11520 18068
rect 11388 18028 11394 18040
rect 11514 18028 11520 18040
rect 11572 18028 11578 18080
rect 14182 18068 14188 18080
rect 14143 18040 14188 18068
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 14458 18028 14464 18080
rect 14516 18068 14522 18080
rect 14936 18068 14964 18176
rect 15749 18173 15761 18176
rect 15795 18173 15807 18207
rect 15948 18204 15976 18235
rect 16942 18232 16948 18284
rect 17000 18272 17006 18284
rect 17402 18272 17408 18284
rect 17000 18244 17408 18272
rect 17000 18232 17006 18244
rect 17402 18232 17408 18244
rect 17460 18232 17466 18284
rect 18230 18232 18236 18284
rect 18288 18272 18294 18284
rect 18325 18275 18383 18281
rect 18325 18272 18337 18275
rect 18288 18244 18337 18272
rect 18288 18232 18294 18244
rect 18325 18241 18337 18244
rect 18371 18241 18383 18275
rect 20732 18272 20760 18368
rect 21358 18340 21364 18352
rect 21319 18312 21364 18340
rect 21358 18300 21364 18312
rect 21416 18300 21422 18352
rect 22462 18272 22468 18284
rect 20732 18244 22468 18272
rect 18325 18235 18383 18241
rect 22462 18232 22468 18244
rect 22520 18272 22526 18284
rect 23017 18275 23075 18281
rect 23017 18272 23029 18275
rect 22520 18244 23029 18272
rect 22520 18232 22526 18244
rect 23017 18241 23029 18244
rect 23063 18272 23075 18275
rect 23290 18272 23296 18284
rect 23063 18244 23296 18272
rect 23063 18241 23075 18244
rect 23017 18235 23075 18241
rect 23290 18232 23296 18244
rect 23348 18232 23354 18284
rect 15749 18167 15807 18173
rect 15856 18176 15976 18204
rect 15856 18148 15884 18176
rect 16574 18164 16580 18216
rect 16632 18204 16638 18216
rect 17678 18204 17684 18216
rect 16632 18176 17684 18204
rect 16632 18164 16638 18176
rect 17678 18164 17684 18176
rect 17736 18204 17742 18216
rect 17773 18207 17831 18213
rect 17773 18204 17785 18207
rect 17736 18176 17785 18204
rect 17736 18164 17742 18176
rect 17773 18173 17785 18176
rect 17819 18173 17831 18207
rect 17773 18167 17831 18173
rect 21177 18207 21235 18213
rect 21177 18173 21189 18207
rect 21223 18204 21235 18207
rect 21223 18176 21864 18204
rect 21223 18173 21235 18176
rect 21177 18167 21235 18173
rect 15838 18096 15844 18148
rect 15896 18096 15902 18148
rect 16853 18139 16911 18145
rect 16853 18105 16865 18139
rect 16899 18136 16911 18139
rect 17497 18139 17555 18145
rect 16899 18108 17448 18136
rect 16899 18105 16911 18108
rect 16853 18099 16911 18105
rect 15378 18068 15384 18080
rect 14516 18040 14964 18068
rect 15339 18040 15384 18068
rect 14516 18028 14522 18040
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 16942 18068 16948 18080
rect 16903 18040 16948 18068
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 17420 18068 17448 18108
rect 17497 18105 17509 18139
rect 17543 18136 17555 18139
rect 18414 18136 18420 18148
rect 17543 18108 18420 18136
rect 17543 18105 17555 18108
rect 17497 18099 17555 18105
rect 18414 18096 18420 18108
rect 18472 18136 18478 18148
rect 18592 18139 18650 18145
rect 18592 18136 18604 18139
rect 18472 18108 18604 18136
rect 18472 18096 18478 18108
rect 18592 18105 18604 18108
rect 18638 18136 18650 18139
rect 20349 18139 20407 18145
rect 18638 18108 19288 18136
rect 18638 18105 18650 18108
rect 18592 18099 18650 18105
rect 19260 18080 19288 18108
rect 20349 18105 20361 18139
rect 20395 18136 20407 18139
rect 20990 18136 20996 18148
rect 20395 18108 20996 18136
rect 20395 18105 20407 18108
rect 20349 18099 20407 18105
rect 20990 18096 20996 18108
rect 21048 18136 21054 18148
rect 21048 18108 21220 18136
rect 21048 18096 21054 18108
rect 21192 18080 21220 18108
rect 17678 18068 17684 18080
rect 17420 18040 17684 18068
rect 17678 18028 17684 18040
rect 17736 18028 17742 18080
rect 19242 18028 19248 18080
rect 19300 18028 19306 18080
rect 21082 18068 21088 18080
rect 21043 18040 21088 18068
rect 21082 18028 21088 18040
rect 21140 18028 21146 18080
rect 21174 18028 21180 18080
rect 21232 18028 21238 18080
rect 21836 18077 21864 18176
rect 22094 18164 22100 18216
rect 22152 18204 22158 18216
rect 22281 18207 22339 18213
rect 22281 18204 22293 18207
rect 22152 18176 22293 18204
rect 22152 18164 22158 18176
rect 22281 18173 22293 18176
rect 22327 18173 22339 18207
rect 22281 18167 22339 18173
rect 23661 18207 23719 18213
rect 23661 18173 23673 18207
rect 23707 18173 23719 18207
rect 23661 18167 23719 18173
rect 23928 18207 23986 18213
rect 23928 18173 23940 18207
rect 23974 18204 23986 18207
rect 24486 18204 24492 18216
rect 23974 18176 24492 18204
rect 23974 18173 23986 18176
rect 23928 18167 23986 18173
rect 22557 18139 22615 18145
rect 22557 18105 22569 18139
rect 22603 18136 22615 18139
rect 23290 18136 23296 18148
rect 22603 18108 23296 18136
rect 22603 18105 22615 18108
rect 22557 18099 22615 18105
rect 23290 18096 23296 18108
rect 23348 18096 23354 18148
rect 23676 18136 23704 18167
rect 24486 18164 24492 18176
rect 24544 18204 24550 18216
rect 24854 18204 24860 18216
rect 24544 18176 24860 18204
rect 24544 18164 24550 18176
rect 24854 18164 24860 18176
rect 24912 18164 24918 18216
rect 24946 18136 24952 18148
rect 23676 18108 24952 18136
rect 24946 18096 24952 18108
rect 25004 18096 25010 18148
rect 21821 18071 21879 18077
rect 21821 18037 21833 18071
rect 21867 18068 21879 18071
rect 21910 18068 21916 18080
rect 21867 18040 21916 18068
rect 21867 18037 21879 18040
rect 21821 18031 21879 18037
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 23474 18068 23480 18080
rect 23435 18040 23480 18068
rect 23474 18028 23480 18040
rect 23532 18028 23538 18080
rect 25041 18071 25099 18077
rect 25041 18037 25053 18071
rect 25087 18068 25099 18071
rect 25130 18068 25136 18080
rect 25087 18040 25136 18068
rect 25087 18037 25099 18040
rect 25041 18031 25099 18037
rect 25130 18028 25136 18040
rect 25188 18028 25194 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 9401 17867 9459 17873
rect 9401 17833 9413 17867
rect 9447 17864 9459 17867
rect 9490 17864 9496 17876
rect 9447 17836 9496 17864
rect 9447 17833 9459 17836
rect 9401 17827 9459 17833
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 10413 17867 10471 17873
rect 10413 17833 10425 17867
rect 10459 17864 10471 17867
rect 10962 17864 10968 17876
rect 10459 17836 10968 17864
rect 10459 17833 10471 17836
rect 10413 17827 10471 17833
rect 10962 17824 10968 17836
rect 11020 17824 11026 17876
rect 12066 17864 12072 17876
rect 12027 17836 12072 17864
rect 12066 17824 12072 17836
rect 12124 17824 12130 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 13081 17867 13139 17873
rect 13081 17864 13093 17867
rect 12492 17836 13093 17864
rect 12492 17824 12498 17836
rect 13081 17833 13093 17836
rect 13127 17833 13139 17867
rect 13081 17827 13139 17833
rect 13633 17867 13691 17873
rect 13633 17833 13645 17867
rect 13679 17864 13691 17867
rect 14182 17864 14188 17876
rect 13679 17836 14188 17864
rect 13679 17833 13691 17836
rect 13633 17827 13691 17833
rect 14182 17824 14188 17836
rect 14240 17864 14246 17876
rect 14645 17867 14703 17873
rect 14645 17864 14657 17867
rect 14240 17836 14657 17864
rect 14240 17824 14246 17836
rect 14645 17833 14657 17836
rect 14691 17833 14703 17867
rect 14645 17827 14703 17833
rect 14734 17824 14740 17876
rect 14792 17864 14798 17876
rect 15013 17867 15071 17873
rect 15013 17864 15025 17867
rect 14792 17836 15025 17864
rect 14792 17824 14798 17836
rect 15013 17833 15025 17836
rect 15059 17833 15071 17867
rect 15013 17827 15071 17833
rect 18141 17867 18199 17873
rect 18141 17833 18153 17867
rect 18187 17864 18199 17867
rect 18230 17864 18236 17876
rect 18187 17836 18236 17864
rect 18187 17833 18199 17836
rect 18141 17827 18199 17833
rect 18230 17824 18236 17836
rect 18288 17824 18294 17876
rect 19334 17824 19340 17876
rect 19392 17864 19398 17876
rect 19613 17867 19671 17873
rect 19613 17864 19625 17867
rect 19392 17836 19625 17864
rect 19392 17824 19398 17836
rect 19613 17833 19625 17836
rect 19659 17833 19671 17867
rect 24486 17864 24492 17876
rect 24447 17836 24492 17864
rect 19613 17827 19671 17833
rect 24486 17824 24492 17836
rect 24544 17824 24550 17876
rect 25222 17864 25228 17876
rect 25183 17836 25228 17864
rect 25222 17824 25228 17836
rect 25280 17824 25286 17876
rect 10134 17756 10140 17808
rect 10192 17796 10198 17808
rect 10873 17799 10931 17805
rect 10873 17796 10885 17799
rect 10192 17768 10885 17796
rect 10192 17756 10198 17768
rect 10873 17765 10885 17768
rect 10919 17765 10931 17799
rect 10873 17759 10931 17765
rect 14093 17799 14151 17805
rect 14093 17765 14105 17799
rect 14139 17796 14151 17799
rect 14366 17796 14372 17808
rect 14139 17768 14372 17796
rect 14139 17765 14151 17768
rect 14093 17759 14151 17765
rect 14366 17756 14372 17768
rect 14424 17756 14430 17808
rect 16666 17796 16672 17808
rect 15764 17768 16672 17796
rect 9858 17688 9864 17740
rect 9916 17728 9922 17740
rect 10778 17728 10784 17740
rect 9916 17700 10784 17728
rect 9916 17688 9922 17700
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 11977 17731 12035 17737
rect 11977 17697 11989 17731
rect 12023 17728 12035 17731
rect 12437 17731 12495 17737
rect 12437 17728 12449 17731
rect 12023 17700 12449 17728
rect 12023 17697 12035 17700
rect 11977 17691 12035 17697
rect 12437 17697 12449 17700
rect 12483 17728 12495 17731
rect 12894 17728 12900 17740
rect 12483 17700 12900 17728
rect 12483 17697 12495 17700
rect 12437 17691 12495 17697
rect 12894 17688 12900 17700
rect 12952 17728 12958 17740
rect 13078 17728 13084 17740
rect 12952 17700 13084 17728
rect 12952 17688 12958 17700
rect 13078 17688 13084 17700
rect 13136 17688 13142 17740
rect 14001 17731 14059 17737
rect 14001 17697 14013 17731
rect 14047 17728 14059 17731
rect 14274 17728 14280 17740
rect 14047 17700 14280 17728
rect 14047 17697 14059 17700
rect 14001 17691 14059 17697
rect 14274 17688 14280 17700
rect 14332 17728 14338 17740
rect 14734 17728 14740 17740
rect 14332 17700 14740 17728
rect 14332 17688 14338 17700
rect 14734 17688 14740 17700
rect 14792 17688 14798 17740
rect 15286 17688 15292 17740
rect 15344 17728 15350 17740
rect 15764 17737 15792 17768
rect 16666 17756 16672 17768
rect 16724 17756 16730 17808
rect 18248 17796 18276 17824
rect 20165 17799 20223 17805
rect 20165 17796 20177 17799
rect 18248 17768 20177 17796
rect 20165 17765 20177 17768
rect 20211 17765 20223 17799
rect 20165 17759 20223 17765
rect 15749 17731 15807 17737
rect 15749 17728 15761 17731
rect 15344 17700 15761 17728
rect 15344 17688 15350 17700
rect 15749 17697 15761 17700
rect 15795 17697 15807 17731
rect 15749 17691 15807 17697
rect 15838 17688 15844 17740
rect 15896 17728 15902 17740
rect 16005 17731 16063 17737
rect 16005 17728 16017 17731
rect 15896 17700 16017 17728
rect 15896 17688 15902 17700
rect 16005 17697 16017 17700
rect 16051 17697 16063 17731
rect 16005 17691 16063 17697
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 18322 17728 18328 17740
rect 17184 17700 18328 17728
rect 17184 17688 17190 17700
rect 18322 17688 18328 17700
rect 18380 17728 18386 17740
rect 21174 17737 21180 17740
rect 18489 17731 18547 17737
rect 18489 17728 18501 17731
rect 18380 17700 18501 17728
rect 18380 17688 18386 17700
rect 18489 17697 18501 17700
rect 18535 17697 18547 17731
rect 21168 17728 21180 17737
rect 21135 17700 21180 17728
rect 18489 17691 18547 17697
rect 21168 17691 21180 17700
rect 21174 17688 21180 17691
rect 21232 17688 21238 17740
rect 22646 17688 22652 17740
rect 22704 17728 22710 17740
rect 23845 17731 23903 17737
rect 23845 17728 23857 17731
rect 22704 17700 23857 17728
rect 22704 17688 22710 17700
rect 23845 17697 23857 17700
rect 23891 17728 23903 17731
rect 24854 17728 24860 17740
rect 23891 17700 24860 17728
rect 23891 17697 23903 17700
rect 23845 17691 23903 17697
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 25038 17728 25044 17740
rect 24999 17700 25044 17728
rect 25038 17688 25044 17700
rect 25096 17688 25102 17740
rect 10962 17620 10968 17672
rect 11020 17660 11026 17672
rect 11020 17632 11065 17660
rect 11020 17620 11026 17632
rect 12250 17620 12256 17672
rect 12308 17660 12314 17672
rect 12529 17663 12587 17669
rect 12529 17660 12541 17663
rect 12308 17632 12541 17660
rect 12308 17620 12314 17632
rect 12529 17629 12541 17632
rect 12575 17629 12587 17663
rect 12529 17623 12587 17629
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17660 12771 17663
rect 13630 17660 13636 17672
rect 12759 17632 13636 17660
rect 12759 17629 12771 17632
rect 12713 17623 12771 17629
rect 11609 17595 11667 17601
rect 11609 17561 11621 17595
rect 11655 17592 11667 17595
rect 12728 17592 12756 17623
rect 13630 17620 13636 17632
rect 13688 17660 13694 17672
rect 14185 17663 14243 17669
rect 14185 17660 14197 17663
rect 13688 17632 14197 17660
rect 13688 17620 13694 17632
rect 14185 17629 14197 17632
rect 14231 17660 14243 17663
rect 14826 17660 14832 17672
rect 14231 17632 14832 17660
rect 14231 17629 14243 17632
rect 14185 17623 14243 17629
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 18230 17660 18236 17672
rect 18191 17632 18236 17660
rect 18230 17620 18236 17632
rect 18288 17620 18294 17672
rect 20901 17663 20959 17669
rect 20901 17660 20913 17663
rect 20548 17632 20913 17660
rect 13449 17595 13507 17601
rect 13449 17592 13461 17595
rect 11655 17564 12756 17592
rect 12912 17564 13461 17592
rect 11655 17561 11667 17564
rect 11609 17555 11667 17561
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 9953 17527 10011 17533
rect 9953 17524 9965 17527
rect 9732 17496 9965 17524
rect 9732 17484 9738 17496
rect 9953 17493 9965 17496
rect 9999 17524 10011 17527
rect 10870 17524 10876 17536
rect 9999 17496 10876 17524
rect 9999 17493 10011 17496
rect 9953 17487 10011 17493
rect 10870 17484 10876 17496
rect 10928 17524 10934 17536
rect 12158 17524 12164 17536
rect 10928 17496 12164 17524
rect 10928 17484 10934 17496
rect 12158 17484 12164 17496
rect 12216 17524 12222 17536
rect 12912 17524 12940 17564
rect 13449 17561 13461 17564
rect 13495 17561 13507 17595
rect 13449 17555 13507 17561
rect 16758 17552 16764 17604
rect 16816 17592 16822 17604
rect 17681 17595 17739 17601
rect 17681 17592 17693 17595
rect 16816 17564 17693 17592
rect 16816 17552 16822 17564
rect 17681 17561 17693 17564
rect 17727 17592 17739 17595
rect 17862 17592 17868 17604
rect 17727 17564 17868 17592
rect 17727 17561 17739 17564
rect 17681 17555 17739 17561
rect 17862 17552 17868 17564
rect 17920 17552 17926 17604
rect 12216 17496 12940 17524
rect 15565 17527 15623 17533
rect 12216 17484 12222 17496
rect 15565 17493 15577 17527
rect 15611 17524 15623 17527
rect 15746 17524 15752 17536
rect 15611 17496 15752 17524
rect 15611 17493 15623 17496
rect 15565 17487 15623 17493
rect 15746 17484 15752 17496
rect 15804 17484 15810 17536
rect 16022 17484 16028 17536
rect 16080 17524 16086 17536
rect 16390 17524 16396 17536
rect 16080 17496 16396 17524
rect 16080 17484 16086 17496
rect 16390 17484 16396 17496
rect 16448 17484 16454 17536
rect 17126 17524 17132 17536
rect 17087 17496 17132 17524
rect 17126 17484 17132 17496
rect 17184 17484 17190 17536
rect 20070 17484 20076 17536
rect 20128 17524 20134 17536
rect 20548 17533 20576 17632
rect 20901 17629 20913 17632
rect 20947 17629 20959 17663
rect 20901 17623 20959 17629
rect 23658 17620 23664 17672
rect 23716 17660 23722 17672
rect 23937 17663 23995 17669
rect 23937 17660 23949 17663
rect 23716 17632 23949 17660
rect 23716 17620 23722 17632
rect 23937 17629 23949 17632
rect 23983 17629 23995 17663
rect 23937 17623 23995 17629
rect 24121 17663 24179 17669
rect 24121 17629 24133 17663
rect 24167 17660 24179 17663
rect 24670 17660 24676 17672
rect 24167 17632 24676 17660
rect 24167 17629 24179 17632
rect 24121 17623 24179 17629
rect 24670 17620 24676 17632
rect 24728 17660 24734 17672
rect 25130 17660 25136 17672
rect 24728 17632 25136 17660
rect 24728 17620 24734 17632
rect 25130 17620 25136 17632
rect 25188 17620 25194 17672
rect 23017 17595 23075 17601
rect 23017 17561 23029 17595
rect 23063 17592 23075 17595
rect 23474 17592 23480 17604
rect 23063 17564 23480 17592
rect 23063 17561 23075 17564
rect 23017 17555 23075 17561
rect 23474 17552 23480 17564
rect 23532 17552 23538 17604
rect 20533 17527 20591 17533
rect 20533 17524 20545 17527
rect 20128 17496 20545 17524
rect 20128 17484 20134 17496
rect 20533 17493 20545 17496
rect 20579 17493 20591 17527
rect 22278 17524 22284 17536
rect 22239 17496 22284 17524
rect 20533 17487 20591 17493
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 23382 17524 23388 17536
rect 23343 17496 23388 17524
rect 23382 17484 23388 17496
rect 23440 17484 23446 17536
rect 24946 17524 24952 17536
rect 24907 17496 24952 17524
rect 24946 17484 24952 17496
rect 25004 17484 25010 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 10137 17323 10195 17329
rect 10137 17289 10149 17323
rect 10183 17320 10195 17323
rect 10962 17320 10968 17332
rect 10183 17292 10968 17320
rect 10183 17289 10195 17292
rect 10137 17283 10195 17289
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 12161 17323 12219 17329
rect 12161 17289 12173 17323
rect 12207 17320 12219 17323
rect 12250 17320 12256 17332
rect 12207 17292 12256 17320
rect 12207 17289 12219 17292
rect 12161 17283 12219 17289
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 14734 17320 14740 17332
rect 14695 17292 14740 17320
rect 14734 17280 14740 17292
rect 14792 17280 14798 17332
rect 16025 17323 16083 17329
rect 16025 17289 16037 17323
rect 16071 17320 16083 17323
rect 16482 17320 16488 17332
rect 16071 17292 16488 17320
rect 16071 17289 16083 17292
rect 16025 17283 16083 17289
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 20165 17323 20223 17329
rect 20165 17289 20177 17323
rect 20211 17320 20223 17323
rect 21174 17320 21180 17332
rect 20211 17292 21180 17320
rect 20211 17289 20223 17292
rect 20165 17283 20223 17289
rect 21174 17280 21180 17292
rect 21232 17320 21238 17332
rect 21450 17320 21456 17332
rect 21232 17292 21456 17320
rect 21232 17280 21238 17292
rect 21450 17280 21456 17292
rect 21508 17320 21514 17332
rect 21637 17323 21695 17329
rect 21637 17320 21649 17323
rect 21508 17292 21649 17320
rect 21508 17280 21514 17292
rect 21637 17289 21649 17292
rect 21683 17289 21695 17323
rect 22646 17320 22652 17332
rect 22607 17292 22652 17320
rect 21637 17283 21695 17289
rect 22646 17280 22652 17292
rect 22704 17280 22710 17332
rect 23477 17323 23535 17329
rect 23477 17289 23489 17323
rect 23523 17320 23535 17323
rect 23658 17320 23664 17332
rect 23523 17292 23664 17320
rect 23523 17289 23535 17292
rect 23477 17283 23535 17289
rect 23658 17280 23664 17292
rect 23716 17280 23722 17332
rect 25130 17320 25136 17332
rect 25091 17292 25136 17320
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 10778 17252 10784 17264
rect 10739 17224 10784 17252
rect 10778 17212 10784 17224
rect 10836 17212 10842 17264
rect 17037 17255 17095 17261
rect 17037 17252 17049 17255
rect 16500 17224 17049 17252
rect 10134 17144 10140 17196
rect 10192 17184 10198 17196
rect 10413 17187 10471 17193
rect 10413 17184 10425 17187
rect 10192 17156 10425 17184
rect 10192 17144 10198 17156
rect 10413 17153 10425 17156
rect 10459 17153 10471 17187
rect 11330 17184 11336 17196
rect 11291 17156 11336 17184
rect 10413 17147 10471 17153
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 12158 17144 12164 17196
rect 12216 17184 12222 17196
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12216 17156 12449 17184
rect 12216 17144 12222 17156
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 16500 17193 16528 17224
rect 17037 17221 17049 17224
rect 17083 17221 17095 17255
rect 17037 17215 17095 17221
rect 17862 17212 17868 17264
rect 17920 17252 17926 17264
rect 17920 17224 20300 17252
rect 17920 17212 17926 17224
rect 16485 17187 16543 17193
rect 16485 17184 16497 17187
rect 15436 17156 16497 17184
rect 15436 17144 15442 17156
rect 16485 17153 16497 17156
rect 16531 17153 16543 17187
rect 16485 17147 16543 17153
rect 16577 17187 16635 17193
rect 16577 17153 16589 17187
rect 16623 17184 16635 17187
rect 17126 17184 17132 17196
rect 16623 17156 17132 17184
rect 16623 17153 16635 17156
rect 16577 17147 16635 17153
rect 11054 17116 11060 17128
rect 11015 17088 11060 17116
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 15473 17119 15531 17125
rect 15473 17085 15485 17119
rect 15519 17116 15531 17119
rect 16592 17116 16620 17147
rect 17126 17144 17132 17156
rect 17184 17144 17190 17196
rect 17497 17187 17555 17193
rect 17497 17153 17509 17187
rect 17543 17184 17555 17187
rect 18046 17184 18052 17196
rect 17543 17156 18052 17184
rect 17543 17153 17555 17156
rect 17497 17147 17555 17153
rect 18046 17144 18052 17156
rect 18104 17184 18110 17196
rect 18874 17184 18880 17196
rect 18104 17156 18880 17184
rect 18104 17144 18110 17156
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 20272 17184 20300 17224
rect 20272 17156 20392 17184
rect 15519 17088 16620 17116
rect 15519 17085 15531 17088
rect 15473 17079 15531 17085
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 18230 17116 18236 17128
rect 18012 17088 18236 17116
rect 18012 17076 18018 17088
rect 18230 17076 18236 17088
rect 18288 17116 18294 17128
rect 18598 17116 18604 17128
rect 18288 17088 18604 17116
rect 18288 17076 18294 17088
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 20070 17116 20076 17128
rect 19392 17088 20076 17116
rect 19392 17076 19398 17088
rect 20070 17076 20076 17088
rect 20128 17116 20134 17128
rect 20257 17119 20315 17125
rect 20257 17116 20269 17119
rect 20128 17088 20269 17116
rect 20128 17076 20134 17088
rect 20257 17085 20269 17088
rect 20303 17085 20315 17119
rect 20364 17116 20392 17156
rect 23382 17144 23388 17196
rect 23440 17184 23446 17196
rect 23658 17184 23664 17196
rect 23440 17156 23664 17184
rect 23440 17144 23446 17156
rect 23658 17144 23664 17156
rect 23716 17184 23722 17196
rect 24121 17187 24179 17193
rect 24121 17184 24133 17187
rect 23716 17156 24133 17184
rect 23716 17144 23722 17156
rect 24121 17153 24133 17156
rect 24167 17153 24179 17187
rect 24121 17147 24179 17153
rect 24210 17144 24216 17196
rect 24268 17184 24274 17196
rect 24673 17187 24731 17193
rect 24673 17184 24685 17187
rect 24268 17156 24685 17184
rect 24268 17144 24274 17156
rect 24673 17153 24685 17156
rect 24719 17153 24731 17187
rect 24673 17147 24731 17153
rect 22281 17119 22339 17125
rect 22281 17116 22293 17119
rect 20364 17088 22293 17116
rect 20257 17079 20315 17085
rect 22281 17085 22293 17088
rect 22327 17116 22339 17119
rect 22925 17119 22983 17125
rect 22925 17116 22937 17119
rect 22327 17088 22937 17116
rect 22327 17085 22339 17088
rect 22281 17079 22339 17085
rect 22925 17085 22937 17088
rect 22971 17085 22983 17119
rect 22925 17079 22983 17085
rect 23474 17076 23480 17128
rect 23532 17116 23538 17128
rect 24029 17119 24087 17125
rect 24029 17116 24041 17119
rect 23532 17088 24041 17116
rect 23532 17076 23538 17088
rect 24029 17085 24041 17088
rect 24075 17085 24087 17119
rect 25222 17116 25228 17128
rect 25183 17088 25228 17116
rect 24029 17079 24087 17085
rect 25222 17076 25228 17088
rect 25280 17116 25286 17128
rect 25961 17119 26019 17125
rect 25961 17116 25973 17119
rect 25280 17088 25973 17116
rect 25280 17076 25286 17088
rect 25961 17085 25973 17088
rect 26007 17085 26019 17119
rect 25961 17079 26019 17085
rect 12704 17051 12762 17057
rect 12704 17017 12716 17051
rect 12750 17048 12762 17051
rect 13170 17048 13176 17060
rect 12750 17020 13176 17048
rect 12750 17017 12762 17020
rect 12704 17011 12762 17017
rect 13170 17008 13176 17020
rect 13228 17008 13234 17060
rect 17865 17051 17923 17057
rect 17865 17017 17877 17051
rect 17911 17048 17923 17051
rect 17911 17020 18736 17048
rect 17911 17017 17923 17020
rect 17865 17011 17923 17017
rect 18708 16992 18736 17020
rect 19150 17008 19156 17060
rect 19208 17048 19214 17060
rect 19613 17051 19671 17057
rect 19613 17048 19625 17051
rect 19208 17020 19625 17048
rect 19208 17008 19214 17020
rect 19613 17017 19625 17020
rect 19659 17017 19671 17051
rect 19613 17011 19671 17017
rect 20346 17008 20352 17060
rect 20404 17048 20410 17060
rect 20502 17051 20560 17057
rect 20502 17048 20514 17051
rect 20404 17020 20514 17048
rect 20404 17008 20410 17020
rect 20502 17017 20514 17020
rect 20548 17017 20560 17051
rect 25498 17048 25504 17060
rect 25459 17020 25504 17048
rect 20502 17011 20560 17017
rect 25498 17008 25504 17020
rect 25556 17008 25562 17060
rect 13817 16983 13875 16989
rect 13817 16949 13829 16983
rect 13863 16980 13875 16983
rect 14182 16980 14188 16992
rect 13863 16952 14188 16980
rect 13863 16949 13875 16952
rect 13817 16943 13875 16949
rect 14182 16940 14188 16952
rect 14240 16940 14246 16992
rect 14274 16940 14280 16992
rect 14332 16980 14338 16992
rect 14369 16983 14427 16989
rect 14369 16980 14381 16983
rect 14332 16952 14381 16980
rect 14332 16940 14338 16952
rect 14369 16949 14381 16952
rect 14415 16949 14427 16983
rect 15838 16980 15844 16992
rect 15799 16952 15844 16980
rect 14369 16943 14427 16949
rect 15838 16940 15844 16952
rect 15896 16940 15902 16992
rect 16390 16980 16396 16992
rect 16351 16952 16396 16980
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 18233 16983 18291 16989
rect 18233 16949 18245 16983
rect 18279 16980 18291 16983
rect 18506 16980 18512 16992
rect 18279 16952 18512 16980
rect 18279 16949 18291 16952
rect 18233 16943 18291 16949
rect 18506 16940 18512 16952
rect 18564 16940 18570 16992
rect 18690 16980 18696 16992
rect 18651 16952 18696 16980
rect 18690 16940 18696 16952
rect 18748 16940 18754 16992
rect 19242 16980 19248 16992
rect 19203 16952 19248 16980
rect 19242 16940 19248 16952
rect 19300 16940 19306 16992
rect 22738 16980 22744 16992
rect 22699 16952 22744 16980
rect 22738 16940 22744 16952
rect 22796 16940 22802 16992
rect 23661 16983 23719 16989
rect 23661 16949 23673 16983
rect 23707 16980 23719 16983
rect 23750 16980 23756 16992
rect 23707 16952 23756 16980
rect 23707 16949 23719 16952
rect 23661 16943 23719 16949
rect 23750 16940 23756 16952
rect 23808 16940 23814 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 10505 16779 10563 16785
rect 10505 16745 10517 16779
rect 10551 16776 10563 16779
rect 10778 16776 10784 16788
rect 10551 16748 10784 16776
rect 10551 16745 10563 16748
rect 10505 16739 10563 16745
rect 10778 16736 10784 16748
rect 10836 16776 10842 16788
rect 11054 16776 11060 16788
rect 10836 16748 11060 16776
rect 10836 16736 10842 16748
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 13170 16776 13176 16788
rect 13131 16748 13176 16776
rect 13170 16736 13176 16748
rect 13228 16736 13234 16788
rect 13541 16779 13599 16785
rect 13541 16745 13553 16779
rect 13587 16776 13599 16779
rect 13630 16776 13636 16788
rect 13587 16748 13636 16776
rect 13587 16745 13599 16748
rect 13541 16739 13599 16745
rect 13630 16736 13636 16748
rect 13688 16736 13694 16788
rect 13998 16776 14004 16788
rect 13832 16748 14004 16776
rect 12250 16668 12256 16720
rect 12308 16708 12314 16720
rect 13832 16708 13860 16748
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 15105 16779 15163 16785
rect 15105 16745 15117 16779
rect 15151 16776 15163 16779
rect 15286 16776 15292 16788
rect 15151 16748 15292 16776
rect 15151 16745 15163 16748
rect 15105 16739 15163 16745
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 15657 16779 15715 16785
rect 15657 16745 15669 16779
rect 15703 16776 15715 16779
rect 16390 16776 16396 16788
rect 15703 16748 16396 16776
rect 15703 16745 15715 16748
rect 15657 16739 15715 16745
rect 16390 16736 16396 16748
rect 16448 16776 16454 16788
rect 16669 16779 16727 16785
rect 16669 16776 16681 16779
rect 16448 16748 16681 16776
rect 16448 16736 16454 16748
rect 16669 16745 16681 16748
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 17129 16779 17187 16785
rect 17129 16745 17141 16779
rect 17175 16776 17187 16779
rect 17221 16779 17279 16785
rect 17221 16776 17233 16779
rect 17175 16748 17233 16776
rect 17175 16745 17187 16748
rect 17129 16739 17187 16745
rect 17221 16745 17233 16748
rect 17267 16776 17279 16779
rect 17862 16776 17868 16788
rect 17267 16748 17868 16776
rect 17267 16745 17279 16748
rect 17221 16739 17279 16745
rect 17862 16736 17868 16748
rect 17920 16736 17926 16788
rect 18230 16776 18236 16788
rect 18191 16748 18236 16776
rect 18230 16736 18236 16748
rect 18288 16736 18294 16788
rect 18322 16736 18328 16788
rect 18380 16776 18386 16788
rect 18598 16776 18604 16788
rect 18380 16748 18604 16776
rect 18380 16736 18386 16748
rect 18598 16736 18604 16748
rect 18656 16736 18662 16788
rect 19242 16776 19248 16788
rect 19203 16748 19248 16776
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 20346 16776 20352 16788
rect 20307 16748 20352 16776
rect 20346 16736 20352 16748
rect 20404 16736 20410 16788
rect 20901 16779 20959 16785
rect 20901 16745 20913 16779
rect 20947 16776 20959 16779
rect 22278 16776 22284 16788
rect 20947 16748 22284 16776
rect 20947 16745 20959 16748
rect 20901 16739 20959 16745
rect 22278 16736 22284 16748
rect 22336 16736 22342 16788
rect 22738 16736 22744 16788
rect 22796 16736 22802 16788
rect 24121 16779 24179 16785
rect 24121 16745 24133 16779
rect 24167 16776 24179 16779
rect 24210 16776 24216 16788
rect 24167 16748 24216 16776
rect 24167 16745 24179 16748
rect 24121 16739 24179 16745
rect 24210 16736 24216 16748
rect 24268 16736 24274 16788
rect 25038 16776 25044 16788
rect 24999 16748 25044 16776
rect 25038 16736 25044 16748
rect 25096 16736 25102 16788
rect 25406 16776 25412 16788
rect 25367 16748 25412 16776
rect 25406 16736 25412 16748
rect 25464 16736 25470 16788
rect 14093 16711 14151 16717
rect 14093 16708 14105 16711
rect 12308 16680 13860 16708
rect 13924 16680 14105 16708
rect 12308 16668 12314 16680
rect 10962 16600 10968 16652
rect 11020 16640 11026 16652
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 11020 16612 11161 16640
rect 11020 16600 11026 16612
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 11149 16603 11207 16609
rect 11416 16643 11474 16649
rect 11416 16609 11428 16643
rect 11462 16640 11474 16643
rect 11882 16640 11888 16652
rect 11462 16612 11888 16640
rect 11462 16609 11474 16612
rect 11416 16603 11474 16609
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 13924 16640 13952 16680
rect 14093 16677 14105 16680
rect 14139 16677 14151 16711
rect 14093 16671 14151 16677
rect 16025 16711 16083 16717
rect 16025 16677 16037 16711
rect 16071 16708 16083 16711
rect 16114 16708 16120 16720
rect 16071 16680 16120 16708
rect 16071 16677 16083 16680
rect 16025 16671 16083 16677
rect 16114 16668 16120 16680
rect 16172 16668 16178 16720
rect 16942 16668 16948 16720
rect 17000 16708 17006 16720
rect 17589 16711 17647 16717
rect 17589 16708 17601 16711
rect 17000 16680 17601 16708
rect 17000 16668 17006 16680
rect 17589 16677 17601 16680
rect 17635 16708 17647 16711
rect 17770 16708 17776 16720
rect 17635 16680 17776 16708
rect 17635 16677 17647 16680
rect 17589 16671 17647 16677
rect 17770 16668 17776 16680
rect 17828 16668 17834 16720
rect 18506 16668 18512 16720
rect 18564 16708 18570 16720
rect 19797 16711 19855 16717
rect 19797 16708 19809 16711
rect 18564 16680 19809 16708
rect 18564 16668 18570 16680
rect 19797 16677 19809 16680
rect 19843 16677 19855 16711
rect 19797 16671 19855 16677
rect 21726 16668 21732 16720
rect 21784 16708 21790 16720
rect 22005 16711 22063 16717
rect 22005 16708 22017 16711
rect 21784 16680 22017 16708
rect 21784 16668 21790 16680
rect 22005 16677 22017 16680
rect 22051 16708 22063 16711
rect 22756 16708 22784 16736
rect 24946 16708 24952 16720
rect 22051 16680 24952 16708
rect 22051 16677 22063 16680
rect 22005 16671 22063 16677
rect 13740 16612 13952 16640
rect 13740 16584 13768 16612
rect 13998 16600 14004 16652
rect 14056 16640 14062 16652
rect 15470 16640 15476 16652
rect 14056 16612 14101 16640
rect 15431 16612 15476 16640
rect 14056 16600 14062 16612
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 15838 16600 15844 16652
rect 15896 16640 15902 16652
rect 18046 16640 18052 16652
rect 15896 16612 18052 16640
rect 15896 16600 15902 16612
rect 13262 16532 13268 16584
rect 13320 16572 13326 16584
rect 13722 16572 13728 16584
rect 13320 16544 13728 16572
rect 13320 16532 13326 16544
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 14182 16572 14188 16584
rect 14143 16544 14188 16572
rect 14182 16532 14188 16544
rect 14240 16532 14246 16584
rect 16022 16532 16028 16584
rect 16080 16572 16086 16584
rect 16316 16581 16344 16612
rect 17880 16584 17908 16612
rect 18046 16600 18052 16612
rect 18104 16600 18110 16652
rect 19150 16640 19156 16652
rect 19111 16612 19156 16640
rect 19150 16600 19156 16612
rect 19208 16600 19214 16652
rect 22756 16649 22784 16680
rect 24946 16668 24952 16680
rect 25004 16668 25010 16720
rect 23014 16649 23020 16652
rect 21269 16643 21327 16649
rect 21269 16640 21281 16643
rect 20640 16612 21281 16640
rect 16117 16575 16175 16581
rect 16117 16572 16129 16575
rect 16080 16544 16129 16572
rect 16080 16532 16086 16544
rect 16117 16541 16129 16544
rect 16163 16541 16175 16575
rect 16117 16535 16175 16541
rect 16301 16575 16359 16581
rect 16301 16541 16313 16575
rect 16347 16541 16359 16575
rect 16301 16535 16359 16541
rect 17494 16532 17500 16584
rect 17552 16572 17558 16584
rect 17681 16575 17739 16581
rect 17681 16572 17693 16575
rect 17552 16544 17693 16572
rect 17552 16532 17558 16544
rect 17681 16541 17693 16544
rect 17727 16541 17739 16575
rect 17862 16572 17868 16584
rect 17775 16544 17868 16572
rect 17681 16535 17739 16541
rect 17862 16532 17868 16544
rect 17920 16532 17926 16584
rect 19337 16575 19395 16581
rect 19337 16541 19349 16575
rect 19383 16541 19395 16575
rect 19337 16535 19395 16541
rect 18874 16464 18880 16516
rect 18932 16504 18938 16516
rect 19352 16504 19380 16535
rect 18932 16476 19380 16504
rect 18932 16464 18938 16476
rect 10873 16439 10931 16445
rect 10873 16405 10885 16439
rect 10919 16436 10931 16439
rect 11146 16436 11152 16448
rect 10919 16408 11152 16436
rect 10919 16405 10931 16408
rect 10873 16399 10931 16405
rect 11146 16396 11152 16408
rect 11204 16396 11210 16448
rect 12526 16436 12532 16448
rect 12487 16408 12532 16436
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 13630 16436 13636 16448
rect 13591 16408 13636 16436
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 14458 16396 14464 16448
rect 14516 16436 14522 16448
rect 14645 16439 14703 16445
rect 14645 16436 14657 16439
rect 14516 16408 14657 16436
rect 14516 16396 14522 16408
rect 14645 16405 14657 16408
rect 14691 16405 14703 16439
rect 18782 16436 18788 16448
rect 18743 16408 18788 16436
rect 14645 16399 14703 16405
rect 18782 16396 18788 16408
rect 18840 16396 18846 16448
rect 20530 16396 20536 16448
rect 20588 16436 20594 16448
rect 20640 16445 20668 16612
rect 21269 16609 21281 16612
rect 21315 16609 21327 16643
rect 21269 16603 21327 16609
rect 22741 16643 22799 16649
rect 22741 16609 22753 16643
rect 22787 16609 22799 16643
rect 23008 16640 23020 16649
rect 22975 16612 23020 16640
rect 22741 16603 22799 16609
rect 23008 16603 23020 16612
rect 23014 16600 23020 16603
rect 23072 16600 23078 16652
rect 25225 16643 25283 16649
rect 25225 16609 25237 16643
rect 25271 16640 25283 16643
rect 25498 16640 25504 16652
rect 25271 16612 25504 16640
rect 25271 16609 25283 16612
rect 25225 16603 25283 16609
rect 25498 16600 25504 16612
rect 25556 16640 25562 16652
rect 25958 16640 25964 16652
rect 25556 16612 25964 16640
rect 25556 16600 25562 16612
rect 25958 16600 25964 16612
rect 26016 16600 26022 16652
rect 21358 16572 21364 16584
rect 21319 16544 21364 16572
rect 21358 16532 21364 16544
rect 21416 16532 21422 16584
rect 21450 16532 21456 16584
rect 21508 16572 21514 16584
rect 21508 16544 21553 16572
rect 21508 16532 21514 16544
rect 20625 16439 20683 16445
rect 20625 16436 20637 16439
rect 20588 16408 20637 16436
rect 20588 16396 20594 16408
rect 20625 16405 20637 16408
rect 20671 16405 20683 16439
rect 20625 16399 20683 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 10778 16232 10784 16244
rect 10739 16204 10784 16232
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 11882 16232 11888 16244
rect 11843 16204 11888 16232
rect 11882 16192 11888 16204
rect 11940 16192 11946 16244
rect 13722 16232 13728 16244
rect 13683 16204 13728 16232
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 17494 16232 17500 16244
rect 17455 16204 17500 16232
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 17770 16232 17776 16244
rect 17731 16204 17776 16232
rect 17770 16192 17776 16204
rect 17828 16192 17834 16244
rect 19978 16192 19984 16244
rect 20036 16232 20042 16244
rect 20346 16232 20352 16244
rect 20036 16204 20352 16232
rect 20036 16192 20042 16204
rect 20346 16192 20352 16204
rect 20404 16232 20410 16244
rect 21085 16235 21143 16241
rect 21085 16232 21097 16235
rect 20404 16204 21097 16232
rect 20404 16192 20410 16204
rect 21085 16201 21097 16204
rect 21131 16201 21143 16235
rect 21085 16195 21143 16201
rect 21542 16192 21548 16244
rect 21600 16232 21606 16244
rect 21637 16235 21695 16241
rect 21637 16232 21649 16235
rect 21600 16204 21649 16232
rect 21600 16192 21606 16204
rect 21637 16201 21649 16204
rect 21683 16201 21695 16235
rect 23474 16232 23480 16244
rect 23435 16204 23480 16232
rect 21637 16195 21695 16201
rect 23474 16192 23480 16204
rect 23532 16192 23538 16244
rect 23658 16232 23664 16244
rect 23619 16204 23664 16232
rect 23658 16192 23664 16204
rect 23716 16192 23722 16244
rect 25958 16232 25964 16244
rect 25919 16204 25964 16232
rect 25958 16192 25964 16204
rect 26016 16192 26022 16244
rect 10870 16124 10876 16176
rect 10928 16164 10934 16176
rect 12253 16167 12311 16173
rect 10928 16136 11376 16164
rect 10928 16124 10934 16136
rect 11146 16056 11152 16108
rect 11204 16096 11210 16108
rect 11348 16105 11376 16136
rect 12253 16133 12265 16167
rect 12299 16164 12311 16167
rect 12299 16136 13216 16164
rect 12299 16133 12311 16136
rect 12253 16127 12311 16133
rect 11241 16099 11299 16105
rect 11241 16096 11253 16099
rect 11204 16068 11253 16096
rect 11204 16056 11210 16068
rect 11241 16065 11253 16068
rect 11287 16065 11299 16099
rect 11241 16059 11299 16065
rect 11333 16099 11391 16105
rect 11333 16065 11345 16099
rect 11379 16065 11391 16099
rect 11333 16059 11391 16065
rect 11256 16028 11284 16059
rect 12526 16056 12532 16108
rect 12584 16096 12590 16108
rect 12894 16096 12900 16108
rect 12584 16068 12900 16096
rect 12584 16056 12590 16068
rect 12894 16056 12900 16068
rect 12952 16096 12958 16108
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 12952 16068 13001 16096
rect 12952 16056 12958 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 13078 16028 13084 16040
rect 11256 16000 13084 16028
rect 13078 15988 13084 16000
rect 13136 15988 13142 16040
rect 10321 15963 10379 15969
rect 10321 15929 10333 15963
rect 10367 15960 10379 15963
rect 11149 15963 11207 15969
rect 11149 15960 11161 15963
rect 10367 15932 11161 15960
rect 10367 15929 10379 15932
rect 10321 15923 10379 15929
rect 11149 15929 11161 15932
rect 11195 15960 11207 15963
rect 12897 15963 12955 15969
rect 11195 15932 12480 15960
rect 11195 15929 11207 15932
rect 11149 15923 11207 15929
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 10870 15892 10876 15904
rect 10735 15864 10876 15892
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 12452 15901 12480 15932
rect 12897 15929 12909 15963
rect 12943 15960 12955 15963
rect 13188 15960 13216 16136
rect 17678 16124 17684 16176
rect 17736 16164 17742 16176
rect 18049 16167 18107 16173
rect 18049 16164 18061 16167
rect 17736 16136 18061 16164
rect 17736 16124 17742 16136
rect 18049 16133 18061 16136
rect 18095 16133 18107 16167
rect 18049 16127 18107 16133
rect 16850 16096 16856 16108
rect 16811 16068 16856 16096
rect 16850 16056 16856 16068
rect 16908 16056 16914 16108
rect 18506 16096 18512 16108
rect 18467 16068 18512 16096
rect 18506 16056 18512 16068
rect 18564 16056 18570 16108
rect 18598 16056 18604 16108
rect 18656 16096 18662 16108
rect 19061 16099 19119 16105
rect 19061 16096 19073 16099
rect 18656 16068 19073 16096
rect 18656 16056 18662 16068
rect 19061 16065 19073 16068
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 21910 16056 21916 16108
rect 21968 16096 21974 16108
rect 22465 16099 22523 16105
rect 22465 16096 22477 16099
rect 21968 16068 22477 16096
rect 21968 16056 21974 16068
rect 22465 16065 22477 16068
rect 22511 16065 22523 16099
rect 23492 16096 23520 16192
rect 24121 16099 24179 16105
rect 24121 16096 24133 16099
rect 23492 16068 24133 16096
rect 22465 16059 22523 16065
rect 24121 16065 24133 16068
rect 24167 16065 24179 16099
rect 24121 16059 24179 16065
rect 24305 16099 24363 16105
rect 24305 16065 24317 16099
rect 24351 16096 24363 16099
rect 24670 16096 24676 16108
rect 24351 16068 24676 16096
rect 24351 16065 24363 16068
rect 24305 16059 24363 16065
rect 13814 15988 13820 16040
rect 13872 16028 13878 16040
rect 14458 16037 14464 16040
rect 14185 16031 14243 16037
rect 14185 16028 14197 16031
rect 13872 16000 14197 16028
rect 13872 15988 13878 16000
rect 14185 15997 14197 16000
rect 14231 15997 14243 16031
rect 14452 16028 14464 16037
rect 14419 16000 14464 16028
rect 14185 15991 14243 15997
rect 14452 15991 14464 16000
rect 14458 15988 14464 15991
rect 14516 15988 14522 16040
rect 16114 15988 16120 16040
rect 16172 16028 16178 16040
rect 16485 16031 16543 16037
rect 16485 16028 16497 16031
rect 16172 16000 16497 16028
rect 16172 15988 16178 16000
rect 16485 15997 16497 16000
rect 16531 15997 16543 16031
rect 16666 16028 16672 16040
rect 16627 16000 16672 16028
rect 16485 15991 16543 15997
rect 16666 15988 16672 16000
rect 16724 15988 16730 16040
rect 17954 15988 17960 16040
rect 18012 16028 18018 16040
rect 18417 16031 18475 16037
rect 18417 16028 18429 16031
rect 18012 16000 18429 16028
rect 18012 15988 18018 16000
rect 18417 15997 18429 16000
rect 18463 15997 18475 16031
rect 18417 15991 18475 15997
rect 19334 15988 19340 16040
rect 19392 16028 19398 16040
rect 19705 16031 19763 16037
rect 19705 16028 19717 16031
rect 19392 16000 19717 16028
rect 19392 15988 19398 16000
rect 19705 15997 19717 16000
rect 19751 15997 19763 16031
rect 22278 16028 22284 16040
rect 22239 16000 22284 16028
rect 19705 15991 19763 15997
rect 22278 15988 22284 16000
rect 22336 15988 22342 16040
rect 23014 15988 23020 16040
rect 23072 16028 23078 16040
rect 23109 16031 23167 16037
rect 23109 16028 23121 16031
rect 23072 16000 23121 16028
rect 23072 15988 23078 16000
rect 23109 15997 23121 16000
rect 23155 16028 23167 16031
rect 24320 16028 24348 16059
rect 24670 16056 24676 16068
rect 24728 16056 24734 16108
rect 25406 16096 25412 16108
rect 25367 16068 25412 16096
rect 25406 16056 25412 16068
rect 25464 16056 25470 16108
rect 25225 16031 25283 16037
rect 25225 16028 25237 16031
rect 23155 16000 24348 16028
rect 25056 16000 25237 16028
rect 23155 15997 23167 16000
rect 23109 15991 23167 15997
rect 14090 15960 14096 15972
rect 12943 15932 14096 15960
rect 12943 15929 12955 15932
rect 12897 15923 12955 15929
rect 14090 15920 14096 15932
rect 14148 15920 14154 15972
rect 19950 15963 20008 15969
rect 19950 15929 19962 15963
rect 19996 15929 20008 15963
rect 19950 15923 20008 15929
rect 22189 15963 22247 15969
rect 22189 15929 22201 15963
rect 22235 15960 22247 15963
rect 23032 15960 23060 15988
rect 22235 15932 23060 15960
rect 22235 15929 22247 15932
rect 22189 15923 22247 15929
rect 12437 15895 12495 15901
rect 12437 15861 12449 15895
rect 12483 15861 12495 15895
rect 12437 15855 12495 15861
rect 12710 15852 12716 15904
rect 12768 15892 12774 15904
rect 12805 15895 12863 15901
rect 12805 15892 12817 15895
rect 12768 15864 12817 15892
rect 12768 15852 12774 15864
rect 12805 15861 12817 15864
rect 12851 15861 12863 15895
rect 13998 15892 14004 15904
rect 13959 15864 14004 15892
rect 12805 15855 12863 15861
rect 13998 15852 14004 15864
rect 14056 15852 14062 15904
rect 15562 15892 15568 15904
rect 15523 15864 15568 15892
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 16022 15852 16028 15904
rect 16080 15892 16086 15904
rect 16117 15895 16175 15901
rect 16117 15892 16129 15895
rect 16080 15864 16129 15892
rect 16080 15852 16086 15864
rect 16117 15861 16129 15864
rect 16163 15861 16175 15895
rect 16117 15855 16175 15861
rect 17954 15852 17960 15904
rect 18012 15892 18018 15904
rect 19521 15895 19579 15901
rect 19521 15892 19533 15895
rect 18012 15864 19533 15892
rect 18012 15852 18018 15864
rect 19521 15861 19533 15864
rect 19567 15892 19579 15895
rect 19965 15892 19993 15923
rect 23842 15920 23848 15972
rect 23900 15960 23906 15972
rect 24029 15963 24087 15969
rect 24029 15960 24041 15963
rect 23900 15932 24041 15960
rect 23900 15920 23906 15932
rect 24029 15929 24041 15932
rect 24075 15929 24087 15963
rect 24029 15923 24087 15929
rect 24765 15963 24823 15969
rect 24765 15929 24777 15963
rect 24811 15960 24823 15963
rect 24946 15960 24952 15972
rect 24811 15932 24952 15960
rect 24811 15929 24823 15932
rect 24765 15923 24823 15929
rect 24946 15920 24952 15932
rect 25004 15920 25010 15972
rect 25056 15904 25084 16000
rect 25225 15997 25237 16000
rect 25271 15997 25283 16031
rect 25225 15991 25283 15997
rect 22278 15892 22284 15904
rect 19567 15864 22284 15892
rect 19567 15861 19579 15864
rect 19521 15855 19579 15861
rect 22278 15852 22284 15864
rect 22336 15852 22342 15904
rect 25038 15892 25044 15904
rect 24999 15864 25044 15892
rect 25038 15852 25044 15864
rect 25096 15852 25102 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 12526 15688 12532 15700
rect 10980 15660 12532 15688
rect 10686 15580 10692 15632
rect 10744 15620 10750 15632
rect 10864 15623 10922 15629
rect 10864 15620 10876 15623
rect 10744 15592 10876 15620
rect 10744 15580 10750 15592
rect 10864 15589 10876 15592
rect 10910 15620 10922 15623
rect 10980 15620 11008 15660
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 12621 15691 12679 15697
rect 12621 15657 12633 15691
rect 12667 15688 12679 15691
rect 12710 15688 12716 15700
rect 12667 15660 12716 15688
rect 12667 15657 12679 15660
rect 12621 15651 12679 15657
rect 12710 15648 12716 15660
rect 12768 15648 12774 15700
rect 13078 15688 13084 15700
rect 13039 15660 13084 15688
rect 13078 15648 13084 15660
rect 13136 15648 13142 15700
rect 13354 15648 13360 15700
rect 13412 15688 13418 15700
rect 13541 15691 13599 15697
rect 13541 15688 13553 15691
rect 13412 15660 13553 15688
rect 13412 15648 13418 15660
rect 13541 15657 13553 15660
rect 13587 15688 13599 15691
rect 13630 15688 13636 15700
rect 13587 15660 13636 15688
rect 13587 15657 13599 15660
rect 13541 15651 13599 15657
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 14182 15688 14188 15700
rect 14143 15660 14188 15688
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 14458 15688 14464 15700
rect 14419 15660 14464 15688
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 15749 15691 15807 15697
rect 15749 15657 15761 15691
rect 15795 15688 15807 15691
rect 15838 15688 15844 15700
rect 15795 15660 15844 15688
rect 15795 15657 15807 15660
rect 15749 15651 15807 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 17678 15688 17684 15700
rect 17639 15660 17684 15688
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 18138 15688 18144 15700
rect 18099 15660 18144 15688
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 18785 15691 18843 15697
rect 18785 15657 18797 15691
rect 18831 15688 18843 15691
rect 18874 15688 18880 15700
rect 18831 15660 18880 15688
rect 18831 15657 18843 15660
rect 18785 15651 18843 15657
rect 18874 15648 18880 15660
rect 18932 15648 18938 15700
rect 19245 15691 19303 15697
rect 19245 15657 19257 15691
rect 19291 15688 19303 15691
rect 21177 15691 21235 15697
rect 21177 15688 21189 15691
rect 19291 15660 21189 15688
rect 19291 15657 19303 15660
rect 19245 15651 19303 15657
rect 21177 15657 21189 15660
rect 21223 15688 21235 15691
rect 21358 15688 21364 15700
rect 21223 15660 21364 15688
rect 21223 15657 21235 15660
rect 21177 15651 21235 15657
rect 21358 15648 21364 15660
rect 21416 15648 21422 15700
rect 21726 15648 21732 15700
rect 21784 15648 21790 15700
rect 22278 15648 22284 15700
rect 22336 15688 22342 15700
rect 22833 15691 22891 15697
rect 22833 15688 22845 15691
rect 22336 15660 22845 15688
rect 22336 15648 22342 15660
rect 22833 15657 22845 15660
rect 22879 15657 22891 15691
rect 22833 15651 22891 15657
rect 23753 15691 23811 15697
rect 23753 15657 23765 15691
rect 23799 15688 23811 15691
rect 23842 15688 23848 15700
rect 23799 15660 23848 15688
rect 23799 15657 23811 15660
rect 23753 15651 23811 15657
rect 23842 15648 23848 15660
rect 23900 15648 23906 15700
rect 23937 15691 23995 15697
rect 23937 15657 23949 15691
rect 23983 15688 23995 15691
rect 25038 15688 25044 15700
rect 23983 15660 25044 15688
rect 23983 15657 23995 15660
rect 23937 15651 23995 15657
rect 25038 15648 25044 15660
rect 25096 15648 25102 15700
rect 10910 15592 11008 15620
rect 10910 15589 10922 15592
rect 10864 15583 10922 15589
rect 11054 15580 11060 15632
rect 11112 15620 11118 15632
rect 16022 15620 16028 15632
rect 11112 15592 16028 15620
rect 11112 15580 11118 15592
rect 16022 15580 16028 15592
rect 16080 15620 16086 15632
rect 16666 15620 16672 15632
rect 16080 15592 16672 15620
rect 16080 15580 16086 15592
rect 16666 15580 16672 15592
rect 16724 15580 16730 15632
rect 17313 15623 17371 15629
rect 17313 15589 17325 15623
rect 17359 15620 17371 15623
rect 17862 15620 17868 15632
rect 17359 15592 17868 15620
rect 17359 15589 17371 15592
rect 17313 15583 17371 15589
rect 17862 15580 17868 15592
rect 17920 15580 17926 15632
rect 19613 15623 19671 15629
rect 19613 15589 19625 15623
rect 19659 15620 19671 15623
rect 20714 15620 20720 15632
rect 19659 15592 20576 15620
rect 20675 15592 20720 15620
rect 19659 15589 19671 15592
rect 19613 15583 19671 15589
rect 12894 15552 12900 15564
rect 12855 15524 12900 15552
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 13170 15512 13176 15564
rect 13228 15552 13234 15564
rect 13449 15555 13507 15561
rect 13449 15552 13461 15555
rect 13228 15524 13461 15552
rect 13228 15512 13234 15524
rect 13449 15521 13461 15524
rect 13495 15521 13507 15555
rect 16482 15552 16488 15564
rect 16443 15524 16488 15552
rect 13449 15515 13507 15521
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 17402 15512 17408 15564
rect 17460 15552 17466 15564
rect 18049 15555 18107 15561
rect 18049 15552 18061 15555
rect 17460 15524 18061 15552
rect 17460 15512 17466 15524
rect 18049 15521 18061 15524
rect 18095 15521 18107 15555
rect 18049 15515 18107 15521
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15552 19763 15555
rect 20548 15552 20576 15592
rect 20714 15580 20720 15592
rect 20772 15580 20778 15632
rect 21744 15620 21772 15648
rect 21468 15592 21772 15620
rect 20806 15552 20812 15564
rect 19751 15524 20392 15552
rect 20548 15524 20812 15552
rect 19751 15521 19763 15524
rect 19705 15515 19763 15521
rect 10594 15484 10600 15496
rect 10555 15456 10600 15484
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 12912 15484 12940 15512
rect 13633 15487 13691 15493
rect 13633 15484 13645 15487
rect 12912 15456 13645 15484
rect 13633 15453 13645 15456
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 16298 15444 16304 15496
rect 16356 15484 16362 15496
rect 16577 15487 16635 15493
rect 16577 15484 16589 15487
rect 16356 15456 16589 15484
rect 16356 15444 16362 15456
rect 16577 15453 16589 15456
rect 16623 15453 16635 15487
rect 16758 15484 16764 15496
rect 16719 15456 16764 15484
rect 16577 15447 16635 15453
rect 16758 15444 16764 15456
rect 16816 15444 16822 15496
rect 18233 15487 18291 15493
rect 18233 15453 18245 15487
rect 18279 15453 18291 15487
rect 18233 15447 18291 15453
rect 19153 15487 19211 15493
rect 19153 15453 19165 15487
rect 19199 15484 19211 15487
rect 19889 15487 19947 15493
rect 19889 15484 19901 15487
rect 19199 15456 19901 15484
rect 19199 15453 19211 15456
rect 19153 15447 19211 15453
rect 19889 15453 19901 15456
rect 19935 15484 19947 15487
rect 19978 15484 19984 15496
rect 19935 15456 19984 15484
rect 19935 15453 19947 15456
rect 19889 15447 19947 15453
rect 14366 15376 14372 15428
rect 14424 15416 14430 15428
rect 14829 15419 14887 15425
rect 14829 15416 14841 15419
rect 14424 15388 14841 15416
rect 14424 15376 14430 15388
rect 14829 15385 14841 15388
rect 14875 15385 14887 15419
rect 14829 15379 14887 15385
rect 17954 15376 17960 15428
rect 18012 15416 18018 15428
rect 18248 15416 18276 15447
rect 19978 15444 19984 15456
rect 20036 15444 20042 15496
rect 20364 15493 20392 15524
rect 20806 15512 20812 15524
rect 20864 15512 20870 15564
rect 21468 15561 21496 15592
rect 21726 15561 21732 15564
rect 21453 15555 21511 15561
rect 21453 15521 21465 15555
rect 21499 15521 21511 15555
rect 21720 15552 21732 15561
rect 21687 15524 21732 15552
rect 21453 15515 21511 15521
rect 21720 15515 21732 15524
rect 21726 15512 21732 15515
rect 21784 15512 21790 15564
rect 23842 15512 23848 15564
rect 23900 15552 23906 15564
rect 24305 15555 24363 15561
rect 24305 15552 24317 15555
rect 23900 15524 24317 15552
rect 23900 15512 23906 15524
rect 24305 15521 24317 15524
rect 24351 15521 24363 15555
rect 24305 15515 24363 15521
rect 24397 15555 24455 15561
rect 24397 15521 24409 15555
rect 24443 15552 24455 15555
rect 24670 15552 24676 15564
rect 24443 15524 24676 15552
rect 24443 15521 24455 15524
rect 24397 15515 24455 15521
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15484 20407 15487
rect 20622 15484 20628 15496
rect 20395 15456 20628 15484
rect 20395 15453 20407 15456
rect 20349 15447 20407 15453
rect 20622 15444 20628 15456
rect 20680 15444 20686 15496
rect 23474 15444 23480 15496
rect 23532 15484 23538 15496
rect 24412 15484 24440 15515
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 23532 15456 24440 15484
rect 24489 15487 24547 15493
rect 23532 15444 23538 15456
rect 24489 15453 24501 15487
rect 24535 15453 24547 15487
rect 24489 15447 24547 15453
rect 18012 15388 18276 15416
rect 18012 15376 18018 15388
rect 23750 15376 23756 15428
rect 23808 15416 23814 15428
rect 24504 15416 24532 15447
rect 23808 15388 24532 15416
rect 23808 15376 23814 15388
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 11977 15351 12035 15357
rect 11977 15348 11989 15351
rect 10928 15320 11989 15348
rect 10928 15308 10934 15320
rect 11977 15317 11989 15320
rect 12023 15317 12035 15351
rect 11977 15311 12035 15317
rect 15746 15308 15752 15360
rect 15804 15348 15810 15360
rect 16117 15351 16175 15357
rect 16117 15348 16129 15351
rect 15804 15320 16129 15348
rect 15804 15308 15810 15320
rect 16117 15317 16129 15320
rect 16163 15317 16175 15351
rect 24946 15348 24952 15360
rect 24907 15320 24952 15348
rect 16117 15311 16175 15317
rect 24946 15308 24952 15320
rect 25004 15308 25010 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 10686 15144 10692 15156
rect 10647 15116 10692 15144
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 12253 15147 12311 15153
rect 12253 15113 12265 15147
rect 12299 15144 12311 15147
rect 13354 15144 13360 15156
rect 12299 15116 13360 15144
rect 12299 15113 12311 15116
rect 12253 15107 12311 15113
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 15378 15144 15384 15156
rect 15291 15116 15384 15144
rect 15378 15104 15384 15116
rect 15436 15144 15442 15156
rect 16482 15144 16488 15156
rect 15436 15116 16488 15144
rect 15436 15104 15442 15116
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 19889 15147 19947 15153
rect 19889 15113 19901 15147
rect 19935 15144 19947 15147
rect 20530 15144 20536 15156
rect 19935 15116 20536 15144
rect 19935 15113 19947 15116
rect 19889 15107 19947 15113
rect 20530 15104 20536 15116
rect 20588 15104 20594 15156
rect 23109 15147 23167 15153
rect 23109 15113 23121 15147
rect 23155 15144 23167 15147
rect 23382 15144 23388 15156
rect 23155 15116 23388 15144
rect 23155 15113 23167 15116
rect 23109 15107 23167 15113
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 23750 15104 23756 15156
rect 23808 15144 23814 15156
rect 23845 15147 23903 15153
rect 23845 15144 23857 15147
rect 23808 15116 23857 15144
rect 23808 15104 23814 15116
rect 23845 15113 23857 15116
rect 23891 15144 23903 15147
rect 25409 15147 25467 15153
rect 25409 15144 25421 15147
rect 23891 15116 25421 15144
rect 23891 15113 23903 15116
rect 23845 15107 23903 15113
rect 25409 15113 25421 15116
rect 25455 15113 25467 15147
rect 25409 15107 25467 15113
rect 11606 15036 11612 15088
rect 11664 15076 11670 15088
rect 11885 15079 11943 15085
rect 11885 15076 11897 15079
rect 11664 15048 11897 15076
rect 11664 15036 11670 15048
rect 11885 15045 11897 15048
rect 11931 15076 11943 15079
rect 13538 15076 13544 15088
rect 11931 15048 13544 15076
rect 11931 15045 11943 15048
rect 11885 15039 11943 15045
rect 13538 15036 13544 15048
rect 13596 15036 13602 15088
rect 16853 15079 16911 15085
rect 16853 15045 16865 15079
rect 16899 15045 16911 15079
rect 16853 15039 16911 15045
rect 12437 15011 12495 15017
rect 12437 14977 12449 15011
rect 12483 15008 12495 15011
rect 12710 15008 12716 15020
rect 12483 14980 12716 15008
rect 12483 14977 12495 14980
rect 12437 14971 12495 14977
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 14366 15008 14372 15020
rect 14327 14980 14372 15008
rect 14366 14968 14372 14980
rect 14424 14968 14430 15020
rect 14458 14968 14464 15020
rect 14516 15008 14522 15020
rect 14516 14980 14561 15008
rect 14516 14968 14522 14980
rect 15286 14968 15292 15020
rect 15344 15008 15350 15020
rect 15473 15011 15531 15017
rect 15473 15008 15485 15011
rect 15344 14980 15485 15008
rect 15344 14968 15350 14980
rect 15473 14977 15485 14980
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 12618 14900 12624 14952
rect 12676 14940 12682 14952
rect 14921 14943 14979 14949
rect 14921 14940 14933 14943
rect 12676 14912 14933 14940
rect 12676 14900 12682 14912
rect 14921 14909 14933 14912
rect 14967 14909 14979 14943
rect 15488 14940 15516 14971
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 16868 15008 16896 15039
rect 19978 15036 19984 15088
rect 20036 15076 20042 15088
rect 20036 15048 20484 15076
rect 20036 15036 20042 15048
rect 18598 15008 18604 15020
rect 16816 14980 18604 15008
rect 16816 14968 16822 14980
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 20346 15008 20352 15020
rect 20307 14980 20352 15008
rect 20346 14968 20352 14980
rect 20404 14968 20410 15020
rect 20456 15017 20484 15048
rect 20806 15036 20812 15088
rect 20864 15076 20870 15088
rect 21453 15079 21511 15085
rect 21453 15076 21465 15079
rect 20864 15048 21465 15076
rect 20864 15036 20870 15048
rect 21453 15045 21465 15048
rect 21499 15045 21511 15079
rect 21453 15039 21511 15045
rect 20441 15011 20499 15017
rect 20441 14977 20453 15011
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 15008 22155 15011
rect 22278 15008 22284 15020
rect 22143 14980 22284 15008
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 22278 14968 22284 14980
rect 22336 15008 22342 15020
rect 22557 15011 22615 15017
rect 22557 15008 22569 15011
rect 22336 14980 22569 15008
rect 22336 14968 22342 14980
rect 22557 14977 22569 14980
rect 22603 14977 22615 15011
rect 23934 15008 23940 15020
rect 22557 14971 22615 14977
rect 23676 14980 23940 15008
rect 23676 14952 23704 14980
rect 23934 14968 23940 14980
rect 23992 14968 23998 15020
rect 16942 14940 16948 14952
rect 15488 14912 16948 14940
rect 14921 14903 14979 14909
rect 10594 14832 10600 14884
rect 10652 14832 10658 14884
rect 11333 14875 11391 14881
rect 11333 14841 11345 14875
rect 11379 14872 11391 14875
rect 13817 14875 13875 14881
rect 13817 14872 13829 14875
rect 11379 14844 13829 14872
rect 11379 14841 11391 14844
rect 11333 14835 11391 14841
rect 13817 14841 13829 14844
rect 13863 14872 13875 14875
rect 14277 14875 14335 14881
rect 14277 14872 14289 14875
rect 13863 14844 14289 14872
rect 13863 14841 13875 14844
rect 13817 14835 13875 14841
rect 14277 14841 14289 14844
rect 14323 14841 14335 14875
rect 14936 14872 14964 14903
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 19521 14943 19579 14949
rect 19521 14909 19533 14943
rect 19567 14940 19579 14943
rect 22462 14940 22468 14952
rect 19567 14912 22468 14940
rect 19567 14909 19579 14912
rect 19521 14903 19579 14909
rect 22462 14900 22468 14912
rect 22520 14940 22526 14952
rect 23014 14940 23020 14952
rect 22520 14912 23020 14940
rect 22520 14900 22526 14912
rect 23014 14900 23020 14912
rect 23072 14900 23078 14952
rect 23658 14900 23664 14952
rect 23716 14900 23722 14952
rect 24029 14943 24087 14949
rect 24029 14909 24041 14943
rect 24075 14940 24087 14943
rect 24075 14912 24992 14940
rect 24075 14909 24087 14912
rect 24029 14903 24087 14909
rect 24964 14884 24992 14912
rect 15562 14872 15568 14884
rect 14936 14844 15568 14872
rect 14277 14835 14335 14841
rect 15562 14832 15568 14844
rect 15620 14872 15626 14884
rect 15718 14875 15776 14881
rect 15718 14872 15730 14875
rect 15620 14844 15730 14872
rect 15620 14832 15626 14844
rect 15718 14841 15730 14844
rect 15764 14841 15776 14875
rect 18414 14872 18420 14884
rect 15718 14835 15776 14841
rect 17788 14844 18420 14872
rect 9858 14764 9864 14816
rect 9916 14804 9922 14816
rect 10229 14807 10287 14813
rect 10229 14804 10241 14807
rect 9916 14776 10241 14804
rect 9916 14764 9922 14776
rect 10229 14773 10241 14776
rect 10275 14804 10287 14807
rect 10612 14804 10640 14832
rect 17788 14816 17816 14844
rect 18414 14832 18420 14844
rect 18472 14832 18478 14884
rect 20990 14872 20996 14884
rect 20903 14844 20996 14872
rect 20990 14832 20996 14844
rect 21048 14872 21054 14884
rect 21174 14872 21180 14884
rect 21048 14844 21180 14872
rect 21048 14832 21054 14844
rect 21174 14832 21180 14844
rect 21232 14872 21238 14884
rect 21821 14875 21879 14881
rect 21821 14872 21833 14875
rect 21232 14844 21833 14872
rect 21232 14832 21238 14844
rect 21821 14841 21833 14844
rect 21867 14841 21879 14875
rect 21821 14835 21879 14841
rect 23106 14832 23112 14884
rect 23164 14872 23170 14884
rect 23477 14875 23535 14881
rect 23477 14872 23489 14875
rect 23164 14844 23489 14872
rect 23164 14832 23170 14844
rect 23477 14841 23489 14844
rect 23523 14872 23535 14875
rect 24296 14875 24354 14881
rect 24296 14872 24308 14875
rect 23523 14844 24308 14872
rect 23523 14841 23535 14844
rect 23477 14835 23535 14841
rect 24296 14841 24308 14844
rect 24342 14872 24354 14875
rect 24486 14872 24492 14884
rect 24342 14844 24492 14872
rect 24342 14841 24354 14844
rect 24296 14835 24354 14841
rect 24486 14832 24492 14844
rect 24544 14832 24550 14884
rect 24946 14832 24952 14884
rect 25004 14832 25010 14884
rect 10962 14804 10968 14816
rect 10275 14776 10968 14804
rect 10275 14773 10287 14776
rect 10229 14767 10287 14773
rect 10962 14764 10968 14776
rect 11020 14804 11026 14816
rect 11149 14807 11207 14813
rect 11149 14804 11161 14807
rect 11020 14776 11161 14804
rect 11020 14764 11026 14776
rect 11149 14773 11161 14776
rect 11195 14773 11207 14807
rect 13170 14804 13176 14816
rect 13131 14776 13176 14804
rect 11149 14767 11207 14773
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 13906 14804 13912 14816
rect 13867 14776 13912 14804
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 17402 14804 17408 14816
rect 17363 14776 17408 14804
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 17770 14804 17776 14816
rect 17731 14776 17776 14804
rect 17770 14764 17776 14776
rect 17828 14764 17834 14816
rect 18046 14804 18052 14816
rect 18007 14776 18052 14804
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 18506 14804 18512 14816
rect 18467 14776 18512 14804
rect 18506 14764 18512 14776
rect 18564 14804 18570 14816
rect 19061 14807 19119 14813
rect 19061 14804 19073 14807
rect 18564 14776 19073 14804
rect 18564 14764 18570 14776
rect 19061 14773 19073 14776
rect 19107 14773 19119 14807
rect 19061 14767 19119 14773
rect 20257 14807 20315 14813
rect 20257 14773 20269 14807
rect 20303 14804 20315 14807
rect 20622 14804 20628 14816
rect 20303 14776 20628 14804
rect 20303 14773 20315 14776
rect 20257 14767 20315 14773
rect 20622 14764 20628 14776
rect 20680 14764 20686 14816
rect 21266 14804 21272 14816
rect 21227 14776 21272 14804
rect 21266 14764 21272 14776
rect 21324 14804 21330 14816
rect 21913 14807 21971 14813
rect 21913 14804 21925 14807
rect 21324 14776 21925 14804
rect 21324 14764 21330 14776
rect 21913 14773 21925 14776
rect 21959 14773 21971 14807
rect 21913 14767 21971 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 10597 14603 10655 14609
rect 10597 14600 10609 14603
rect 9824 14572 10609 14600
rect 9824 14560 9830 14572
rect 10597 14569 10609 14572
rect 10643 14600 10655 14603
rect 10962 14600 10968 14612
rect 10643 14572 10968 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 11606 14600 11612 14612
rect 11567 14572 11612 14600
rect 11606 14560 11612 14572
rect 11664 14560 11670 14612
rect 11977 14603 12035 14609
rect 11977 14569 11989 14603
rect 12023 14600 12035 14603
rect 12437 14603 12495 14609
rect 12437 14600 12449 14603
rect 12023 14572 12449 14600
rect 12023 14569 12035 14572
rect 11977 14563 12035 14569
rect 12437 14569 12449 14572
rect 12483 14600 12495 14603
rect 13906 14600 13912 14612
rect 12483 14572 13912 14600
rect 12483 14569 12495 14572
rect 12437 14563 12495 14569
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 14093 14603 14151 14609
rect 14093 14569 14105 14603
rect 14139 14600 14151 14603
rect 14182 14600 14188 14612
rect 14139 14572 14188 14600
rect 14139 14569 14151 14572
rect 14093 14563 14151 14569
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 15289 14603 15347 14609
rect 15289 14569 15301 14603
rect 15335 14569 15347 14603
rect 15289 14563 15347 14569
rect 12342 14492 12348 14544
rect 12400 14532 12406 14544
rect 12529 14535 12587 14541
rect 12529 14532 12541 14535
rect 12400 14504 12541 14532
rect 12400 14492 12406 14504
rect 12529 14501 12541 14504
rect 12575 14532 12587 14535
rect 15304 14532 15332 14563
rect 15562 14560 15568 14612
rect 15620 14600 15626 14612
rect 15838 14600 15844 14612
rect 15620 14572 15844 14600
rect 15620 14560 15626 14572
rect 15838 14560 15844 14572
rect 15896 14560 15902 14612
rect 16758 14600 16764 14612
rect 16719 14572 16764 14600
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 16942 14560 16948 14612
rect 17000 14600 17006 14612
rect 17037 14603 17095 14609
rect 17037 14600 17049 14603
rect 17000 14572 17049 14600
rect 17000 14560 17006 14572
rect 17037 14569 17049 14572
rect 17083 14569 17095 14603
rect 17037 14563 17095 14569
rect 17681 14603 17739 14609
rect 17681 14569 17693 14603
rect 17727 14600 17739 14603
rect 17862 14600 17868 14612
rect 17727 14572 17868 14600
rect 17727 14569 17739 14572
rect 17681 14563 17739 14569
rect 12575 14504 15332 14532
rect 12575 14501 12587 14504
rect 12529 14495 12587 14501
rect 10778 14464 10784 14476
rect 10739 14436 10784 14464
rect 10778 14424 10784 14436
rect 10836 14464 10842 14476
rect 11606 14464 11612 14476
rect 10836 14436 11612 14464
rect 10836 14424 10842 14436
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 12894 14424 12900 14476
rect 12952 14464 12958 14476
rect 13081 14467 13139 14473
rect 13081 14464 13093 14467
rect 12952 14436 13093 14464
rect 12952 14424 12958 14436
rect 13081 14433 13093 14436
rect 13127 14433 13139 14467
rect 13081 14427 13139 14433
rect 13354 14424 13360 14476
rect 13412 14464 13418 14476
rect 13814 14464 13820 14476
rect 13412 14436 13820 14464
rect 13412 14424 13418 14436
rect 13814 14424 13820 14436
rect 13872 14464 13878 14476
rect 14001 14467 14059 14473
rect 14001 14464 14013 14467
rect 13872 14436 14013 14464
rect 13872 14424 13878 14436
rect 14001 14433 14013 14436
rect 14047 14433 14059 14467
rect 15657 14467 15715 14473
rect 15657 14464 15669 14467
rect 14001 14427 14059 14433
rect 14660 14436 15669 14464
rect 11054 14396 11060 14408
rect 11015 14368 11060 14396
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 12618 14396 12624 14408
rect 12579 14368 12624 14396
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 13906 14396 13912 14408
rect 13587 14368 13912 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 13906 14356 13912 14368
rect 13964 14396 13970 14408
rect 14185 14399 14243 14405
rect 14185 14396 14197 14399
rect 13964 14368 14197 14396
rect 13964 14356 13970 14368
rect 14185 14365 14197 14368
rect 14231 14365 14243 14399
rect 14185 14359 14243 14365
rect 12066 14328 12072 14340
rect 12027 14300 12072 14328
rect 12066 14288 12072 14300
rect 12124 14288 12130 14340
rect 13633 14331 13691 14337
rect 13633 14297 13645 14331
rect 13679 14328 13691 14331
rect 14366 14328 14372 14340
rect 13679 14300 14372 14328
rect 13679 14297 13691 14300
rect 13633 14291 13691 14297
rect 14366 14288 14372 14300
rect 14424 14288 14430 14340
rect 13814 14220 13820 14272
rect 13872 14260 13878 14272
rect 14660 14269 14688 14436
rect 15657 14433 15669 14436
rect 15703 14433 15715 14467
rect 15657 14427 15715 14433
rect 15749 14467 15807 14473
rect 15749 14433 15761 14467
rect 15795 14464 15807 14467
rect 17052 14464 17080 14563
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 18874 14560 18880 14612
rect 18932 14600 18938 14612
rect 19153 14603 19211 14609
rect 19153 14600 19165 14603
rect 18932 14572 19165 14600
rect 18932 14560 18938 14572
rect 19153 14569 19165 14572
rect 19199 14569 19211 14603
rect 19153 14563 19211 14569
rect 19978 14560 19984 14612
rect 20036 14600 20042 14612
rect 20257 14603 20315 14609
rect 20257 14600 20269 14603
rect 20036 14572 20269 14600
rect 20036 14560 20042 14572
rect 20257 14569 20269 14572
rect 20303 14569 20315 14603
rect 20257 14563 20315 14569
rect 20714 14560 20720 14612
rect 20772 14600 20778 14612
rect 20901 14603 20959 14609
rect 20901 14600 20913 14603
rect 20772 14572 20913 14600
rect 20772 14560 20778 14572
rect 20901 14569 20913 14572
rect 20947 14569 20959 14603
rect 20901 14563 20959 14569
rect 21726 14560 21732 14612
rect 21784 14600 21790 14612
rect 21913 14603 21971 14609
rect 21913 14600 21925 14603
rect 21784 14572 21925 14600
rect 21784 14560 21790 14572
rect 21913 14569 21925 14572
rect 21959 14569 21971 14603
rect 21913 14563 21971 14569
rect 23753 14603 23811 14609
rect 23753 14569 23765 14603
rect 23799 14600 23811 14603
rect 23842 14600 23848 14612
rect 23799 14572 23848 14600
rect 23799 14569 23811 14572
rect 23753 14563 23811 14569
rect 23842 14560 23848 14572
rect 23900 14560 23906 14612
rect 24854 14560 24860 14612
rect 24912 14600 24918 14612
rect 25409 14603 25467 14609
rect 25409 14600 25421 14603
rect 24912 14572 25421 14600
rect 24912 14560 24918 14572
rect 25409 14569 25421 14572
rect 25455 14569 25467 14603
rect 25409 14563 25467 14569
rect 18040 14535 18098 14541
rect 18040 14501 18052 14535
rect 18086 14532 18098 14535
rect 18230 14532 18236 14544
rect 18086 14504 18236 14532
rect 18086 14501 18098 14504
rect 18040 14495 18098 14501
rect 18230 14492 18236 14504
rect 18288 14492 18294 14544
rect 20806 14532 20812 14544
rect 20732 14504 20812 14532
rect 17773 14467 17831 14473
rect 17773 14464 17785 14467
rect 15795 14436 15976 14464
rect 17052 14436 17785 14464
rect 15795 14433 15807 14436
rect 15749 14427 15807 14433
rect 15838 14396 15844 14408
rect 15799 14368 15844 14396
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 15105 14331 15163 14337
rect 15105 14297 15117 14331
rect 15151 14328 15163 14331
rect 15286 14328 15292 14340
rect 15151 14300 15292 14328
rect 15151 14297 15163 14300
rect 15105 14291 15163 14297
rect 15286 14288 15292 14300
rect 15344 14328 15350 14340
rect 15948 14328 15976 14436
rect 17773 14433 17785 14436
rect 17819 14464 17831 14467
rect 17862 14464 17868 14476
rect 17819 14436 17868 14464
rect 17819 14433 17831 14436
rect 17773 14427 17831 14433
rect 17862 14424 17868 14436
rect 17920 14424 17926 14476
rect 20732 14473 20760 14504
rect 20806 14492 20812 14504
rect 20864 14492 20870 14544
rect 21269 14535 21327 14541
rect 21269 14501 21281 14535
rect 21315 14532 21327 14535
rect 21358 14532 21364 14544
rect 21315 14504 21364 14532
rect 21315 14501 21327 14504
rect 21269 14495 21327 14501
rect 21358 14492 21364 14504
rect 21416 14492 21422 14544
rect 22370 14492 22376 14544
rect 22428 14532 22434 14544
rect 22741 14535 22799 14541
rect 22741 14532 22753 14535
rect 22428 14504 22753 14532
rect 22428 14492 22434 14504
rect 22741 14501 22753 14504
rect 22787 14501 22799 14535
rect 24946 14532 24952 14544
rect 24907 14504 24952 14532
rect 22741 14495 22799 14501
rect 24946 14492 24952 14504
rect 25004 14492 25010 14544
rect 20717 14467 20775 14473
rect 20717 14433 20729 14467
rect 20763 14433 20775 14467
rect 20717 14427 20775 14433
rect 21818 14424 21824 14476
rect 21876 14464 21882 14476
rect 22465 14467 22523 14473
rect 22465 14464 22477 14467
rect 21876 14436 22477 14464
rect 21876 14424 21882 14436
rect 22465 14433 22477 14436
rect 22511 14464 22523 14467
rect 23201 14467 23259 14473
rect 23201 14464 23213 14467
rect 22511 14436 23213 14464
rect 22511 14433 22523 14436
rect 22465 14427 22523 14433
rect 23201 14433 23213 14436
rect 23247 14433 23259 14467
rect 23201 14427 23259 14433
rect 24026 14424 24032 14476
rect 24084 14464 24090 14476
rect 24213 14467 24271 14473
rect 24213 14464 24225 14467
rect 24084 14436 24225 14464
rect 24084 14424 24090 14436
rect 24213 14433 24225 14436
rect 24259 14433 24271 14467
rect 24213 14427 24271 14433
rect 17310 14356 17316 14408
rect 17368 14396 17374 14408
rect 17678 14396 17684 14408
rect 17368 14368 17684 14396
rect 17368 14356 17374 14368
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 19981 14399 20039 14405
rect 19981 14365 19993 14399
rect 20027 14396 20039 14399
rect 20622 14396 20628 14408
rect 20027 14368 20628 14396
rect 20027 14365 20039 14368
rect 19981 14359 20039 14365
rect 20622 14356 20628 14368
rect 20680 14356 20686 14408
rect 20806 14356 20812 14408
rect 20864 14396 20870 14408
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 20864 14368 21373 14396
rect 20864 14356 20870 14368
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 21545 14399 21603 14405
rect 21545 14365 21557 14399
rect 21591 14396 21603 14399
rect 21634 14396 21640 14408
rect 21591 14368 21640 14396
rect 21591 14365 21603 14368
rect 21545 14359 21603 14365
rect 21634 14356 21640 14368
rect 21692 14396 21698 14408
rect 22278 14396 22284 14408
rect 21692 14368 22284 14396
rect 21692 14356 21698 14368
rect 22278 14356 22284 14368
rect 22336 14356 22342 14408
rect 23842 14356 23848 14408
rect 23900 14396 23906 14408
rect 24305 14399 24363 14405
rect 24305 14396 24317 14399
rect 23900 14368 24317 14396
rect 23900 14356 23906 14368
rect 24305 14365 24317 14368
rect 24351 14365 24363 14399
rect 24486 14396 24492 14408
rect 24399 14368 24492 14396
rect 24305 14359 24363 14365
rect 24486 14356 24492 14368
rect 24544 14356 24550 14408
rect 15344 14300 15976 14328
rect 15344 14288 15350 14300
rect 23198 14288 23204 14340
rect 23256 14328 23262 14340
rect 23860 14328 23888 14356
rect 23256 14300 23888 14328
rect 24504 14328 24532 14356
rect 25498 14328 25504 14340
rect 24504 14300 25504 14328
rect 23256 14288 23262 14300
rect 25498 14288 25504 14300
rect 25556 14288 25562 14340
rect 14645 14263 14703 14269
rect 14645 14260 14657 14263
rect 13872 14232 14657 14260
rect 13872 14220 13878 14232
rect 14645 14229 14657 14232
rect 14691 14229 14703 14263
rect 16298 14260 16304 14272
rect 16259 14232 16304 14260
rect 14645 14223 14703 14229
rect 16298 14220 16304 14232
rect 16356 14220 16362 14272
rect 22278 14260 22284 14272
rect 22239 14232 22284 14260
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 10597 14059 10655 14065
rect 10597 14025 10609 14059
rect 10643 14056 10655 14059
rect 11238 14056 11244 14068
rect 10643 14028 11244 14056
rect 10643 14025 10655 14028
rect 10597 14019 10655 14025
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 11606 14056 11612 14068
rect 11567 14028 11612 14056
rect 11606 14016 11612 14028
rect 11664 14016 11670 14068
rect 12161 14059 12219 14065
rect 12161 14025 12173 14059
rect 12207 14056 12219 14059
rect 12618 14056 12624 14068
rect 12207 14028 12624 14056
rect 12207 14025 12219 14028
rect 12161 14019 12219 14025
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 14921 14059 14979 14065
rect 14921 14056 14933 14059
rect 14516 14028 14933 14056
rect 14516 14016 14522 14028
rect 14921 14025 14933 14028
rect 14967 14056 14979 14059
rect 15473 14059 15531 14065
rect 15473 14056 15485 14059
rect 14967 14028 15485 14056
rect 14967 14025 14979 14028
rect 14921 14019 14979 14025
rect 15473 14025 15485 14028
rect 15519 14056 15531 14059
rect 15838 14056 15844 14068
rect 15519 14028 15844 14056
rect 15519 14025 15531 14028
rect 15473 14019 15531 14025
rect 15838 14016 15844 14028
rect 15896 14016 15902 14068
rect 16390 14056 16396 14068
rect 16351 14028 16396 14056
rect 16390 14016 16396 14028
rect 16448 14016 16454 14068
rect 17497 14059 17555 14065
rect 17497 14056 17509 14059
rect 16868 14028 17509 14056
rect 13354 13988 13360 14000
rect 13315 13960 13360 13988
rect 13354 13948 13360 13960
rect 13412 13948 13418 14000
rect 10962 13880 10968 13932
rect 11020 13920 11026 13932
rect 11057 13923 11115 13929
rect 11057 13920 11069 13923
rect 11020 13892 11069 13920
rect 11020 13880 11026 13892
rect 11057 13889 11069 13892
rect 11103 13889 11115 13923
rect 11057 13883 11115 13889
rect 11149 13923 11207 13929
rect 11149 13889 11161 13923
rect 11195 13889 11207 13923
rect 13538 13920 13544 13932
rect 13499 13892 13544 13920
rect 11149 13883 11207 13889
rect 10134 13852 10140 13864
rect 10095 13824 10140 13852
rect 10134 13812 10140 13824
rect 10192 13852 10198 13864
rect 10192 13824 10456 13852
rect 10192 13812 10198 13824
rect 10428 13716 10456 13824
rect 10505 13787 10563 13793
rect 10505 13753 10517 13787
rect 10551 13784 10563 13787
rect 10686 13784 10692 13796
rect 10551 13756 10692 13784
rect 10551 13753 10563 13756
rect 10505 13747 10563 13753
rect 10686 13744 10692 13756
rect 10744 13784 10750 13796
rect 10965 13787 11023 13793
rect 10965 13784 10977 13787
rect 10744 13756 10977 13784
rect 10744 13744 10750 13756
rect 10965 13753 10977 13756
rect 11011 13753 11023 13787
rect 10965 13747 11023 13753
rect 11164 13716 11192 13883
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 16868 13929 16896 14028
rect 17497 14025 17509 14028
rect 17543 14056 17555 14059
rect 18046 14056 18052 14068
rect 17543 14028 18052 14056
rect 17543 14025 17555 14028
rect 17497 14019 17555 14025
rect 18046 14016 18052 14028
rect 18104 14016 18110 14068
rect 18325 14059 18383 14065
rect 18325 14025 18337 14059
rect 18371 14056 18383 14059
rect 18598 14056 18604 14068
rect 18371 14028 18604 14056
rect 18371 14025 18383 14028
rect 18325 14019 18383 14025
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 18874 14056 18880 14068
rect 18835 14028 18880 14056
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 21634 14056 21640 14068
rect 21595 14028 21640 14056
rect 21634 14016 21640 14028
rect 21692 14016 21698 14068
rect 21818 14056 21824 14068
rect 21779 14028 21824 14056
rect 21818 14016 21824 14028
rect 21876 14016 21882 14068
rect 23106 14056 23112 14068
rect 23067 14028 23112 14056
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 23842 14056 23848 14068
rect 23803 14028 23848 14056
rect 23842 14016 23848 14028
rect 23900 14016 23906 14068
rect 16209 13923 16267 13929
rect 16209 13920 16221 13923
rect 15212 13892 16221 13920
rect 15212 13852 15240 13892
rect 16209 13889 16221 13892
rect 16255 13889 16267 13923
rect 16209 13883 16267 13889
rect 16853 13923 16911 13929
rect 16853 13889 16865 13923
rect 16899 13889 16911 13923
rect 16853 13883 16911 13889
rect 16945 13923 17003 13929
rect 16945 13889 16957 13923
rect 16991 13889 17003 13923
rect 18892 13920 18920 14016
rect 20349 13991 20407 13997
rect 20349 13957 20361 13991
rect 20395 13988 20407 13991
rect 20438 13988 20444 14000
rect 20395 13960 20444 13988
rect 20395 13957 20407 13960
rect 20349 13951 20407 13957
rect 20438 13948 20444 13960
rect 20496 13948 20502 14000
rect 18892 13892 19104 13920
rect 16945 13883 17003 13889
rect 15838 13852 15844 13864
rect 13740 13824 15240 13852
rect 15799 13824 15844 13852
rect 12529 13787 12587 13793
rect 12529 13753 12541 13787
rect 12575 13784 12587 13787
rect 13740 13784 13768 13824
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 16224 13852 16252 13883
rect 16224 13824 16528 13852
rect 12575 13756 13768 13784
rect 13808 13787 13866 13793
rect 12575 13753 12587 13756
rect 12529 13747 12587 13753
rect 13808 13753 13820 13787
rect 13854 13784 13866 13787
rect 13906 13784 13912 13796
rect 13854 13756 13912 13784
rect 13854 13753 13866 13756
rect 13808 13747 13866 13753
rect 13906 13744 13912 13756
rect 13964 13744 13970 13796
rect 16500 13784 16528 13824
rect 16574 13812 16580 13864
rect 16632 13852 16638 13864
rect 16960 13852 16988 13883
rect 17773 13855 17831 13861
rect 17773 13852 17785 13855
rect 16632 13824 17785 13852
rect 16632 13812 16638 13824
rect 17773 13821 17785 13824
rect 17819 13852 17831 13855
rect 18230 13852 18236 13864
rect 17819 13824 18236 13852
rect 17819 13821 17831 13824
rect 17773 13815 17831 13821
rect 18230 13812 18236 13824
rect 18288 13812 18294 13864
rect 18969 13855 19027 13861
rect 18969 13821 18981 13855
rect 19015 13821 19027 13855
rect 19076 13852 19104 13892
rect 22094 13880 22100 13932
rect 22152 13920 22158 13932
rect 22373 13923 22431 13929
rect 22373 13920 22385 13923
rect 22152 13892 22385 13920
rect 22152 13880 22158 13892
rect 22373 13889 22385 13892
rect 22419 13920 22431 13923
rect 23382 13920 23388 13932
rect 22419 13892 23388 13920
rect 22419 13889 22431 13892
rect 22373 13883 22431 13889
rect 23382 13880 23388 13892
rect 23440 13880 23446 13932
rect 23658 13880 23664 13932
rect 23716 13920 23722 13932
rect 23842 13920 23848 13932
rect 23716 13892 23848 13920
rect 23716 13880 23722 13892
rect 23842 13880 23848 13892
rect 23900 13880 23906 13932
rect 19225 13855 19283 13861
rect 19225 13852 19237 13855
rect 19076 13824 19237 13852
rect 18969 13815 19027 13821
rect 19225 13821 19237 13824
rect 19271 13821 19283 13855
rect 19225 13815 19283 13821
rect 16761 13787 16819 13793
rect 16761 13784 16773 13787
rect 16500 13756 16773 13784
rect 16761 13753 16773 13756
rect 16807 13753 16819 13787
rect 18984 13784 19012 13815
rect 20806 13812 20812 13864
rect 20864 13852 20870 13864
rect 20901 13855 20959 13861
rect 20901 13852 20913 13855
rect 20864 13824 20913 13852
rect 20864 13812 20870 13824
rect 20901 13821 20913 13824
rect 20947 13821 20959 13855
rect 21358 13852 21364 13864
rect 21319 13824 21364 13852
rect 20901 13815 20959 13821
rect 21358 13812 21364 13824
rect 21416 13812 21422 13864
rect 22278 13852 22284 13864
rect 22239 13824 22284 13852
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 23477 13855 23535 13861
rect 23477 13821 23489 13855
rect 23523 13852 23535 13855
rect 24026 13852 24032 13864
rect 23523 13824 24032 13852
rect 23523 13821 23535 13824
rect 23477 13815 23535 13821
rect 24026 13812 24032 13824
rect 24084 13812 24090 13864
rect 24121 13855 24179 13861
rect 24121 13821 24133 13855
rect 24167 13852 24179 13855
rect 24946 13852 24952 13864
rect 24167 13824 24952 13852
rect 24167 13821 24179 13824
rect 24121 13815 24179 13821
rect 24946 13812 24952 13824
rect 25004 13812 25010 13864
rect 19058 13784 19064 13796
rect 18984 13756 19064 13784
rect 16761 13747 16819 13753
rect 19058 13744 19064 13756
rect 19116 13744 19122 13796
rect 24394 13793 24400 13796
rect 24388 13784 24400 13793
rect 24355 13756 24400 13784
rect 24388 13747 24400 13756
rect 24394 13744 24400 13747
rect 24452 13744 24458 13796
rect 11698 13716 11704 13728
rect 10428 13688 11704 13716
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 13078 13716 13084 13728
rect 13039 13688 13084 13716
rect 13078 13676 13084 13688
rect 13136 13716 13142 13728
rect 14182 13716 14188 13728
rect 13136 13688 14188 13716
rect 13136 13676 13142 13688
rect 14182 13676 14188 13688
rect 14240 13676 14246 13728
rect 22186 13716 22192 13728
rect 22147 13688 22192 13716
rect 22186 13676 22192 13688
rect 22244 13676 22250 13728
rect 25498 13716 25504 13728
rect 25459 13688 25504 13716
rect 25498 13676 25504 13688
rect 25556 13676 25562 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 11698 13512 11704 13524
rect 11659 13484 11704 13512
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 12342 13512 12348 13524
rect 12303 13484 12348 13512
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 12713 13515 12771 13521
rect 12713 13481 12725 13515
rect 12759 13512 12771 13515
rect 13906 13512 13912 13524
rect 12759 13484 13912 13512
rect 12759 13481 12771 13484
rect 12713 13475 12771 13481
rect 13906 13472 13912 13484
rect 13964 13512 13970 13524
rect 14826 13512 14832 13524
rect 13964 13484 14832 13512
rect 13964 13472 13970 13484
rect 14826 13472 14832 13484
rect 14884 13512 14890 13524
rect 15013 13515 15071 13521
rect 15013 13512 15025 13515
rect 14884 13484 15025 13512
rect 14884 13472 14890 13484
rect 15013 13481 15025 13484
rect 15059 13481 15071 13515
rect 15286 13512 15292 13524
rect 15247 13484 15292 13512
rect 15013 13475 15071 13481
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 18230 13512 18236 13524
rect 18191 13484 18236 13512
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 19058 13472 19064 13524
rect 19116 13512 19122 13524
rect 19153 13515 19211 13521
rect 19153 13512 19165 13515
rect 19116 13484 19165 13512
rect 19116 13472 19122 13484
rect 19153 13481 19165 13484
rect 19199 13481 19211 13515
rect 20898 13512 20904 13524
rect 20859 13484 20904 13512
rect 19153 13475 19211 13481
rect 20898 13472 20904 13484
rect 20956 13472 20962 13524
rect 21545 13515 21603 13521
rect 21545 13481 21557 13515
rect 21591 13512 21603 13515
rect 22186 13512 22192 13524
rect 21591 13484 22192 13512
rect 21591 13481 21603 13484
rect 21545 13475 21603 13481
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 23474 13512 23480 13524
rect 23435 13484 23480 13512
rect 23474 13472 23480 13484
rect 23532 13472 23538 13524
rect 24581 13515 24639 13521
rect 24581 13481 24593 13515
rect 24627 13512 24639 13515
rect 24670 13512 24676 13524
rect 24627 13484 24676 13512
rect 24627 13481 24639 13484
rect 24581 13475 24639 13481
rect 24670 13472 24676 13484
rect 24728 13472 24734 13524
rect 16758 13404 16764 13456
rect 16816 13444 16822 13456
rect 17098 13447 17156 13453
rect 17098 13444 17110 13447
rect 16816 13416 17110 13444
rect 16816 13404 16822 13416
rect 17098 13413 17110 13416
rect 17144 13413 17156 13447
rect 17098 13407 17156 13413
rect 17954 13404 17960 13456
rect 18012 13444 18018 13456
rect 18785 13447 18843 13453
rect 18785 13444 18797 13447
rect 18012 13416 18797 13444
rect 18012 13404 18018 13416
rect 18785 13413 18797 13416
rect 18831 13413 18843 13447
rect 18785 13407 18843 13413
rect 19426 13404 19432 13456
rect 19484 13444 19490 13456
rect 19613 13447 19671 13453
rect 19613 13444 19625 13447
rect 19484 13416 19625 13444
rect 19484 13404 19490 13416
rect 19613 13413 19625 13416
rect 19659 13413 19671 13447
rect 19613 13407 19671 13413
rect 21913 13447 21971 13453
rect 21913 13413 21925 13447
rect 21959 13444 21971 13447
rect 22094 13444 22100 13456
rect 21959 13416 22100 13444
rect 21959 13413 21971 13416
rect 21913 13407 21971 13413
rect 22094 13404 22100 13416
rect 22152 13404 22158 13456
rect 10410 13336 10416 13388
rect 10468 13376 10474 13388
rect 10577 13379 10635 13385
rect 10577 13376 10589 13379
rect 10468 13348 10589 13376
rect 10468 13336 10474 13348
rect 10577 13345 10589 13348
rect 10623 13376 10635 13379
rect 10870 13376 10876 13388
rect 10623 13348 10876 13376
rect 10623 13345 10635 13348
rect 10577 13339 10635 13345
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 12802 13376 12808 13388
rect 12763 13348 12808 13376
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 15654 13376 15660 13388
rect 15615 13348 15660 13376
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 15749 13379 15807 13385
rect 15749 13345 15761 13379
rect 15795 13376 15807 13379
rect 16022 13376 16028 13388
rect 15795 13348 16028 13376
rect 15795 13345 15807 13348
rect 15749 13339 15807 13345
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16853 13379 16911 13385
rect 16853 13345 16865 13379
rect 16899 13376 16911 13379
rect 16942 13376 16948 13388
rect 16899 13348 16948 13376
rect 16899 13345 16911 13348
rect 16853 13339 16911 13345
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 19242 13336 19248 13388
rect 19300 13376 19306 13388
rect 22370 13385 22376 13388
rect 19337 13379 19395 13385
rect 19337 13376 19349 13379
rect 19300 13348 19349 13376
rect 19300 13336 19306 13348
rect 19337 13345 19349 13348
rect 19383 13376 19395 13379
rect 20073 13379 20131 13385
rect 20073 13376 20085 13379
rect 19383 13348 20085 13376
rect 19383 13345 19395 13348
rect 19337 13339 19395 13345
rect 20073 13345 20085 13348
rect 20119 13345 20131 13379
rect 20073 13339 20131 13345
rect 22364 13339 22376 13385
rect 22428 13376 22434 13388
rect 24946 13376 24952 13388
rect 22428 13348 22464 13376
rect 24859 13348 24952 13376
rect 22370 13336 22376 13339
rect 22428 13336 22434 13348
rect 24946 13336 24952 13348
rect 25004 13376 25010 13388
rect 25682 13376 25688 13388
rect 25004 13348 25688 13376
rect 25004 13336 25010 13348
rect 25682 13336 25688 13348
rect 25740 13336 25746 13388
rect 9674 13308 9680 13320
rect 9635 13280 9680 13308
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 9858 13268 9864 13320
rect 9916 13308 9922 13320
rect 10318 13308 10324 13320
rect 9916 13280 10324 13308
rect 9916 13268 9922 13280
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 14568 13240 14596 13271
rect 14826 13268 14832 13320
rect 14884 13308 14890 13320
rect 15841 13311 15899 13317
rect 15841 13308 15853 13311
rect 14884 13280 15853 13308
rect 14884 13268 14890 13280
rect 15841 13277 15853 13280
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 22002 13268 22008 13320
rect 22060 13308 22066 13320
rect 22097 13311 22155 13317
rect 22097 13308 22109 13311
rect 22060 13280 22109 13308
rect 22060 13268 22066 13280
rect 22097 13277 22109 13280
rect 22143 13277 22155 13311
rect 25038 13308 25044 13320
rect 24999 13280 25044 13308
rect 22097 13271 22155 13277
rect 25038 13268 25044 13280
rect 25096 13268 25102 13320
rect 25133 13311 25191 13317
rect 25133 13277 25145 13311
rect 25179 13308 25191 13311
rect 25498 13308 25504 13320
rect 25179 13280 25504 13308
rect 25179 13277 25191 13280
rect 25133 13271 25191 13277
rect 25498 13268 25504 13280
rect 25556 13308 25562 13320
rect 25958 13308 25964 13320
rect 25556 13280 25964 13308
rect 25556 13268 25562 13280
rect 25958 13268 25964 13280
rect 26016 13268 26022 13320
rect 24213 13243 24271 13249
rect 14568 13212 16896 13240
rect 16868 13184 16896 13212
rect 24213 13209 24225 13243
rect 24259 13240 24271 13243
rect 24394 13240 24400 13252
rect 24259 13212 24400 13240
rect 24259 13209 24271 13212
rect 24213 13203 24271 13209
rect 24394 13200 24400 13212
rect 24452 13240 24458 13252
rect 25222 13240 25228 13252
rect 24452 13212 25228 13240
rect 24452 13200 24458 13212
rect 25222 13200 25228 13212
rect 25280 13200 25286 13252
rect 9858 13132 9864 13184
rect 9916 13172 9922 13184
rect 10137 13175 10195 13181
rect 10137 13172 10149 13175
rect 9916 13144 10149 13172
rect 9916 13132 9922 13144
rect 10137 13141 10149 13144
rect 10183 13141 10195 13175
rect 16390 13172 16396 13184
rect 16351 13144 16396 13172
rect 10137 13135 10195 13141
rect 16390 13132 16396 13144
rect 16448 13172 16454 13184
rect 16574 13172 16580 13184
rect 16448 13144 16580 13172
rect 16448 13132 16454 13144
rect 16574 13132 16580 13144
rect 16632 13132 16638 13184
rect 16850 13132 16856 13184
rect 16908 13132 16914 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 9732 12940 10609 12968
rect 9732 12928 9738 12940
rect 10597 12937 10609 12940
rect 10643 12937 10655 12971
rect 10778 12968 10784 12980
rect 10739 12940 10784 12968
rect 10597 12931 10655 12937
rect 10321 12903 10379 12909
rect 10321 12869 10333 12903
rect 10367 12900 10379 12903
rect 10410 12900 10416 12912
rect 10367 12872 10416 12900
rect 10367 12869 10379 12872
rect 10321 12863 10379 12869
rect 10410 12860 10416 12872
rect 10468 12860 10474 12912
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12832 9827 12835
rect 10042 12832 10048 12844
rect 9815 12804 10048 12832
rect 9815 12801 9827 12804
rect 9769 12795 9827 12801
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 9401 12767 9459 12773
rect 9401 12733 9413 12767
rect 9447 12764 9459 12767
rect 9490 12764 9496 12776
rect 9447 12736 9496 12764
rect 9447 12733 9459 12736
rect 9401 12727 9459 12733
rect 9490 12724 9496 12736
rect 9548 12724 9554 12776
rect 10612 12764 10640 12931
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 14458 12928 14464 12980
rect 14516 12968 14522 12980
rect 14826 12968 14832 12980
rect 14516 12940 14832 12968
rect 14516 12928 14522 12940
rect 14826 12928 14832 12940
rect 14884 12968 14890 12980
rect 15105 12971 15163 12977
rect 15105 12968 15117 12971
rect 14884 12940 15117 12968
rect 14884 12928 14890 12940
rect 15105 12937 15117 12940
rect 15151 12937 15163 12971
rect 16022 12968 16028 12980
rect 15983 12940 16028 12968
rect 15105 12931 15163 12937
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 16758 12928 16764 12980
rect 16816 12968 16822 12980
rect 17402 12968 17408 12980
rect 16816 12940 17408 12968
rect 16816 12928 16822 12940
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 22005 12971 22063 12977
rect 22005 12937 22017 12971
rect 22051 12968 22063 12971
rect 22186 12968 22192 12980
rect 22051 12940 22192 12968
rect 22051 12937 22063 12940
rect 22005 12931 22063 12937
rect 22186 12928 22192 12940
rect 22244 12928 22250 12980
rect 23474 12968 23480 12980
rect 23435 12940 23480 12968
rect 23474 12928 23480 12940
rect 23532 12928 23538 12980
rect 24762 12928 24768 12980
rect 24820 12968 24826 12980
rect 25038 12968 25044 12980
rect 24820 12940 25044 12968
rect 24820 12928 24826 12940
rect 25038 12928 25044 12940
rect 25096 12968 25102 12980
rect 26329 12971 26387 12977
rect 26329 12968 26341 12971
rect 25096 12940 26341 12968
rect 25096 12928 25102 12940
rect 26329 12937 26341 12940
rect 26375 12937 26387 12971
rect 26329 12931 26387 12937
rect 12161 12903 12219 12909
rect 12161 12900 12173 12903
rect 11256 12872 12173 12900
rect 11256 12844 11284 12872
rect 12161 12869 12173 12872
rect 12207 12869 12219 12903
rect 12161 12863 12219 12869
rect 15194 12860 15200 12912
rect 15252 12900 15258 12912
rect 16206 12900 16212 12912
rect 15252 12872 16212 12900
rect 15252 12860 15258 12872
rect 16206 12860 16212 12872
rect 16264 12860 16270 12912
rect 16393 12903 16451 12909
rect 16393 12869 16405 12903
rect 16439 12869 16451 12903
rect 16393 12863 16451 12869
rect 11238 12832 11244 12844
rect 11199 12804 11244 12832
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 11425 12835 11483 12841
rect 11425 12801 11437 12835
rect 11471 12832 11483 12835
rect 11790 12832 11796 12844
rect 11471 12804 11796 12832
rect 11471 12801 11483 12804
rect 11425 12795 11483 12801
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12832 12771 12835
rect 12986 12832 12992 12844
rect 12759 12804 12992 12832
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 15470 12792 15476 12844
rect 15528 12792 15534 12844
rect 11149 12767 11207 12773
rect 11149 12764 11161 12767
rect 10612 12736 11161 12764
rect 11149 12733 11161 12736
rect 11195 12733 11207 12767
rect 11149 12727 11207 12733
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12764 12495 12767
rect 12618 12764 12624 12776
rect 12483 12736 12624 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 12618 12724 12624 12736
rect 12676 12724 12682 12776
rect 13725 12767 13783 12773
rect 13725 12733 13737 12767
rect 13771 12764 13783 12767
rect 14550 12764 14556 12776
rect 13771 12736 14556 12764
rect 13771 12733 13783 12736
rect 13725 12727 13783 12733
rect 14550 12724 14556 12736
rect 14608 12724 14614 12776
rect 15488 12764 15516 12792
rect 16408 12776 16436 12863
rect 16574 12792 16580 12844
rect 16632 12832 16638 12844
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16632 12804 16957 12832
rect 16632 12792 16638 12804
rect 16945 12801 16957 12804
rect 16991 12801 17003 12835
rect 18322 12832 18328 12844
rect 18283 12804 18328 12832
rect 16945 12795 17003 12801
rect 18322 12792 18328 12804
rect 18380 12792 18386 12844
rect 19334 12792 19340 12844
rect 19392 12832 19398 12844
rect 19981 12835 20039 12841
rect 19981 12832 19993 12835
rect 19392 12804 19993 12832
rect 19392 12792 19398 12804
rect 19981 12801 19993 12804
rect 20027 12832 20039 12835
rect 20441 12835 20499 12841
rect 20441 12832 20453 12835
rect 20027 12804 20453 12832
rect 20027 12801 20039 12804
rect 19981 12795 20039 12801
rect 20441 12801 20453 12804
rect 20487 12801 20499 12835
rect 20441 12795 20499 12801
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 20993 12835 21051 12841
rect 20993 12832 21005 12835
rect 20772 12804 21005 12832
rect 20772 12792 20778 12804
rect 20993 12801 21005 12804
rect 21039 12801 21051 12835
rect 20993 12795 21051 12801
rect 21545 12835 21603 12841
rect 21545 12801 21557 12835
rect 21591 12832 21603 12835
rect 22370 12832 22376 12844
rect 21591 12804 22376 12832
rect 21591 12801 21603 12804
rect 21545 12795 21603 12801
rect 22370 12792 22376 12804
rect 22428 12832 22434 12844
rect 22557 12835 22615 12841
rect 22557 12832 22569 12835
rect 22428 12804 22569 12832
rect 22428 12792 22434 12804
rect 22557 12801 22569 12804
rect 22603 12832 22615 12835
rect 22646 12832 22652 12844
rect 22603 12804 22652 12832
rect 22603 12801 22615 12804
rect 22557 12795 22615 12801
rect 22646 12792 22652 12804
rect 22704 12832 22710 12844
rect 23017 12835 23075 12841
rect 23017 12832 23029 12835
rect 22704 12804 23029 12832
rect 22704 12792 22710 12804
rect 23017 12801 23029 12804
rect 23063 12801 23075 12835
rect 23492 12832 23520 12928
rect 25682 12900 25688 12912
rect 25643 12872 25688 12900
rect 25682 12860 25688 12872
rect 25740 12860 25746 12912
rect 25958 12900 25964 12912
rect 25919 12872 25964 12900
rect 25958 12860 25964 12872
rect 26016 12860 26022 12912
rect 23492 12804 23796 12832
rect 23017 12795 23075 12801
rect 15488 12736 15884 12764
rect 10042 12656 10048 12708
rect 10100 12696 10106 12708
rect 10318 12696 10324 12708
rect 10100 12668 10324 12696
rect 10100 12656 10106 12668
rect 10318 12656 10324 12668
rect 10376 12656 10382 12708
rect 13633 12699 13691 12705
rect 13633 12665 13645 12699
rect 13679 12696 13691 12699
rect 13992 12699 14050 12705
rect 13992 12696 14004 12699
rect 13679 12668 14004 12696
rect 13679 12665 13691 12668
rect 13633 12659 13691 12665
rect 13992 12665 14004 12668
rect 14038 12696 14050 12699
rect 15470 12696 15476 12708
rect 14038 12668 15476 12696
rect 14038 12665 14050 12668
rect 13992 12659 14050 12665
rect 15470 12656 15476 12668
rect 15528 12656 15534 12708
rect 12250 12588 12256 12640
rect 12308 12628 12314 12640
rect 12802 12628 12808 12640
rect 12308 12600 12808 12628
rect 12308 12588 12314 12600
rect 12802 12588 12808 12600
rect 12860 12628 12866 12640
rect 13173 12631 13231 12637
rect 13173 12628 13185 12631
rect 12860 12600 13185 12628
rect 12860 12588 12866 12600
rect 13173 12597 13185 12600
rect 13219 12597 13231 12631
rect 15654 12628 15660 12640
rect 15615 12600 15660 12628
rect 13173 12591 13231 12597
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 15856 12628 15884 12736
rect 16390 12724 16396 12776
rect 16448 12724 16454 12776
rect 17862 12764 17868 12776
rect 16776 12736 17868 12764
rect 16776 12640 16804 12736
rect 17862 12724 17868 12736
rect 17920 12724 17926 12776
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12764 18107 12767
rect 18230 12764 18236 12776
rect 18095 12736 18236 12764
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 18230 12724 18236 12736
rect 18288 12764 18294 12776
rect 18782 12764 18788 12776
rect 18288 12736 18788 12764
rect 18288 12724 18294 12736
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 19245 12767 19303 12773
rect 19245 12733 19257 12767
rect 19291 12764 19303 12767
rect 19889 12767 19947 12773
rect 19889 12764 19901 12767
rect 19291 12736 19901 12764
rect 19291 12733 19303 12736
rect 19245 12727 19303 12733
rect 19889 12733 19901 12736
rect 19935 12764 19947 12767
rect 20162 12764 20168 12776
rect 19935 12736 20168 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 20162 12724 20168 12736
rect 20220 12724 20226 12776
rect 20898 12724 20904 12776
rect 20956 12764 20962 12776
rect 21913 12767 21971 12773
rect 21913 12764 21925 12767
rect 20956 12736 21925 12764
rect 20956 12724 20962 12736
rect 21913 12733 21925 12736
rect 21959 12764 21971 12767
rect 22465 12767 22523 12773
rect 22465 12764 22477 12767
rect 21959 12736 22477 12764
rect 21959 12733 21971 12736
rect 21913 12727 21971 12733
rect 22465 12733 22477 12736
rect 22511 12764 22523 12767
rect 22830 12764 22836 12776
rect 22511 12736 22836 12764
rect 22511 12733 22523 12736
rect 22465 12727 22523 12733
rect 22830 12724 22836 12736
rect 22888 12724 22894 12776
rect 23658 12764 23664 12776
rect 23619 12736 23664 12764
rect 23658 12724 23664 12736
rect 23716 12724 23722 12776
rect 23768 12764 23796 12804
rect 23917 12767 23975 12773
rect 23917 12764 23929 12767
rect 23768 12736 23929 12764
rect 23917 12733 23929 12736
rect 23963 12733 23975 12767
rect 23917 12727 23975 12733
rect 16853 12699 16911 12705
rect 16853 12665 16865 12699
rect 16899 12696 16911 12699
rect 17770 12696 17776 12708
rect 16899 12668 17776 12696
rect 16899 12665 16911 12668
rect 16853 12659 16911 12665
rect 17770 12656 17776 12668
rect 17828 12656 17834 12708
rect 18969 12699 19027 12705
rect 18969 12665 18981 12699
rect 19015 12696 19027 12699
rect 19797 12699 19855 12705
rect 19797 12696 19809 12699
rect 19015 12668 19809 12696
rect 19015 12665 19027 12668
rect 18969 12659 19027 12665
rect 19797 12665 19809 12668
rect 19843 12696 19855 12699
rect 20714 12696 20720 12708
rect 19843 12668 20720 12696
rect 19843 12665 19855 12668
rect 19797 12659 19855 12665
rect 20714 12656 20720 12668
rect 20772 12656 20778 12708
rect 24118 12656 24124 12708
rect 24176 12696 24182 12708
rect 24670 12696 24676 12708
rect 24176 12668 24676 12696
rect 24176 12656 24182 12668
rect 24670 12656 24676 12668
rect 24728 12656 24734 12708
rect 16114 12628 16120 12640
rect 15856 12600 16120 12628
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 16758 12628 16764 12640
rect 16719 12600 16764 12628
rect 16758 12588 16764 12600
rect 16816 12588 16822 12640
rect 19426 12628 19432 12640
rect 19387 12600 19432 12628
rect 19426 12588 19432 12600
rect 19484 12588 19490 12640
rect 20898 12628 20904 12640
rect 20859 12600 20904 12628
rect 20898 12588 20904 12600
rect 20956 12588 20962 12640
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 22373 12631 22431 12637
rect 22373 12628 22385 12631
rect 22152 12600 22385 12628
rect 22152 12588 22158 12600
rect 22373 12597 22385 12600
rect 22419 12597 22431 12631
rect 22373 12591 22431 12597
rect 25041 12631 25099 12637
rect 25041 12597 25053 12631
rect 25087 12628 25099 12631
rect 25222 12628 25228 12640
rect 25087 12600 25228 12628
rect 25087 12597 25099 12600
rect 25041 12591 25099 12597
rect 25222 12588 25228 12600
rect 25280 12588 25286 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10321 12427 10379 12433
rect 10321 12424 10333 12427
rect 10100 12396 10333 12424
rect 10100 12384 10106 12396
rect 10321 12393 10333 12396
rect 10367 12393 10379 12427
rect 12618 12424 12624 12436
rect 12579 12396 12624 12424
rect 10321 12387 10379 12393
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 12805 12427 12863 12433
rect 12805 12393 12817 12427
rect 12851 12424 12863 12427
rect 13446 12424 13452 12436
rect 12851 12396 13452 12424
rect 12851 12393 12863 12396
rect 12805 12387 12863 12393
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 13633 12427 13691 12433
rect 13633 12393 13645 12427
rect 13679 12424 13691 12427
rect 13722 12424 13728 12436
rect 13679 12396 13728 12424
rect 13679 12393 13691 12396
rect 13633 12387 13691 12393
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 15286 12424 15292 12436
rect 15247 12396 15292 12424
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 16482 12424 16488 12436
rect 15528 12396 15976 12424
rect 16443 12396 16488 12424
rect 15528 12384 15534 12396
rect 1578 12316 1584 12368
rect 1636 12365 1642 12368
rect 1636 12359 1700 12365
rect 1636 12325 1654 12359
rect 1688 12325 1700 12359
rect 1636 12319 1700 12325
rect 1636 12316 1642 12319
rect 10134 12316 10140 12368
rect 10192 12356 10198 12368
rect 10934 12359 10992 12365
rect 10934 12356 10946 12359
rect 10192 12328 10946 12356
rect 10192 12316 10198 12328
rect 10934 12325 10946 12328
rect 10980 12325 10992 12359
rect 10934 12319 10992 12325
rect 15838 12316 15844 12368
rect 15896 12316 15902 12368
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 2038 12288 2044 12300
rect 1443 12260 2044 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 9916 12260 10057 12288
rect 9916 12248 9922 12260
rect 10045 12257 10057 12260
rect 10091 12288 10103 12291
rect 10689 12291 10747 12297
rect 10689 12288 10701 12291
rect 10091 12260 10701 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10689 12257 10701 12260
rect 10735 12288 10747 12291
rect 12434 12288 12440 12300
rect 10735 12260 12440 12288
rect 10735 12257 10747 12260
rect 10689 12251 10747 12257
rect 12434 12248 12440 12260
rect 12492 12248 12498 12300
rect 13170 12288 13176 12300
rect 13131 12260 13176 12288
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 14001 12291 14059 12297
rect 14001 12257 14013 12291
rect 14047 12288 14059 12291
rect 14366 12288 14372 12300
rect 14047 12260 14372 12288
rect 14047 12257 14059 12260
rect 14001 12251 14059 12257
rect 14366 12248 14372 12260
rect 14424 12248 14430 12300
rect 15470 12248 15476 12300
rect 15528 12288 15534 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15528 12260 15669 12288
rect 15528 12248 15534 12260
rect 15657 12257 15669 12260
rect 15703 12288 15715 12291
rect 15856 12288 15884 12316
rect 15703 12260 15884 12288
rect 15703 12257 15715 12260
rect 15657 12251 15715 12257
rect 12342 12180 12348 12232
rect 12400 12220 12406 12232
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 12400 12192 13277 12220
rect 12400 12180 12406 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 13354 12180 13360 12232
rect 13412 12220 13418 12232
rect 14093 12223 14151 12229
rect 13412 12192 13457 12220
rect 13412 12180 13418 12192
rect 14093 12189 14105 12223
rect 14139 12220 14151 12223
rect 14182 12220 14188 12232
rect 14139 12192 14188 12220
rect 14139 12189 14151 12192
rect 14093 12183 14151 12189
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12220 14335 12223
rect 14458 12220 14464 12232
rect 14323 12192 14464 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 15746 12220 15752 12232
rect 14783 12192 15752 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 15948 12220 15976 12396
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 17218 12424 17224 12436
rect 17131 12396 17224 12424
rect 17218 12384 17224 12396
rect 17276 12424 17282 12436
rect 17494 12424 17500 12436
rect 17276 12396 17500 12424
rect 17276 12384 17282 12396
rect 17494 12384 17500 12396
rect 17552 12384 17558 12436
rect 17862 12384 17868 12436
rect 17920 12424 17926 12436
rect 17957 12427 18015 12433
rect 17957 12424 17969 12427
rect 17920 12396 17969 12424
rect 17920 12384 17926 12396
rect 17957 12393 17969 12396
rect 18003 12393 18015 12427
rect 18230 12424 18236 12436
rect 18191 12396 18236 12424
rect 17957 12387 18015 12393
rect 18230 12384 18236 12396
rect 18288 12384 18294 12436
rect 19242 12424 19248 12436
rect 19203 12396 19248 12424
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 21177 12427 21235 12433
rect 21177 12393 21189 12427
rect 21223 12424 21235 12427
rect 22094 12424 22100 12436
rect 21223 12396 22100 12424
rect 21223 12393 21235 12396
rect 21177 12387 21235 12393
rect 22094 12384 22100 12396
rect 22152 12424 22158 12436
rect 22152 12396 22245 12424
rect 22152 12384 22158 12396
rect 22646 12384 22652 12436
rect 22704 12424 22710 12436
rect 23569 12427 23627 12433
rect 23569 12424 23581 12427
rect 22704 12396 23581 12424
rect 22704 12384 22710 12396
rect 23569 12393 23581 12396
rect 23615 12393 23627 12427
rect 23569 12387 23627 12393
rect 23842 12384 23848 12436
rect 23900 12424 23906 12436
rect 24673 12427 24731 12433
rect 23900 12396 24624 12424
rect 23900 12384 23906 12396
rect 20806 12316 20812 12368
rect 20864 12356 20870 12368
rect 20990 12356 20996 12368
rect 20864 12328 20996 12356
rect 20864 12316 20870 12328
rect 20990 12316 20996 12328
rect 21048 12316 21054 12368
rect 23658 12356 23664 12368
rect 22204 12328 23664 12356
rect 19150 12288 19156 12300
rect 19111 12260 19156 12288
rect 19150 12248 19156 12260
rect 19208 12248 19214 12300
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 19613 12291 19671 12297
rect 19613 12288 19625 12291
rect 19484 12260 19625 12288
rect 19484 12248 19490 12260
rect 19613 12257 19625 12260
rect 19659 12288 19671 12291
rect 19978 12288 19984 12300
rect 19659 12260 19984 12288
rect 19659 12257 19671 12260
rect 19613 12251 19671 12257
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 20717 12291 20775 12297
rect 20717 12257 20729 12291
rect 20763 12288 20775 12291
rect 20898 12288 20904 12300
rect 20763 12260 20904 12288
rect 20763 12257 20775 12260
rect 20717 12251 20775 12257
rect 17310 12220 17316 12232
rect 15896 12192 15976 12220
rect 17271 12192 17316 12220
rect 15896 12180 15902 12192
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12220 17555 12223
rect 17862 12220 17868 12232
rect 17543 12192 17868 12220
rect 17543 12189 17555 12192
rect 17497 12183 17555 12189
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 19518 12180 19524 12232
rect 19576 12220 19582 12232
rect 19705 12223 19763 12229
rect 19705 12220 19717 12223
rect 19576 12192 19717 12220
rect 19576 12180 19582 12192
rect 19705 12189 19717 12192
rect 19751 12189 19763 12223
rect 19886 12220 19892 12232
rect 19847 12192 19892 12220
rect 19705 12183 19763 12189
rect 19886 12180 19892 12192
rect 19944 12180 19950 12232
rect 18598 12112 18604 12164
rect 18656 12152 18662 12164
rect 18969 12155 19027 12161
rect 18969 12152 18981 12155
rect 18656 12124 18981 12152
rect 18656 12112 18662 12124
rect 18969 12121 18981 12124
rect 19015 12152 19027 12155
rect 20732 12152 20760 12251
rect 20898 12248 20904 12260
rect 20956 12288 20962 12300
rect 21729 12291 21787 12297
rect 21729 12288 21741 12291
rect 20956 12260 21741 12288
rect 20956 12248 20962 12260
rect 21729 12257 21741 12260
rect 21775 12288 21787 12291
rect 22002 12288 22008 12300
rect 21775 12260 22008 12288
rect 21775 12257 21787 12260
rect 21729 12251 21787 12257
rect 22002 12248 22008 12260
rect 22060 12288 22066 12300
rect 22204 12297 22232 12328
rect 23658 12316 23664 12328
rect 23716 12356 23722 12368
rect 24489 12359 24547 12365
rect 24489 12356 24501 12359
rect 23716 12328 24501 12356
rect 23716 12316 23722 12328
rect 24489 12325 24501 12328
rect 24535 12325 24547 12359
rect 24596 12356 24624 12396
rect 24673 12393 24685 12427
rect 24719 12424 24731 12427
rect 24762 12424 24768 12436
rect 24719 12396 24768 12424
rect 24719 12393 24731 12396
rect 24673 12387 24731 12393
rect 24762 12384 24768 12396
rect 24820 12384 24826 12436
rect 25498 12356 25504 12368
rect 24596 12328 25504 12356
rect 24489 12319 24547 12325
rect 25498 12316 25504 12328
rect 25556 12316 25562 12368
rect 22462 12297 22468 12300
rect 22189 12291 22247 12297
rect 22189 12288 22201 12291
rect 22060 12260 22201 12288
rect 22060 12248 22066 12260
rect 22189 12257 22201 12260
rect 22235 12257 22247 12291
rect 22189 12251 22247 12257
rect 22456 12251 22468 12297
rect 22520 12288 22526 12300
rect 22520 12260 22556 12288
rect 22462 12248 22468 12251
rect 22520 12248 22526 12260
rect 22922 12248 22928 12300
rect 22980 12288 22986 12300
rect 23842 12288 23848 12300
rect 22980 12260 23848 12288
rect 22980 12248 22986 12260
rect 23842 12248 23848 12260
rect 23900 12248 23906 12300
rect 25038 12288 25044 12300
rect 24999 12260 25044 12288
rect 25038 12248 25044 12260
rect 25096 12248 25102 12300
rect 25133 12291 25191 12297
rect 25133 12257 25145 12291
rect 25179 12288 25191 12291
rect 25314 12288 25320 12300
rect 25179 12260 25320 12288
rect 25179 12257 25191 12260
rect 25133 12251 25191 12257
rect 25314 12248 25320 12260
rect 25372 12248 25378 12300
rect 25222 12180 25228 12232
rect 25280 12220 25286 12232
rect 25280 12192 25325 12220
rect 25280 12180 25286 12192
rect 19015 12124 20760 12152
rect 19015 12121 19027 12124
rect 18969 12115 19027 12121
rect 2774 12044 2780 12096
rect 2832 12084 2838 12096
rect 9309 12087 9367 12093
rect 2832 12056 2877 12084
rect 2832 12044 2838 12056
rect 9309 12053 9321 12087
rect 9355 12084 9367 12087
rect 9582 12084 9588 12096
rect 9355 12056 9588 12084
rect 9355 12053 9367 12056
rect 9309 12047 9367 12053
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 11422 12044 11428 12096
rect 11480 12084 11486 12096
rect 11790 12084 11796 12096
rect 11480 12056 11796 12084
rect 11480 12044 11486 12056
rect 11790 12044 11796 12056
rect 11848 12084 11854 12096
rect 12069 12087 12127 12093
rect 12069 12084 12081 12087
rect 11848 12056 12081 12084
rect 11848 12044 11854 12056
rect 12069 12053 12081 12056
rect 12115 12053 12127 12087
rect 12069 12047 12127 12053
rect 15105 12087 15163 12093
rect 15105 12053 15117 12087
rect 15151 12084 15163 12087
rect 15378 12084 15384 12096
rect 15151 12056 15384 12084
rect 15151 12053 15163 12056
rect 15105 12047 15163 12053
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 16853 12087 16911 12093
rect 16853 12084 16865 12087
rect 16632 12056 16865 12084
rect 16632 12044 16638 12056
rect 16853 12053 16865 12056
rect 16899 12053 16911 12087
rect 18690 12084 18696 12096
rect 18651 12056 18696 12084
rect 16853 12047 16911 12053
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 18782 12044 18788 12096
rect 18840 12084 18846 12096
rect 20257 12087 20315 12093
rect 20257 12084 20269 12087
rect 18840 12056 20269 12084
rect 18840 12044 18846 12056
rect 20257 12053 20269 12056
rect 20303 12053 20315 12087
rect 24210 12084 24216 12096
rect 24171 12056 24216 12084
rect 20257 12047 20315 12053
rect 24210 12044 24216 12056
rect 24268 12044 24274 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 10229 11883 10287 11889
rect 10229 11880 10241 11883
rect 10192 11852 10241 11880
rect 10192 11840 10198 11852
rect 10229 11849 10241 11852
rect 10275 11849 10287 11883
rect 10229 11843 10287 11849
rect 12253 11883 12311 11889
rect 12253 11849 12265 11883
rect 12299 11880 12311 11883
rect 13354 11880 13360 11892
rect 12299 11852 13360 11880
rect 12299 11849 12311 11852
rect 12253 11843 12311 11849
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 13538 11880 13544 11892
rect 13499 11852 13544 11880
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 17129 11883 17187 11889
rect 15120 11852 16988 11880
rect 14550 11772 14556 11824
rect 14608 11812 14614 11824
rect 15120 11812 15148 11852
rect 16960 11824 16988 11852
rect 17129 11849 17141 11883
rect 17175 11880 17187 11883
rect 17310 11880 17316 11892
rect 17175 11852 17316 11880
rect 17175 11849 17187 11852
rect 17129 11843 17187 11849
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 17494 11880 17500 11892
rect 17455 11852 17500 11880
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 17589 11883 17647 11889
rect 17589 11849 17601 11883
rect 17635 11880 17647 11883
rect 18782 11880 18788 11892
rect 17635 11852 18788 11880
rect 17635 11849 17647 11852
rect 17589 11843 17647 11849
rect 14608 11784 15148 11812
rect 14608 11772 14614 11784
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 9640 11716 9781 11744
rect 9640 11704 9646 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 11330 11744 11336 11756
rect 11291 11716 11336 11744
rect 9769 11707 9827 11713
rect 11330 11704 11336 11716
rect 11388 11704 11394 11756
rect 12713 11747 12771 11753
rect 12713 11713 12725 11747
rect 12759 11744 12771 11747
rect 13998 11744 14004 11756
rect 12759 11716 14004 11744
rect 12759 11713 12771 11716
rect 12713 11707 12771 11713
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11744 14243 11747
rect 14826 11744 14832 11756
rect 14231 11716 14832 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 14826 11704 14832 11716
rect 14884 11744 14890 11756
rect 15120 11753 15148 11784
rect 16114 11772 16120 11824
rect 16172 11812 16178 11824
rect 16482 11812 16488 11824
rect 16172 11784 16488 11812
rect 16172 11772 16178 11784
rect 16482 11772 16488 11784
rect 16540 11772 16546 11824
rect 16942 11772 16948 11824
rect 17000 11812 17006 11824
rect 17604 11812 17632 11843
rect 18782 11840 18788 11852
rect 18840 11840 18846 11892
rect 22462 11880 22468 11892
rect 22423 11852 22468 11880
rect 22462 11840 22468 11852
rect 22520 11880 22526 11892
rect 23017 11883 23075 11889
rect 23017 11880 23029 11883
rect 22520 11852 23029 11880
rect 22520 11840 22526 11852
rect 23017 11849 23029 11852
rect 23063 11849 23075 11883
rect 23017 11843 23075 11849
rect 17000 11784 17632 11812
rect 17000 11772 17006 11784
rect 14921 11747 14979 11753
rect 14921 11744 14933 11747
rect 14884 11716 14933 11744
rect 14884 11704 14890 11716
rect 14921 11713 14933 11716
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 15105 11747 15163 11753
rect 15105 11713 15117 11747
rect 15151 11713 15163 11747
rect 18598 11744 18604 11756
rect 18559 11716 18604 11744
rect 15105 11707 15163 11713
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 20898 11704 20904 11756
rect 20956 11744 20962 11756
rect 21085 11747 21143 11753
rect 21085 11744 21097 11747
rect 20956 11716 21097 11744
rect 20956 11704 20962 11716
rect 21085 11713 21097 11716
rect 21131 11713 21143 11747
rect 21085 11707 21143 11713
rect 23658 11704 23664 11756
rect 23716 11744 23722 11756
rect 24581 11747 24639 11753
rect 24581 11744 24593 11747
rect 23716 11716 24593 11744
rect 23716 11704 23722 11716
rect 24581 11713 24593 11716
rect 24627 11713 24639 11747
rect 25590 11744 25596 11756
rect 25551 11716 25596 11744
rect 24581 11707 24639 11713
rect 25590 11704 25596 11716
rect 25648 11704 25654 11756
rect 9122 11636 9128 11688
rect 9180 11676 9186 11688
rect 9677 11679 9735 11685
rect 9677 11676 9689 11679
rect 9180 11648 9689 11676
rect 9180 11636 9186 11648
rect 9677 11645 9689 11648
rect 9723 11645 9735 11679
rect 13906 11676 13912 11688
rect 13867 11648 13912 11676
rect 9677 11639 9735 11645
rect 13906 11636 13912 11648
rect 13964 11676 13970 11688
rect 15378 11685 15384 11688
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 13964 11648 14565 11676
rect 13964 11636 13970 11648
rect 14553 11645 14565 11648
rect 14599 11645 14611 11679
rect 15372 11676 15384 11685
rect 15339 11648 15384 11676
rect 14553 11639 14611 11645
rect 15372 11639 15384 11648
rect 15436 11676 15442 11688
rect 16114 11676 16120 11688
rect 15436 11648 16120 11676
rect 15378 11636 15384 11639
rect 15436 11636 15442 11648
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 16850 11636 16856 11688
rect 16908 11676 16914 11688
rect 17773 11679 17831 11685
rect 17773 11676 17785 11679
rect 16908 11648 17785 11676
rect 16908 11636 16914 11648
rect 17773 11645 17785 11648
rect 17819 11676 17831 11679
rect 17954 11676 17960 11688
rect 17819 11648 17960 11676
rect 17819 11645 17831 11648
rect 17773 11639 17831 11645
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 19150 11636 19156 11688
rect 19208 11676 19214 11688
rect 20533 11679 20591 11685
rect 20533 11676 20545 11679
rect 19208 11648 20545 11676
rect 19208 11636 19214 11648
rect 20533 11645 20545 11648
rect 20579 11645 20591 11679
rect 24118 11676 24124 11688
rect 20533 11639 20591 11645
rect 23860 11648 24124 11676
rect 9033 11611 9091 11617
rect 9033 11577 9045 11611
rect 9079 11608 9091 11611
rect 9079 11580 9628 11608
rect 9079 11577 9091 11580
rect 9033 11571 9091 11577
rect 9600 11552 9628 11580
rect 9950 11568 9956 11620
rect 10008 11608 10014 11620
rect 10597 11611 10655 11617
rect 10597 11608 10609 11611
rect 10008 11580 10609 11608
rect 10008 11568 10014 11580
rect 10597 11577 10609 11580
rect 10643 11608 10655 11611
rect 11149 11611 11207 11617
rect 11149 11608 11161 11611
rect 10643 11580 11161 11608
rect 10643 11577 10655 11580
rect 10597 11571 10655 11577
rect 11149 11577 11161 11580
rect 11195 11577 11207 11611
rect 11149 11571 11207 11577
rect 13449 11611 13507 11617
rect 13449 11577 13461 11611
rect 13495 11608 13507 11611
rect 13998 11608 14004 11620
rect 13495 11580 14004 11608
rect 13495 11577 13507 11580
rect 13449 11571 13507 11577
rect 13998 11568 14004 11580
rect 14056 11608 14062 11620
rect 14182 11608 14188 11620
rect 14056 11580 14188 11608
rect 14056 11568 14062 11580
rect 14182 11568 14188 11580
rect 14240 11568 14246 11620
rect 18690 11568 18696 11620
rect 18748 11608 18754 11620
rect 18868 11611 18926 11617
rect 18868 11608 18880 11611
rect 18748 11580 18880 11608
rect 18748 11568 18754 11580
rect 18868 11577 18880 11580
rect 18914 11608 18926 11611
rect 19242 11608 19248 11620
rect 18914 11580 19248 11608
rect 18914 11577 18926 11580
rect 18868 11571 18926 11577
rect 19242 11568 19248 11580
rect 19300 11568 19306 11620
rect 19886 11568 19892 11620
rect 19944 11608 19950 11620
rect 20901 11611 20959 11617
rect 20901 11608 20913 11611
rect 19944 11580 20913 11608
rect 19944 11568 19950 11580
rect 20901 11577 20913 11580
rect 20947 11608 20959 11611
rect 21330 11611 21388 11617
rect 21330 11608 21342 11611
rect 20947 11580 21342 11608
rect 20947 11577 20959 11580
rect 20901 11571 20959 11577
rect 21330 11577 21342 11580
rect 21376 11577 21388 11611
rect 21330 11571 21388 11577
rect 23106 11568 23112 11620
rect 23164 11608 23170 11620
rect 23860 11617 23888 11648
rect 24118 11636 24124 11648
rect 24176 11676 24182 11688
rect 24489 11679 24547 11685
rect 24489 11676 24501 11679
rect 24176 11648 24501 11676
rect 24176 11636 24182 11648
rect 24489 11645 24501 11648
rect 24535 11645 24547 11679
rect 24489 11639 24547 11645
rect 25038 11636 25044 11688
rect 25096 11676 25102 11688
rect 25409 11679 25467 11685
rect 25409 11676 25421 11679
rect 25096 11648 25421 11676
rect 25096 11636 25102 11648
rect 25409 11645 25421 11648
rect 25455 11645 25467 11679
rect 25409 11639 25467 11645
rect 23845 11611 23903 11617
rect 23845 11608 23857 11611
rect 23164 11580 23857 11608
rect 23164 11568 23170 11580
rect 23845 11577 23857 11580
rect 23891 11577 23903 11611
rect 23845 11571 23903 11577
rect 24210 11568 24216 11620
rect 24268 11608 24274 11620
rect 24397 11611 24455 11617
rect 24397 11608 24409 11611
rect 24268 11580 24409 11608
rect 24268 11568 24274 11580
rect 24397 11577 24409 11580
rect 24443 11608 24455 11611
rect 24762 11608 24768 11620
rect 24443 11580 24768 11608
rect 24443 11577 24455 11580
rect 24397 11571 24455 11577
rect 24762 11568 24768 11580
rect 24820 11568 24826 11620
rect 2038 11540 2044 11552
rect 1999 11512 2044 11540
rect 2038 11500 2044 11512
rect 2096 11500 2102 11552
rect 9214 11540 9220 11552
rect 9175 11512 9220 11540
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 9582 11540 9588 11552
rect 9543 11512 9588 11540
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 10778 11540 10784 11552
rect 10739 11512 10784 11540
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11241 11543 11299 11549
rect 11241 11540 11253 11543
rect 10928 11512 11253 11540
rect 10928 11500 10934 11512
rect 11241 11509 11253 11512
rect 11287 11540 11299 11543
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11287 11512 11805 11540
rect 11287 11509 11299 11512
rect 11241 11503 11299 11509
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 12802 11540 12808 11552
rect 12584 11512 12808 11540
rect 12584 11500 12590 11512
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 13081 11543 13139 11549
rect 13081 11509 13093 11543
rect 13127 11540 13139 11543
rect 14366 11540 14372 11552
rect 13127 11512 14372 11540
rect 13127 11509 13139 11512
rect 13081 11503 13139 11509
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 15838 11540 15844 11552
rect 15160 11512 15844 11540
rect 15160 11500 15166 11512
rect 15838 11500 15844 11512
rect 15896 11540 15902 11552
rect 16485 11543 16543 11549
rect 16485 11540 16497 11543
rect 15896 11512 16497 11540
rect 15896 11500 15902 11512
rect 16485 11509 16497 11512
rect 16531 11509 16543 11543
rect 16485 11503 16543 11509
rect 18509 11543 18567 11549
rect 18509 11509 18521 11543
rect 18555 11540 18567 11543
rect 19904 11540 19932 11568
rect 19981 11543 20039 11549
rect 19981 11540 19993 11543
rect 18555 11512 19993 11540
rect 18555 11509 18567 11512
rect 18509 11503 18567 11509
rect 19981 11509 19993 11512
rect 20027 11509 20039 11543
rect 19981 11503 20039 11509
rect 23477 11543 23535 11549
rect 23477 11509 23489 11543
rect 23523 11540 23535 11543
rect 23658 11540 23664 11552
rect 23523 11512 23664 11540
rect 23523 11509 23535 11512
rect 23477 11503 23535 11509
rect 23658 11500 23664 11512
rect 23716 11500 23722 11552
rect 24026 11540 24032 11552
rect 23987 11512 24032 11540
rect 24026 11500 24032 11512
rect 24084 11500 24090 11552
rect 25133 11543 25191 11549
rect 25133 11509 25145 11543
rect 25179 11540 25191 11543
rect 25314 11540 25320 11552
rect 25179 11512 25320 11540
rect 25179 11509 25191 11512
rect 25133 11503 25191 11509
rect 25314 11500 25320 11512
rect 25372 11500 25378 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 9217 11339 9275 11345
rect 9217 11336 9229 11339
rect 9180 11308 9229 11336
rect 9180 11296 9186 11308
rect 9217 11305 9229 11308
rect 9263 11305 9275 11339
rect 9950 11336 9956 11348
rect 9911 11308 9956 11336
rect 9217 11299 9275 11305
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10505 11339 10563 11345
rect 10505 11305 10517 11339
rect 10551 11336 10563 11339
rect 10778 11336 10784 11348
rect 10551 11308 10784 11336
rect 10551 11305 10563 11308
rect 10505 11299 10563 11305
rect 10778 11296 10784 11308
rect 10836 11336 10842 11348
rect 11333 11339 11391 11345
rect 11333 11336 11345 11339
rect 10836 11308 11345 11336
rect 10836 11296 10842 11308
rect 11333 11305 11345 11308
rect 11379 11305 11391 11339
rect 11333 11299 11391 11305
rect 12069 11339 12127 11345
rect 12069 11305 12081 11339
rect 12115 11336 12127 11339
rect 13170 11336 13176 11348
rect 12115 11308 13176 11336
rect 12115 11305 12127 11308
rect 12069 11299 12127 11305
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 14458 11336 14464 11348
rect 14419 11308 14464 11336
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 15102 11336 15108 11348
rect 15063 11308 15108 11336
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 15470 11336 15476 11348
rect 15431 11308 15476 11336
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 15838 11296 15844 11348
rect 15896 11336 15902 11348
rect 15933 11339 15991 11345
rect 15933 11336 15945 11339
rect 15896 11308 15945 11336
rect 15896 11296 15902 11308
rect 15933 11305 15945 11308
rect 15979 11336 15991 11339
rect 16206 11336 16212 11348
rect 15979 11308 16212 11336
rect 15979 11305 15991 11308
rect 15933 11299 15991 11305
rect 16206 11296 16212 11308
rect 16264 11296 16270 11348
rect 16574 11336 16580 11348
rect 16535 11308 16580 11336
rect 16574 11296 16580 11308
rect 16632 11336 16638 11348
rect 17405 11339 17463 11345
rect 17405 11336 17417 11339
rect 16632 11308 17417 11336
rect 16632 11296 16638 11308
rect 17405 11305 17417 11308
rect 17451 11305 17463 11339
rect 17405 11299 17463 11305
rect 17494 11296 17500 11348
rect 17552 11336 17558 11348
rect 18601 11339 18659 11345
rect 18601 11336 18613 11339
rect 17552 11308 18613 11336
rect 17552 11296 17558 11308
rect 18601 11305 18613 11308
rect 18647 11305 18659 11339
rect 18601 11299 18659 11305
rect 19518 11296 19524 11348
rect 19576 11336 19582 11348
rect 19613 11339 19671 11345
rect 19613 11336 19625 11339
rect 19576 11308 19625 11336
rect 19576 11296 19582 11308
rect 19613 11305 19625 11308
rect 19659 11305 19671 11339
rect 19978 11336 19984 11348
rect 19939 11308 19984 11336
rect 19613 11299 19671 11305
rect 19978 11296 19984 11308
rect 20036 11296 20042 11348
rect 20714 11296 20720 11348
rect 20772 11336 20778 11348
rect 20901 11339 20959 11345
rect 20901 11336 20913 11339
rect 20772 11308 20913 11336
rect 20772 11296 20778 11308
rect 20901 11305 20913 11308
rect 20947 11305 20959 11339
rect 20901 11299 20959 11305
rect 22097 11339 22155 11345
rect 22097 11305 22109 11339
rect 22143 11336 22155 11339
rect 22278 11336 22284 11348
rect 22143 11308 22284 11336
rect 22143 11305 22155 11308
rect 22097 11299 22155 11305
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 23201 11339 23259 11345
rect 23201 11305 23213 11339
rect 23247 11336 23259 11339
rect 23566 11336 23572 11348
rect 23247 11308 23572 11336
rect 23247 11305 23259 11308
rect 23201 11299 23259 11305
rect 23566 11296 23572 11308
rect 23624 11336 23630 11348
rect 23842 11336 23848 11348
rect 23624 11308 23848 11336
rect 23624 11296 23630 11308
rect 23842 11296 23848 11308
rect 23900 11296 23906 11348
rect 24765 11339 24823 11345
rect 24765 11305 24777 11339
rect 24811 11336 24823 11339
rect 25222 11336 25228 11348
rect 24811 11308 25228 11336
rect 24811 11305 24823 11308
rect 24765 11299 24823 11305
rect 25222 11296 25228 11308
rect 25280 11296 25286 11348
rect 25409 11339 25467 11345
rect 25409 11305 25421 11339
rect 25455 11336 25467 11339
rect 25774 11336 25780 11348
rect 25455 11308 25780 11336
rect 25455 11305 25467 11308
rect 25409 11299 25467 11305
rect 25774 11296 25780 11308
rect 25832 11296 25838 11348
rect 12342 11268 12348 11280
rect 12303 11240 12348 11268
rect 12342 11228 12348 11240
rect 12400 11228 12406 11280
rect 12618 11268 12624 11280
rect 12531 11240 12624 11268
rect 12618 11228 12624 11240
rect 12676 11268 12682 11280
rect 14550 11268 14556 11280
rect 12676 11240 14556 11268
rect 12676 11228 12682 11240
rect 14550 11228 14556 11240
rect 14608 11228 14614 11280
rect 17954 11228 17960 11280
rect 18012 11268 18018 11280
rect 18141 11271 18199 11277
rect 18141 11268 18153 11271
rect 18012 11240 18153 11268
rect 18012 11228 18018 11240
rect 18141 11237 18153 11240
rect 18187 11268 18199 11271
rect 19150 11268 19156 11280
rect 18187 11240 19156 11268
rect 18187 11237 18199 11240
rect 18141 11231 18199 11237
rect 19150 11228 19156 11240
rect 19208 11268 19214 11280
rect 19208 11240 19564 11268
rect 19208 11228 19214 11240
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 11425 11135 11483 11141
rect 11425 11132 11437 11135
rect 11112 11104 11437 11132
rect 11112 11092 11118 11104
rect 11425 11101 11437 11104
rect 11471 11101 11483 11135
rect 11606 11132 11612 11144
rect 11567 11104 11612 11132
rect 11425 11095 11483 11101
rect 10962 11064 10968 11076
rect 10923 11036 10968 11064
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 11440 11064 11468 11095
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 12536 11135 12594 11141
rect 12536 11101 12548 11135
rect 12582 11132 12594 11135
rect 12636 11132 12664 11228
rect 19536 11212 19564 11240
rect 21726 11228 21732 11280
rect 21784 11268 21790 11280
rect 22186 11268 22192 11280
rect 21784 11240 22192 11268
rect 21784 11228 21790 11240
rect 22186 11228 22192 11240
rect 22244 11268 22250 11280
rect 22465 11271 22523 11277
rect 22465 11268 22477 11271
rect 22244 11240 22477 11268
rect 22244 11228 22250 11240
rect 22465 11237 22477 11240
rect 22511 11237 22523 11271
rect 22465 11231 22523 11237
rect 12796 11203 12854 11209
rect 12796 11169 12808 11203
rect 12842 11200 12854 11203
rect 13078 11200 13084 11212
rect 12842 11172 13084 11200
rect 12842 11169 12854 11172
rect 12796 11163 12854 11169
rect 13078 11160 13084 11172
rect 13136 11160 13142 11212
rect 15841 11203 15899 11209
rect 15841 11169 15853 11203
rect 15887 11200 15899 11203
rect 16390 11200 16396 11212
rect 15887 11172 16396 11200
rect 15887 11169 15899 11172
rect 15841 11163 15899 11169
rect 16390 11160 16396 11172
rect 16448 11160 16454 11212
rect 18509 11203 18567 11209
rect 18509 11169 18521 11203
rect 18555 11200 18567 11203
rect 18782 11200 18788 11212
rect 18555 11172 18788 11200
rect 18555 11169 18567 11172
rect 18509 11163 18567 11169
rect 18782 11160 18788 11172
rect 18840 11160 18846 11212
rect 18874 11160 18880 11212
rect 18932 11200 18938 11212
rect 18969 11203 19027 11209
rect 18969 11200 18981 11203
rect 18932 11172 18981 11200
rect 18932 11160 18938 11172
rect 18969 11169 18981 11172
rect 19015 11169 19027 11203
rect 18969 11163 19027 11169
rect 19518 11160 19524 11212
rect 19576 11160 19582 11212
rect 20346 11160 20352 11212
rect 20404 11200 20410 11212
rect 20441 11203 20499 11209
rect 20441 11200 20453 11203
rect 20404 11172 20453 11200
rect 20404 11160 20410 11172
rect 20441 11169 20453 11172
rect 20487 11200 20499 11203
rect 20898 11200 20904 11212
rect 20487 11172 20904 11200
rect 20487 11169 20499 11172
rect 20441 11163 20499 11169
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 24026 11200 24032 11212
rect 23987 11172 24032 11200
rect 24026 11160 24032 11172
rect 24084 11160 24090 11212
rect 25130 11160 25136 11212
rect 25188 11200 25194 11212
rect 25225 11203 25283 11209
rect 25225 11200 25237 11203
rect 25188 11172 25237 11200
rect 25188 11160 25194 11172
rect 25225 11169 25237 11172
rect 25271 11169 25283 11203
rect 25225 11163 25283 11169
rect 16114 11132 16120 11144
rect 12582 11104 12664 11132
rect 16075 11104 16120 11132
rect 12582 11101 12594 11104
rect 12536 11095 12594 11101
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 17586 11132 17592 11144
rect 17547 11104 17592 11132
rect 17586 11092 17592 11104
rect 17644 11092 17650 11144
rect 18690 11092 18696 11144
rect 18748 11132 18754 11144
rect 19061 11135 19119 11141
rect 19061 11132 19073 11135
rect 18748 11104 19073 11132
rect 18748 11092 18754 11104
rect 19061 11101 19073 11104
rect 19107 11101 19119 11135
rect 19061 11095 19119 11101
rect 19153 11135 19211 11141
rect 19153 11101 19165 11135
rect 19199 11101 19211 11135
rect 22554 11132 22560 11144
rect 22515 11104 22560 11132
rect 19153 11095 19211 11101
rect 11440 11036 12480 11064
rect 12452 11008 12480 11036
rect 15746 11024 15752 11076
rect 15804 11064 15810 11076
rect 17037 11067 17095 11073
rect 17037 11064 17049 11067
rect 15804 11036 17049 11064
rect 15804 11024 15810 11036
rect 17037 11033 17049 11036
rect 17083 11033 17095 11067
rect 17037 11027 17095 11033
rect 17862 11024 17868 11076
rect 17920 11064 17926 11076
rect 19168 11064 19196 11095
rect 22554 11092 22560 11104
rect 22612 11092 22618 11144
rect 22646 11092 22652 11144
rect 22704 11132 22710 11144
rect 23566 11132 23572 11144
rect 22704 11104 22749 11132
rect 23479 11104 23572 11132
rect 22704 11092 22710 11104
rect 23566 11092 23572 11104
rect 23624 11132 23630 11144
rect 24121 11135 24179 11141
rect 24121 11132 24133 11135
rect 23624 11104 24133 11132
rect 23624 11092 23630 11104
rect 24121 11101 24133 11104
rect 24167 11101 24179 11135
rect 24121 11095 24179 11101
rect 24213 11135 24271 11141
rect 24213 11101 24225 11135
rect 24259 11101 24271 11135
rect 24213 11095 24271 11101
rect 17920 11036 19196 11064
rect 22005 11067 22063 11073
rect 17920 11024 17926 11036
rect 22005 11033 22017 11067
rect 22051 11064 22063 11067
rect 22664 11064 22692 11092
rect 22051 11036 22692 11064
rect 22051 11033 22063 11036
rect 22005 11027 22063 11033
rect 23750 11024 23756 11076
rect 23808 11064 23814 11076
rect 24228 11064 24256 11095
rect 23808 11036 24256 11064
rect 23808 11024 23814 11036
rect 10778 10996 10784 11008
rect 10739 10968 10784 10996
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 12434 10956 12440 11008
rect 12492 10956 12498 11008
rect 13909 10999 13967 11005
rect 13909 10965 13921 10999
rect 13955 10996 13967 10999
rect 14734 10996 14740 11008
rect 13955 10968 14740 10996
rect 13955 10965 13967 10968
rect 13909 10959 13967 10965
rect 14734 10956 14740 10968
rect 14792 10956 14798 11008
rect 16942 10996 16948 11008
rect 16855 10968 16948 10996
rect 16942 10956 16948 10968
rect 17000 10996 17006 11008
rect 17880 10996 17908 11024
rect 17000 10968 17908 10996
rect 21453 10999 21511 11005
rect 17000 10956 17006 10968
rect 21453 10965 21465 10999
rect 21499 10996 21511 10999
rect 21910 10996 21916 11008
rect 21499 10968 21916 10996
rect 21499 10965 21511 10968
rect 21453 10959 21511 10965
rect 21910 10956 21916 10968
rect 21968 10956 21974 11008
rect 23661 10999 23719 11005
rect 23661 10965 23673 10999
rect 23707 10996 23719 10999
rect 24210 10996 24216 11008
rect 23707 10968 24216 10996
rect 23707 10965 23719 10968
rect 23661 10959 23719 10965
rect 24210 10956 24216 10968
rect 24268 10956 24274 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 8938 10792 8944 10804
rect 8899 10764 8944 10792
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 12437 10795 12495 10801
rect 12437 10761 12449 10795
rect 12483 10792 12495 10795
rect 12526 10792 12532 10804
rect 12483 10764 12532 10792
rect 12483 10761 12495 10764
rect 12437 10755 12495 10761
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 13078 10752 13084 10804
rect 13136 10752 13142 10804
rect 15841 10795 15899 10801
rect 15841 10761 15853 10795
rect 15887 10792 15899 10795
rect 16114 10792 16120 10804
rect 15887 10764 16120 10792
rect 15887 10761 15899 10764
rect 15841 10755 15899 10761
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 16390 10792 16396 10804
rect 16351 10764 16396 10792
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 17862 10792 17868 10804
rect 17823 10764 17868 10792
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 18322 10792 18328 10804
rect 18283 10764 18328 10792
rect 18322 10752 18328 10764
rect 18380 10752 18386 10804
rect 21358 10792 21364 10804
rect 21319 10764 21364 10792
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 22186 10752 22192 10804
rect 22244 10792 22250 10804
rect 22373 10795 22431 10801
rect 22373 10792 22385 10795
rect 22244 10764 22385 10792
rect 22244 10752 22250 10764
rect 22373 10761 22385 10764
rect 22419 10761 22431 10795
rect 22373 10755 22431 10761
rect 23109 10795 23167 10801
rect 23109 10761 23121 10795
rect 23155 10792 23167 10795
rect 23658 10792 23664 10804
rect 23155 10764 23664 10792
rect 23155 10761 23167 10764
rect 23109 10755 23167 10761
rect 23658 10752 23664 10764
rect 23716 10792 23722 10804
rect 24118 10792 24124 10804
rect 23716 10764 24124 10792
rect 23716 10752 23722 10764
rect 24118 10752 24124 10764
rect 24176 10752 24182 10804
rect 25130 10752 25136 10804
rect 25188 10792 25194 10804
rect 25777 10795 25835 10801
rect 25777 10792 25789 10795
rect 25188 10764 25789 10792
rect 25188 10752 25194 10764
rect 25777 10761 25789 10764
rect 25823 10761 25835 10795
rect 25777 10755 25835 10761
rect 11517 10727 11575 10733
rect 11517 10693 11529 10727
rect 11563 10724 11575 10727
rect 11606 10724 11612 10736
rect 11563 10696 11612 10724
rect 11563 10693 11575 10696
rect 11517 10687 11575 10693
rect 11606 10684 11612 10696
rect 11664 10724 11670 10736
rect 12250 10724 12256 10736
rect 11664 10696 12256 10724
rect 11664 10684 11670 10696
rect 12250 10684 12256 10696
rect 12308 10724 12314 10736
rect 13096 10724 13124 10752
rect 12308 10696 13124 10724
rect 12308 10684 12314 10696
rect 9306 10656 9312 10668
rect 9267 10628 9312 10656
rect 9306 10616 9312 10628
rect 9364 10656 9370 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 9364 10628 9628 10656
rect 9364 10616 9370 10628
rect 8938 10548 8944 10600
rect 8996 10588 9002 10600
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 8996 10560 9505 10588
rect 8996 10548 9002 10560
rect 9493 10557 9505 10560
rect 9539 10557 9551 10591
rect 9600 10588 9628 10628
rect 11808 10628 13001 10656
rect 9749 10591 9807 10597
rect 9749 10588 9761 10591
rect 9600 10560 9761 10588
rect 9493 10551 9551 10557
rect 9749 10557 9761 10560
rect 9795 10588 9807 10591
rect 10042 10588 10048 10600
rect 9795 10560 10048 10588
rect 9795 10557 9807 10560
rect 9749 10551 9807 10557
rect 10042 10548 10048 10560
rect 10100 10548 10106 10600
rect 10778 10412 10784 10464
rect 10836 10452 10842 10464
rect 10873 10455 10931 10461
rect 10873 10452 10885 10455
rect 10836 10424 10885 10452
rect 10836 10412 10842 10424
rect 10873 10421 10885 10424
rect 10919 10452 10931 10455
rect 10962 10452 10968 10464
rect 10919 10424 10968 10452
rect 10919 10421 10931 10424
rect 10873 10415 10931 10421
rect 10962 10412 10968 10424
rect 11020 10452 11026 10464
rect 11330 10452 11336 10464
rect 11020 10424 11336 10452
rect 11020 10412 11026 10424
rect 11330 10412 11336 10424
rect 11388 10452 11394 10464
rect 11808 10461 11836 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 14369 10659 14427 10665
rect 14369 10625 14381 10659
rect 14415 10656 14427 10659
rect 16408 10656 16436 10752
rect 23842 10684 23848 10736
rect 23900 10684 23906 10736
rect 16945 10659 17003 10665
rect 16945 10656 16957 10659
rect 14415 10628 14596 10656
rect 16408 10628 16957 10656
rect 14415 10625 14427 10628
rect 14369 10619 14427 10625
rect 14458 10588 14464 10600
rect 14419 10560 14464 10588
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 14568 10588 14596 10628
rect 16945 10625 16957 10628
rect 16991 10625 17003 10659
rect 21913 10659 21971 10665
rect 21913 10656 21925 10659
rect 16945 10619 17003 10625
rect 20824 10628 21925 10656
rect 14734 10597 14740 10600
rect 14728 10588 14740 10597
rect 14568 10560 14740 10588
rect 14728 10551 14740 10560
rect 14734 10548 14740 10551
rect 14792 10548 14798 10600
rect 16114 10548 16120 10600
rect 16172 10588 16178 10600
rect 16761 10591 16819 10597
rect 16761 10588 16773 10591
rect 16172 10560 16773 10588
rect 16172 10548 16178 10560
rect 16761 10557 16773 10560
rect 16807 10588 16819 10591
rect 17405 10591 17463 10597
rect 17405 10588 17417 10591
rect 16807 10560 17417 10588
rect 16807 10557 16819 10560
rect 16761 10551 16819 10557
rect 17405 10557 17417 10560
rect 17451 10588 17463 10591
rect 17586 10588 17592 10600
rect 17451 10560 17592 10588
rect 17451 10557 17463 10560
rect 17405 10551 17463 10557
rect 17586 10548 17592 10560
rect 17644 10548 17650 10600
rect 18598 10548 18604 10600
rect 18656 10588 18662 10600
rect 18877 10591 18935 10597
rect 18877 10588 18889 10591
rect 18656 10560 18889 10588
rect 18656 10548 18662 10560
rect 18877 10557 18889 10560
rect 18923 10588 18935 10591
rect 19426 10588 19432 10600
rect 18923 10560 19432 10588
rect 18923 10557 18935 10560
rect 18877 10551 18935 10557
rect 19426 10548 19432 10560
rect 19484 10588 19490 10600
rect 20346 10588 20352 10600
rect 19484 10560 20352 10588
rect 19484 10548 19490 10560
rect 20346 10548 20352 10560
rect 20404 10548 20410 10600
rect 12805 10523 12863 10529
rect 12805 10489 12817 10523
rect 12851 10520 12863 10523
rect 12851 10492 13860 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 13832 10464 13860 10492
rect 15746 10480 15752 10532
rect 15804 10520 15810 10532
rect 16666 10520 16672 10532
rect 15804 10492 16672 10520
rect 15804 10480 15810 10492
rect 16666 10480 16672 10492
rect 16724 10480 16730 10532
rect 19058 10480 19064 10532
rect 19116 10529 19122 10532
rect 19116 10523 19180 10529
rect 19116 10489 19134 10523
rect 19168 10520 19180 10523
rect 20438 10520 20444 10532
rect 19168 10492 20444 10520
rect 19168 10489 19180 10492
rect 19116 10483 19180 10489
rect 19116 10480 19122 10483
rect 20438 10480 20444 10492
rect 20496 10520 20502 10532
rect 20824 10529 20852 10628
rect 21913 10625 21925 10628
rect 21959 10625 21971 10659
rect 21913 10619 21971 10625
rect 21269 10591 21327 10597
rect 21269 10557 21281 10591
rect 21315 10588 21327 10591
rect 21726 10588 21732 10600
rect 21315 10560 21732 10588
rect 21315 10557 21327 10560
rect 21269 10551 21327 10557
rect 21726 10548 21732 10560
rect 21784 10548 21790 10600
rect 23860 10597 23888 10684
rect 24118 10597 24124 10600
rect 23852 10591 23910 10597
rect 23852 10557 23864 10591
rect 23898 10557 23910 10591
rect 24112 10588 24124 10597
rect 24079 10560 24124 10588
rect 23852 10551 23910 10557
rect 24112 10551 24124 10560
rect 24118 10548 24124 10551
rect 24176 10548 24182 10600
rect 20809 10523 20867 10529
rect 20809 10520 20821 10523
rect 20496 10492 20821 10520
rect 20496 10480 20502 10492
rect 20809 10489 20821 10492
rect 20855 10489 20867 10523
rect 20809 10483 20867 10489
rect 23477 10523 23535 10529
rect 23477 10489 23489 10523
rect 23523 10520 23535 10523
rect 23750 10520 23756 10532
rect 23523 10492 23756 10520
rect 23523 10489 23535 10492
rect 23477 10483 23535 10489
rect 23750 10480 23756 10492
rect 23808 10520 23814 10532
rect 23808 10492 25268 10520
rect 23808 10480 23814 10492
rect 11793 10455 11851 10461
rect 11793 10452 11805 10455
rect 11388 10424 11805 10452
rect 11388 10412 11394 10424
rect 11793 10421 11805 10424
rect 11839 10421 11851 10455
rect 12894 10452 12900 10464
rect 12807 10424 12900 10452
rect 11793 10415 11851 10421
rect 12894 10412 12900 10424
rect 12952 10452 12958 10464
rect 13449 10455 13507 10461
rect 13449 10452 13461 10455
rect 12952 10424 13461 10452
rect 12952 10412 12958 10424
rect 13449 10421 13461 10424
rect 13495 10421 13507 10455
rect 13814 10452 13820 10464
rect 13775 10424 13820 10452
rect 13449 10415 13507 10421
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 18690 10452 18696 10464
rect 18651 10424 18696 10452
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 20257 10455 20315 10461
rect 20257 10452 20269 10455
rect 19392 10424 20269 10452
rect 19392 10412 19398 10424
rect 20257 10421 20269 10424
rect 20303 10421 20315 10455
rect 20257 10415 20315 10421
rect 21821 10455 21879 10461
rect 21821 10421 21833 10455
rect 21867 10452 21879 10455
rect 21910 10452 21916 10464
rect 21867 10424 21916 10452
rect 21867 10421 21879 10424
rect 21821 10415 21879 10421
rect 21910 10412 21916 10424
rect 21968 10412 21974 10464
rect 25240 10461 25268 10492
rect 25225 10455 25283 10461
rect 25225 10421 25237 10455
rect 25271 10421 25283 10455
rect 25225 10415 25283 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 10689 10251 10747 10257
rect 10689 10217 10701 10251
rect 10735 10248 10747 10251
rect 11054 10248 11060 10260
rect 10735 10220 11060 10248
rect 10735 10217 10747 10220
rect 10689 10211 10747 10217
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 12161 10251 12219 10257
rect 12161 10217 12173 10251
rect 12207 10248 12219 10251
rect 12250 10248 12256 10260
rect 12207 10220 12256 10248
rect 12207 10217 12219 10220
rect 12161 10211 12219 10217
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 12805 10251 12863 10257
rect 12805 10248 12817 10251
rect 12768 10220 12817 10248
rect 12768 10208 12774 10220
rect 12805 10217 12817 10220
rect 12851 10217 12863 10251
rect 12805 10211 12863 10217
rect 13265 10251 13323 10257
rect 13265 10217 13277 10251
rect 13311 10248 13323 10251
rect 13814 10248 13820 10260
rect 13311 10220 13820 10248
rect 13311 10217 13323 10220
rect 13265 10211 13323 10217
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 17129 10251 17187 10257
rect 17129 10217 17141 10251
rect 17175 10248 17187 10251
rect 17494 10248 17500 10260
rect 17175 10220 17500 10248
rect 17175 10217 17187 10220
rect 17129 10211 17187 10217
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 18598 10248 18604 10260
rect 18559 10220 18604 10248
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 18969 10251 19027 10257
rect 18969 10217 18981 10251
rect 19015 10248 19027 10251
rect 19058 10248 19064 10260
rect 19015 10220 19064 10248
rect 19015 10217 19027 10220
rect 18969 10211 19027 10217
rect 19058 10208 19064 10220
rect 19116 10208 19122 10260
rect 19334 10208 19340 10260
rect 19392 10248 19398 10260
rect 19705 10251 19763 10257
rect 19705 10248 19717 10251
rect 19392 10220 19717 10248
rect 19392 10208 19398 10220
rect 19705 10217 19717 10220
rect 19751 10248 19763 10251
rect 19978 10248 19984 10260
rect 19751 10220 19984 10248
rect 19751 10217 19763 10220
rect 19705 10211 19763 10217
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 20346 10248 20352 10260
rect 20307 10220 20352 10248
rect 20346 10208 20352 10220
rect 20404 10208 20410 10260
rect 22462 10248 22468 10260
rect 22423 10220 22468 10248
rect 22462 10208 22468 10220
rect 22520 10208 22526 10260
rect 23566 10248 23572 10260
rect 23527 10220 23572 10248
rect 23566 10208 23572 10220
rect 23624 10208 23630 10260
rect 24854 10208 24860 10260
rect 24912 10248 24918 10260
rect 25133 10251 25191 10257
rect 25133 10248 25145 10251
rect 24912 10220 25145 10248
rect 24912 10208 24918 10220
rect 25133 10217 25145 10220
rect 25179 10217 25191 10251
rect 25133 10211 25191 10217
rect 14366 10140 14372 10192
rect 14424 10180 14430 10192
rect 15105 10183 15163 10189
rect 15105 10180 15117 10183
rect 14424 10152 15117 10180
rect 14424 10140 14430 10152
rect 15105 10149 15117 10152
rect 15151 10180 15163 10183
rect 16117 10183 16175 10189
rect 16117 10180 16129 10183
rect 15151 10152 16129 10180
rect 15151 10149 15163 10152
rect 15105 10143 15163 10149
rect 16117 10149 16129 10152
rect 16163 10149 16175 10183
rect 16117 10143 16175 10149
rect 17402 10140 17408 10192
rect 17460 10180 17466 10192
rect 17681 10183 17739 10189
rect 17681 10180 17693 10183
rect 17460 10152 17693 10180
rect 17460 10140 17466 10152
rect 17681 10149 17693 10152
rect 17727 10149 17739 10183
rect 17681 10143 17739 10149
rect 23477 10183 23535 10189
rect 23477 10149 23489 10183
rect 23523 10180 23535 10183
rect 24026 10180 24032 10192
rect 23523 10152 24032 10180
rect 23523 10149 23535 10152
rect 23477 10143 23535 10149
rect 24026 10140 24032 10152
rect 24084 10140 24090 10192
rect 11054 10121 11060 10124
rect 11048 10112 11060 10121
rect 11015 10084 11060 10112
rect 11048 10075 11060 10084
rect 11054 10072 11060 10075
rect 11112 10072 11118 10124
rect 11790 10072 11796 10124
rect 11848 10112 11854 10124
rect 12618 10112 12624 10124
rect 11848 10084 12624 10112
rect 11848 10072 11854 10084
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 13630 10112 13636 10124
rect 13591 10084 13636 10112
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 16025 10115 16083 10121
rect 16025 10081 16037 10115
rect 16071 10112 16083 10115
rect 16669 10115 16727 10121
rect 16669 10112 16681 10115
rect 16071 10084 16681 10112
rect 16071 10081 16083 10084
rect 16025 10075 16083 10081
rect 16669 10081 16681 10084
rect 16715 10081 16727 10115
rect 16669 10075 16727 10081
rect 9950 10004 9956 10056
rect 10008 10044 10014 10056
rect 10781 10047 10839 10053
rect 10781 10044 10793 10047
rect 10008 10016 10793 10044
rect 10008 10004 10014 10016
rect 10781 10013 10793 10016
rect 10827 10013 10839 10047
rect 10781 10007 10839 10013
rect 13354 10004 13360 10056
rect 13412 10044 13418 10056
rect 13725 10047 13783 10053
rect 13725 10044 13737 10047
rect 13412 10016 13737 10044
rect 13412 10004 13418 10016
rect 13725 10013 13737 10016
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 13817 10047 13875 10053
rect 13817 10013 13829 10047
rect 13863 10013 13875 10047
rect 16206 10044 16212 10056
rect 16167 10016 16212 10044
rect 13817 10007 13875 10013
rect 13446 9936 13452 9988
rect 13504 9976 13510 9988
rect 13832 9976 13860 10007
rect 16206 10004 16212 10016
rect 16264 10004 16270 10056
rect 15838 9976 15844 9988
rect 13504 9948 13860 9976
rect 15488 9948 15844 9976
rect 13504 9936 13510 9948
rect 15488 9920 15516 9948
rect 15838 9936 15844 9948
rect 15896 9936 15902 9988
rect 16684 9976 16712 10075
rect 17310 10072 17316 10124
rect 17368 10112 17374 10124
rect 17589 10115 17647 10121
rect 17589 10112 17601 10115
rect 17368 10084 17601 10112
rect 17368 10072 17374 10084
rect 17589 10081 17601 10084
rect 17635 10081 17647 10115
rect 19610 10112 19616 10124
rect 19571 10084 19616 10112
rect 17589 10075 17647 10081
rect 19610 10072 19616 10084
rect 19668 10072 19674 10124
rect 21082 10072 21088 10124
rect 21140 10112 21146 10124
rect 21269 10115 21327 10121
rect 21269 10112 21281 10115
rect 21140 10084 21281 10112
rect 21140 10072 21146 10084
rect 21269 10081 21281 10084
rect 21315 10081 21327 10115
rect 21269 10075 21327 10081
rect 22097 10115 22155 10121
rect 22097 10081 22109 10115
rect 22143 10112 22155 10115
rect 23658 10112 23664 10124
rect 22143 10084 23664 10112
rect 22143 10081 22155 10084
rect 22097 10075 22155 10081
rect 23658 10072 23664 10084
rect 23716 10112 23722 10124
rect 23937 10115 23995 10121
rect 23937 10112 23949 10115
rect 23716 10084 23949 10112
rect 23716 10072 23722 10084
rect 23937 10081 23949 10084
rect 23983 10081 23995 10115
rect 23937 10075 23995 10081
rect 17770 10044 17776 10056
rect 17731 10016 17776 10044
rect 17770 10004 17776 10016
rect 17828 10004 17834 10056
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10044 19947 10047
rect 19978 10044 19984 10056
rect 19935 10016 19984 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 19978 10004 19984 10016
rect 20036 10004 20042 10056
rect 21358 10044 21364 10056
rect 21319 10016 21364 10044
rect 21358 10004 21364 10016
rect 21416 10004 21422 10056
rect 21450 10004 21456 10056
rect 21508 10044 21514 10056
rect 22557 10047 22615 10053
rect 21508 10016 21553 10044
rect 21508 10004 21514 10016
rect 22557 10013 22569 10047
rect 22603 10044 22615 10047
rect 23382 10044 23388 10056
rect 22603 10016 23388 10044
rect 22603 10013 22615 10016
rect 22557 10007 22615 10013
rect 23382 10004 23388 10016
rect 23440 10004 23446 10056
rect 23566 10004 23572 10056
rect 23624 10044 23630 10056
rect 24029 10047 24087 10053
rect 24029 10044 24041 10047
rect 23624 10016 24041 10044
rect 23624 10004 23630 10016
rect 24029 10013 24041 10016
rect 24075 10013 24087 10047
rect 24029 10007 24087 10013
rect 24118 10004 24124 10056
rect 24176 10044 24182 10056
rect 24176 10016 24221 10044
rect 24176 10004 24182 10016
rect 17221 9979 17279 9985
rect 17221 9976 17233 9979
rect 16684 9948 17233 9976
rect 17221 9945 17233 9948
rect 17267 9945 17279 9979
rect 17221 9939 17279 9945
rect 14458 9908 14464 9920
rect 14419 9880 14464 9908
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 15470 9908 15476 9920
rect 15431 9880 15476 9908
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 15657 9911 15715 9917
rect 15657 9877 15669 9911
rect 15703 9908 15715 9911
rect 16666 9908 16672 9920
rect 15703 9880 16672 9908
rect 15703 9877 15715 9880
rect 15657 9871 15715 9877
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 19242 9908 19248 9920
rect 19203 9880 19248 9908
rect 19242 9868 19248 9880
rect 19300 9868 19306 9920
rect 20901 9911 20959 9917
rect 20901 9877 20913 9911
rect 20947 9908 20959 9911
rect 21266 9908 21272 9920
rect 20947 9880 21272 9908
rect 20947 9877 20959 9880
rect 20901 9871 20959 9877
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 22186 9868 22192 9920
rect 22244 9908 22250 9920
rect 22554 9908 22560 9920
rect 22244 9880 22560 9908
rect 22244 9868 22250 9880
rect 22554 9868 22560 9880
rect 22612 9908 22618 9920
rect 23017 9911 23075 9917
rect 23017 9908 23029 9911
rect 22612 9880 23029 9908
rect 22612 9868 22618 9880
rect 23017 9877 23029 9880
rect 23063 9877 23075 9911
rect 23017 9871 23075 9877
rect 23750 9868 23756 9920
rect 23808 9908 23814 9920
rect 24581 9911 24639 9917
rect 24581 9908 24593 9911
rect 23808 9880 24593 9908
rect 23808 9868 23814 9880
rect 24581 9877 24593 9880
rect 24627 9877 24639 9911
rect 24581 9871 24639 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 9950 9704 9956 9716
rect 9911 9676 9956 9704
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 10229 9707 10287 9713
rect 10229 9704 10241 9707
rect 10100 9676 10241 9704
rect 10100 9664 10106 9676
rect 10229 9673 10241 9676
rect 10275 9673 10287 9707
rect 10229 9667 10287 9673
rect 12805 9707 12863 9713
rect 12805 9673 12817 9707
rect 12851 9704 12863 9707
rect 12894 9704 12900 9716
rect 12851 9676 12900 9704
rect 12851 9673 12863 9676
rect 12805 9667 12863 9673
rect 10244 9568 10272 9667
rect 12894 9664 12900 9676
rect 12952 9664 12958 9716
rect 14366 9704 14372 9716
rect 14327 9676 14372 9704
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 17310 9704 17316 9716
rect 17271 9676 17316 9704
rect 17310 9664 17316 9676
rect 17368 9664 17374 9716
rect 17402 9664 17408 9716
rect 17460 9704 17466 9716
rect 17589 9707 17647 9713
rect 17589 9704 17601 9707
rect 17460 9676 17601 9704
rect 17460 9664 17466 9676
rect 17589 9673 17601 9676
rect 17635 9673 17647 9707
rect 19610 9704 19616 9716
rect 17589 9667 17647 9673
rect 19352 9676 19616 9704
rect 10781 9639 10839 9645
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 10870 9636 10876 9648
rect 10827 9608 10876 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 10870 9596 10876 9608
rect 10928 9596 10934 9648
rect 11790 9636 11796 9648
rect 11751 9608 11796 9636
rect 11790 9596 11796 9608
rect 11848 9596 11854 9648
rect 13909 9639 13967 9645
rect 12176 9608 13492 9636
rect 12176 9577 12204 9608
rect 13464 9580 13492 9608
rect 13909 9605 13921 9639
rect 13955 9636 13967 9639
rect 13998 9636 14004 9648
rect 13955 9608 14004 9636
rect 13955 9605 13967 9608
rect 13909 9599 13967 9605
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 15841 9639 15899 9645
rect 15841 9605 15853 9639
rect 15887 9636 15899 9639
rect 15930 9636 15936 9648
rect 15887 9608 15936 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 15930 9596 15936 9608
rect 15988 9636 15994 9648
rect 18969 9639 19027 9645
rect 18969 9636 18981 9639
rect 15988 9608 16436 9636
rect 15988 9596 15994 9608
rect 11333 9571 11391 9577
rect 11333 9568 11345 9571
rect 10244 9540 11345 9568
rect 11333 9537 11345 9540
rect 11379 9568 11391 9571
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 11379 9540 12173 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 12161 9537 12173 9540
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 13265 9571 13323 9577
rect 13265 9568 13277 9571
rect 12768 9540 13277 9568
rect 12768 9528 12774 9540
rect 13265 9537 13277 9540
rect 13311 9537 13323 9571
rect 13446 9568 13452 9580
rect 13407 9540 13452 9568
rect 13265 9531 13323 9537
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 14458 9528 14464 9580
rect 14516 9568 14522 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14516 9540 15025 9568
rect 14516 9528 14522 9540
rect 15013 9537 15025 9540
rect 15059 9568 15071 9571
rect 15654 9568 15660 9580
rect 15059 9540 15660 9568
rect 15059 9537 15071 9540
rect 15013 9531 15071 9537
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 16408 9577 16436 9608
rect 18432 9608 18981 9636
rect 18432 9577 18460 9608
rect 18969 9605 18981 9608
rect 19015 9636 19027 9639
rect 19352 9636 19380 9676
rect 19610 9664 19616 9676
rect 19668 9664 19674 9716
rect 20162 9664 20168 9716
rect 20220 9704 20226 9716
rect 20346 9704 20352 9716
rect 20220 9676 20352 9704
rect 20220 9664 20226 9676
rect 20346 9664 20352 9676
rect 20404 9664 20410 9716
rect 22002 9636 22008 9648
rect 19015 9608 19380 9636
rect 21963 9608 22008 9636
rect 19015 9605 19027 9608
rect 18969 9599 19027 9605
rect 22002 9596 22008 9608
rect 22060 9596 22066 9648
rect 23106 9636 23112 9648
rect 22388 9608 23112 9636
rect 16393 9571 16451 9577
rect 16393 9537 16405 9571
rect 16439 9537 16451 9571
rect 16393 9531 16451 9537
rect 16485 9571 16543 9577
rect 16485 9537 16497 9571
rect 16531 9537 16543 9571
rect 16485 9531 16543 9537
rect 18417 9571 18475 9577
rect 18417 9537 18429 9571
rect 18463 9537 18475 9571
rect 19334 9568 19340 9580
rect 19295 9540 19340 9568
rect 18417 9531 18475 9537
rect 10778 9460 10784 9512
rect 10836 9500 10842 9512
rect 11238 9500 11244 9512
rect 10836 9472 11244 9500
rect 10836 9460 10842 9472
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 14277 9503 14335 9509
rect 14277 9469 14289 9503
rect 14323 9500 14335 9503
rect 14734 9500 14740 9512
rect 14323 9472 14740 9500
rect 14323 9469 14335 9472
rect 14277 9463 14335 9469
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 14826 9460 14832 9512
rect 14884 9500 14890 9512
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 14884 9472 15393 9500
rect 14884 9460 14890 9472
rect 15381 9469 15393 9472
rect 15427 9500 15439 9503
rect 16206 9500 16212 9512
rect 15427 9472 16212 9500
rect 15427 9469 15439 9472
rect 15381 9463 15439 9469
rect 16206 9460 16212 9472
rect 16264 9500 16270 9512
rect 16500 9500 16528 9531
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 19484 9540 19529 9568
rect 19484 9528 19490 9540
rect 22388 9509 22416 9608
rect 23106 9596 23112 9608
rect 23164 9596 23170 9648
rect 22462 9528 22468 9580
rect 22520 9568 22526 9580
rect 22557 9571 22615 9577
rect 22557 9568 22569 9571
rect 22520 9540 22569 9568
rect 22520 9528 22526 9540
rect 22557 9537 22569 9540
rect 22603 9537 22615 9571
rect 23750 9568 23756 9580
rect 23711 9540 23756 9568
rect 22557 9531 22615 9537
rect 23750 9528 23756 9540
rect 23808 9528 23814 9580
rect 16264 9472 16528 9500
rect 21913 9503 21971 9509
rect 16264 9460 16270 9472
rect 21913 9469 21925 9503
rect 21959 9500 21971 9503
rect 22373 9503 22431 9509
rect 22373 9500 22385 9503
rect 21959 9472 22385 9500
rect 21959 9469 21971 9472
rect 21913 9463 21971 9469
rect 22373 9469 22385 9472
rect 22419 9469 22431 9503
rect 23658 9500 23664 9512
rect 22373 9463 22431 9469
rect 22480 9472 23664 9500
rect 12713 9435 12771 9441
rect 12713 9401 12725 9435
rect 12759 9432 12771 9435
rect 13170 9432 13176 9444
rect 12759 9404 13176 9432
rect 12759 9401 12771 9404
rect 12713 9395 12771 9401
rect 13170 9392 13176 9404
rect 13228 9392 13234 9444
rect 14366 9392 14372 9444
rect 14424 9432 14430 9444
rect 19696 9435 19754 9441
rect 14424 9404 14872 9432
rect 14424 9392 14430 9404
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 10597 9367 10655 9373
rect 10597 9364 10609 9367
rect 9732 9336 10609 9364
rect 9732 9324 9738 9336
rect 10597 9333 10609 9336
rect 10643 9364 10655 9367
rect 11149 9367 11207 9373
rect 11149 9364 11161 9367
rect 10643 9336 11161 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 11149 9333 11161 9336
rect 11195 9364 11207 9367
rect 12158 9364 12164 9376
rect 11195 9336 12164 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 14844 9373 14872 9404
rect 19696 9401 19708 9435
rect 19742 9432 19754 9435
rect 20070 9432 20076 9444
rect 19742 9404 20076 9432
rect 19742 9401 19754 9404
rect 19696 9395 19754 9401
rect 20070 9392 20076 9404
rect 20128 9392 20134 9444
rect 21358 9432 21364 9444
rect 21319 9404 21364 9432
rect 21358 9392 21364 9404
rect 21416 9392 21422 9444
rect 22480 9441 22508 9472
rect 23658 9460 23664 9472
rect 23716 9460 23722 9512
rect 22465 9435 22523 9441
rect 22465 9401 22477 9435
rect 22511 9401 22523 9435
rect 23566 9432 23572 9444
rect 22465 9395 22523 9401
rect 23032 9404 23572 9432
rect 23032 9376 23060 9404
rect 23566 9392 23572 9404
rect 23624 9392 23630 9444
rect 23934 9392 23940 9444
rect 23992 9441 23998 9444
rect 23992 9435 24056 9441
rect 23992 9401 24010 9435
rect 24044 9401 24056 9435
rect 23992 9395 24056 9401
rect 23992 9392 23998 9395
rect 14829 9367 14887 9373
rect 14829 9333 14841 9367
rect 14875 9333 14887 9367
rect 15930 9364 15936 9376
rect 15891 9336 15936 9364
rect 14829 9327 14887 9333
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 16022 9324 16028 9376
rect 16080 9364 16086 9376
rect 16301 9367 16359 9373
rect 16301 9364 16313 9367
rect 16080 9336 16313 9364
rect 16080 9324 16086 9336
rect 16301 9333 16313 9336
rect 16347 9333 16359 9367
rect 16301 9327 16359 9333
rect 17770 9324 17776 9376
rect 17828 9364 17834 9376
rect 18322 9364 18328 9376
rect 17828 9336 18328 9364
rect 17828 9324 17834 9336
rect 18322 9324 18328 9336
rect 18380 9324 18386 9376
rect 19978 9324 19984 9376
rect 20036 9364 20042 9376
rect 20806 9364 20812 9376
rect 20036 9336 20812 9364
rect 20036 9324 20042 9336
rect 20806 9324 20812 9336
rect 20864 9324 20870 9376
rect 23014 9364 23020 9376
rect 22975 9336 23020 9364
rect 23014 9324 23020 9336
rect 23072 9324 23078 9376
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 23658 9364 23664 9376
rect 23523 9336 23664 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 23658 9324 23664 9336
rect 23716 9324 23722 9376
rect 24118 9324 24124 9376
rect 24176 9364 24182 9376
rect 25133 9367 25191 9373
rect 25133 9364 25145 9367
rect 24176 9336 25145 9364
rect 24176 9324 24182 9336
rect 25133 9333 25145 9336
rect 25179 9333 25191 9367
rect 25133 9327 25191 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 11054 9120 11060 9172
rect 11112 9160 11118 9172
rect 11149 9163 11207 9169
rect 11149 9160 11161 9163
rect 11112 9132 11161 9160
rect 11112 9120 11118 9132
rect 11149 9129 11161 9132
rect 11195 9129 11207 9163
rect 13354 9160 13360 9172
rect 13315 9132 13360 9160
rect 11149 9123 11207 9129
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 13633 9163 13691 9169
rect 13633 9160 13645 9163
rect 13504 9132 13645 9160
rect 13504 9120 13510 9132
rect 13633 9129 13645 9132
rect 13679 9129 13691 9163
rect 13633 9123 13691 9129
rect 14093 9163 14151 9169
rect 14093 9129 14105 9163
rect 14139 9160 14151 9163
rect 14550 9160 14556 9172
rect 14139 9132 14556 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 15289 9163 15347 9169
rect 15289 9129 15301 9163
rect 15335 9160 15347 9163
rect 16022 9160 16028 9172
rect 15335 9132 16028 9160
rect 15335 9129 15347 9132
rect 15289 9123 15347 9129
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 16206 9120 16212 9172
rect 16264 9160 16270 9172
rect 17681 9163 17739 9169
rect 17681 9160 17693 9163
rect 16264 9132 17693 9160
rect 16264 9120 16270 9132
rect 17681 9129 17693 9132
rect 17727 9129 17739 9163
rect 17681 9123 17739 9129
rect 18785 9163 18843 9169
rect 18785 9129 18797 9163
rect 18831 9160 18843 9163
rect 19242 9160 19248 9172
rect 18831 9132 19248 9160
rect 18831 9129 18843 9132
rect 18785 9123 18843 9129
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 20349 9163 20407 9169
rect 20349 9129 20361 9163
rect 20395 9160 20407 9163
rect 21450 9160 21456 9172
rect 20395 9132 21456 9160
rect 20395 9129 20407 9132
rect 20349 9123 20407 9129
rect 14366 9092 14372 9104
rect 14327 9064 14372 9092
rect 14366 9052 14372 9064
rect 14424 9052 14430 9104
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 11330 9024 11336 9036
rect 10008 8996 11336 9024
rect 10008 8984 10014 8996
rect 11330 8984 11336 8996
rect 11388 8984 11394 9036
rect 11422 8984 11428 9036
rect 11480 9024 11486 9036
rect 11589 9027 11647 9033
rect 11589 9024 11601 9027
rect 11480 8996 11601 9024
rect 11480 8984 11486 8996
rect 11589 8993 11601 8996
rect 11635 8993 11647 9027
rect 14568 9024 14596 9120
rect 15654 9052 15660 9104
rect 15712 9092 15718 9104
rect 16568 9095 16626 9101
rect 16568 9092 16580 9095
rect 15712 9064 16580 9092
rect 15712 9052 15718 9064
rect 16568 9061 16580 9064
rect 16614 9092 16626 9095
rect 17770 9092 17776 9104
rect 16614 9064 17776 9092
rect 16614 9061 16626 9064
rect 16568 9055 16626 9061
rect 17770 9052 17776 9064
rect 17828 9052 17834 9104
rect 19153 9095 19211 9101
rect 19153 9061 19165 9095
rect 19199 9092 19211 9095
rect 19978 9092 19984 9104
rect 19199 9064 19984 9092
rect 19199 9061 19211 9064
rect 19153 9055 19211 9061
rect 19978 9052 19984 9064
rect 20036 9052 20042 9104
rect 16301 9027 16359 9033
rect 16301 9024 16313 9027
rect 14568 8996 16313 9024
rect 11589 8987 11647 8993
rect 16301 8993 16313 8996
rect 16347 9024 16359 9027
rect 17586 9024 17592 9036
rect 16347 8996 17592 9024
rect 16347 8993 16359 8996
rect 16301 8987 16359 8993
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 19613 9027 19671 9033
rect 19613 8993 19625 9027
rect 19659 9024 19671 9027
rect 20162 9024 20168 9036
rect 19659 8996 20168 9024
rect 19659 8993 19671 8996
rect 19613 8987 19671 8993
rect 20162 8984 20168 8996
rect 20220 8984 20226 9036
rect 10778 8956 10784 8968
rect 10739 8928 10784 8956
rect 10778 8916 10784 8928
rect 10836 8916 10842 8968
rect 19334 8916 19340 8968
rect 19392 8956 19398 8968
rect 19705 8959 19763 8965
rect 19705 8956 19717 8959
rect 19392 8928 19717 8956
rect 19392 8916 19398 8928
rect 19705 8925 19717 8928
rect 19751 8925 19763 8959
rect 19705 8919 19763 8925
rect 19889 8959 19947 8965
rect 19889 8925 19901 8959
rect 19935 8956 19947 8959
rect 20070 8956 20076 8968
rect 19935 8928 20076 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 20070 8916 20076 8928
rect 20128 8956 20134 8968
rect 20364 8956 20392 9123
rect 21450 9120 21456 9132
rect 21508 9120 21514 9172
rect 24118 9160 24124 9172
rect 24079 9132 24124 9160
rect 24118 9120 24124 9132
rect 24176 9120 24182 9172
rect 21082 9092 21088 9104
rect 21043 9064 21088 9092
rect 21082 9052 21088 9064
rect 21140 9052 21146 9104
rect 24949 9095 25007 9101
rect 24949 9061 24961 9095
rect 24995 9092 25007 9095
rect 25038 9092 25044 9104
rect 24995 9064 25044 9092
rect 24995 9061 25007 9064
rect 24949 9055 25007 9061
rect 25038 9052 25044 9064
rect 25096 9052 25102 9104
rect 22094 9033 22100 9036
rect 22088 8987 22100 9033
rect 22152 9024 22158 9036
rect 22152 8996 22188 9024
rect 22094 8984 22100 8987
rect 22152 8984 22158 8996
rect 24854 8984 24860 9036
rect 24912 9024 24918 9036
rect 24912 8996 25176 9024
rect 24912 8984 24918 8996
rect 20128 8928 20392 8956
rect 20128 8916 20134 8928
rect 21542 8916 21548 8968
rect 21600 8956 21606 8968
rect 21821 8959 21879 8965
rect 21821 8956 21833 8959
rect 21600 8928 21833 8956
rect 21600 8916 21606 8928
rect 21821 8925 21833 8928
rect 21867 8925 21879 8959
rect 21821 8919 21879 8925
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 23934 8956 23940 8968
rect 23891 8928 23940 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 23934 8916 23940 8928
rect 23992 8956 23998 8968
rect 24762 8956 24768 8968
rect 23992 8928 24768 8956
rect 23992 8916 23998 8928
rect 24762 8916 24768 8928
rect 24820 8916 24826 8968
rect 25148 8965 25176 8996
rect 25041 8959 25099 8965
rect 25041 8925 25053 8959
rect 25087 8925 25099 8959
rect 25041 8919 25099 8925
rect 25133 8959 25191 8965
rect 25133 8925 25145 8959
rect 25179 8925 25191 8959
rect 25133 8919 25191 8925
rect 25056 8888 25084 8919
rect 25314 8888 25320 8900
rect 25056 8860 25320 8888
rect 25314 8848 25320 8860
rect 25372 8888 25378 8900
rect 25682 8888 25688 8900
rect 25372 8860 25688 8888
rect 25372 8848 25378 8860
rect 25682 8848 25688 8860
rect 25740 8848 25746 8900
rect 12710 8820 12716 8832
rect 12671 8792 12716 8820
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 14826 8780 14832 8832
rect 14884 8820 14890 8832
rect 15013 8823 15071 8829
rect 15013 8820 15025 8823
rect 14884 8792 15025 8820
rect 14884 8780 14890 8792
rect 15013 8789 15025 8792
rect 15059 8789 15071 8823
rect 15013 8783 15071 8789
rect 19150 8780 19156 8832
rect 19208 8820 19214 8832
rect 19245 8823 19303 8829
rect 19245 8820 19257 8823
rect 19208 8792 19257 8820
rect 19208 8780 19214 8792
rect 19245 8789 19257 8792
rect 19291 8789 19303 8823
rect 19245 8783 19303 8789
rect 20530 8780 20536 8832
rect 20588 8820 20594 8832
rect 20625 8823 20683 8829
rect 20625 8820 20637 8823
rect 20588 8792 20637 8820
rect 20588 8780 20594 8792
rect 20625 8789 20637 8792
rect 20671 8789 20683 8823
rect 20625 8783 20683 8789
rect 23201 8823 23259 8829
rect 23201 8789 23213 8823
rect 23247 8820 23259 8823
rect 23382 8820 23388 8832
rect 23247 8792 23388 8820
rect 23247 8789 23259 8792
rect 23201 8783 23259 8789
rect 23382 8780 23388 8792
rect 23440 8780 23446 8832
rect 24118 8780 24124 8832
rect 24176 8820 24182 8832
rect 24581 8823 24639 8829
rect 24581 8820 24593 8823
rect 24176 8792 24593 8820
rect 24176 8780 24182 8792
rect 24581 8789 24593 8792
rect 24627 8789 24639 8823
rect 24581 8783 24639 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 11422 8616 11428 8628
rect 11383 8588 11428 8616
rect 11422 8576 11428 8588
rect 11480 8576 11486 8628
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 16209 8619 16267 8625
rect 16209 8616 16221 8619
rect 14700 8588 16221 8616
rect 14700 8576 14706 8588
rect 16209 8585 16221 8588
rect 16255 8585 16267 8619
rect 17586 8616 17592 8628
rect 17547 8588 17592 8616
rect 16209 8579 16267 8585
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 21821 8619 21879 8625
rect 21821 8616 21833 8619
rect 19444 8588 21833 8616
rect 11330 8508 11336 8560
rect 11388 8548 11394 8560
rect 11701 8551 11759 8557
rect 11701 8548 11713 8551
rect 11388 8520 11713 8548
rect 11388 8508 11394 8520
rect 11701 8517 11713 8520
rect 11747 8517 11759 8551
rect 11701 8511 11759 8517
rect 11716 8412 11744 8511
rect 14734 8508 14740 8560
rect 14792 8548 14798 8560
rect 15105 8551 15163 8557
rect 15105 8548 15117 8551
rect 14792 8520 15117 8548
rect 14792 8508 14798 8520
rect 15105 8517 15117 8520
rect 15151 8548 15163 8551
rect 16117 8551 16175 8557
rect 16117 8548 16129 8551
rect 15151 8520 16129 8548
rect 15151 8517 15163 8520
rect 15105 8511 15163 8517
rect 16117 8517 16129 8520
rect 16163 8548 16175 8551
rect 18874 8548 18880 8560
rect 16163 8520 16804 8548
rect 18835 8520 18880 8548
rect 16163 8517 16175 8520
rect 16117 8511 16175 8517
rect 15654 8480 15660 8492
rect 15615 8452 15660 8480
rect 15654 8440 15660 8452
rect 15712 8440 15718 8492
rect 16666 8480 16672 8492
rect 16627 8452 16672 8480
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 16776 8489 16804 8520
rect 18874 8508 18880 8520
rect 18932 8508 18938 8560
rect 19444 8489 19472 8588
rect 21821 8585 21833 8588
rect 21867 8616 21879 8619
rect 22094 8616 22100 8628
rect 21867 8588 22100 8616
rect 21867 8585 21879 8588
rect 21821 8579 21879 8585
rect 22094 8576 22100 8588
rect 22152 8616 22158 8628
rect 22373 8619 22431 8625
rect 22373 8616 22385 8619
rect 22152 8588 22385 8616
rect 22152 8576 22158 8588
rect 22373 8585 22385 8588
rect 22419 8585 22431 8619
rect 22373 8579 22431 8585
rect 24762 8508 24768 8560
rect 24820 8548 24826 8560
rect 25041 8551 25099 8557
rect 25041 8548 25053 8551
rect 24820 8520 25053 8548
rect 24820 8508 24826 8520
rect 25041 8517 25053 8520
rect 25087 8517 25099 8551
rect 25041 8511 25099 8517
rect 16761 8483 16819 8489
rect 16761 8449 16773 8483
rect 16807 8449 16819 8483
rect 16761 8443 16819 8449
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8480 18843 8483
rect 19429 8483 19487 8489
rect 19429 8480 19441 8483
rect 18831 8452 19441 8480
rect 18831 8449 18843 8452
rect 18785 8443 18843 8449
rect 19429 8449 19441 8452
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 11716 8384 13737 8412
rect 13556 8288 13584 8384
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 15930 8372 15936 8424
rect 15988 8412 15994 8424
rect 16577 8415 16635 8421
rect 16577 8412 16589 8415
rect 15988 8384 16589 8412
rect 15988 8372 15994 8384
rect 16577 8381 16589 8384
rect 16623 8412 16635 8415
rect 17221 8415 17279 8421
rect 17221 8412 17233 8415
rect 16623 8384 17233 8412
rect 16623 8381 16635 8384
rect 16577 8375 16635 8381
rect 17221 8381 17233 8384
rect 17267 8381 17279 8415
rect 19242 8412 19248 8424
rect 19203 8384 19248 8412
rect 17221 8375 17279 8381
rect 19242 8372 19248 8384
rect 19300 8372 19306 8424
rect 19981 8415 20039 8421
rect 19981 8381 19993 8415
rect 20027 8412 20039 8415
rect 20162 8412 20168 8424
rect 20027 8384 20168 8412
rect 20027 8381 20039 8384
rect 19981 8375 20039 8381
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 20441 8415 20499 8421
rect 20441 8381 20453 8415
rect 20487 8412 20499 8415
rect 20530 8412 20536 8424
rect 20487 8384 20536 8412
rect 20487 8381 20499 8384
rect 20441 8375 20499 8381
rect 20530 8372 20536 8384
rect 20588 8412 20594 8424
rect 21542 8412 21548 8424
rect 20588 8384 21548 8412
rect 20588 8372 20594 8384
rect 21542 8372 21548 8384
rect 21600 8372 21606 8424
rect 23109 8415 23167 8421
rect 23109 8381 23121 8415
rect 23155 8412 23167 8415
rect 23290 8412 23296 8424
rect 23155 8384 23296 8412
rect 23155 8381 23167 8384
rect 23109 8375 23167 8381
rect 23290 8372 23296 8384
rect 23348 8412 23354 8424
rect 23661 8415 23719 8421
rect 23661 8412 23673 8415
rect 23348 8384 23673 8412
rect 23348 8372 23354 8384
rect 23661 8381 23673 8384
rect 23707 8412 23719 8415
rect 23750 8412 23756 8424
rect 23707 8384 23756 8412
rect 23707 8381 23719 8384
rect 23661 8375 23719 8381
rect 23750 8372 23756 8384
rect 23808 8372 23814 8424
rect 24854 8372 24860 8424
rect 24912 8412 24918 8424
rect 25961 8415 26019 8421
rect 25961 8412 25973 8415
rect 24912 8384 25973 8412
rect 24912 8372 24918 8384
rect 25961 8381 25973 8384
rect 26007 8381 26019 8415
rect 25961 8375 26019 8381
rect 13633 8347 13691 8353
rect 13633 8313 13645 8347
rect 13679 8344 13691 8347
rect 13970 8347 14028 8353
rect 13970 8344 13982 8347
rect 13679 8316 13982 8344
rect 13679 8313 13691 8316
rect 13633 8307 13691 8313
rect 13970 8313 13982 8316
rect 14016 8344 14028 8347
rect 14826 8344 14832 8356
rect 14016 8316 14832 8344
rect 14016 8313 14028 8316
rect 13970 8307 14028 8313
rect 14826 8304 14832 8316
rect 14884 8304 14890 8356
rect 18417 8347 18475 8353
rect 18417 8313 18429 8347
rect 18463 8344 18475 8347
rect 20070 8344 20076 8356
rect 18463 8316 20076 8344
rect 18463 8313 18475 8316
rect 18417 8307 18475 8313
rect 20070 8304 20076 8316
rect 20128 8304 20134 8356
rect 20349 8347 20407 8353
rect 20349 8313 20361 8347
rect 20395 8344 20407 8347
rect 20708 8347 20766 8353
rect 20708 8344 20720 8347
rect 20395 8316 20720 8344
rect 20395 8313 20407 8316
rect 20349 8307 20407 8313
rect 20708 8313 20720 8316
rect 20754 8344 20766 8347
rect 20806 8344 20812 8356
rect 20754 8316 20812 8344
rect 20754 8313 20766 8316
rect 20708 8307 20766 8313
rect 20806 8304 20812 8316
rect 20864 8344 20870 8356
rect 21634 8344 21640 8356
rect 20864 8316 21640 8344
rect 20864 8304 20870 8316
rect 21634 8304 21640 8316
rect 21692 8304 21698 8356
rect 23477 8347 23535 8353
rect 23477 8313 23489 8347
rect 23523 8344 23535 8347
rect 23928 8347 23986 8353
rect 23928 8344 23940 8347
rect 23523 8316 23940 8344
rect 23523 8313 23535 8316
rect 23477 8307 23535 8313
rect 23928 8313 23940 8316
rect 23974 8344 23986 8347
rect 24210 8344 24216 8356
rect 23974 8316 24216 8344
rect 23974 8313 23986 8316
rect 23928 8307 23986 8313
rect 24210 8304 24216 8316
rect 24268 8304 24274 8356
rect 25682 8344 25688 8356
rect 25643 8316 25688 8344
rect 25682 8304 25688 8316
rect 25740 8304 25746 8356
rect 13265 8279 13323 8285
rect 13265 8245 13277 8279
rect 13311 8276 13323 8279
rect 13538 8276 13544 8288
rect 13311 8248 13544 8276
rect 13311 8245 13323 8248
rect 13265 8239 13323 8245
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 19242 8236 19248 8288
rect 19300 8276 19306 8288
rect 19337 8279 19395 8285
rect 19337 8276 19349 8279
rect 19300 8248 19349 8276
rect 19300 8236 19306 8248
rect 19337 8245 19349 8248
rect 19383 8245 19395 8279
rect 19337 8239 19395 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 13725 8075 13783 8081
rect 13725 8041 13737 8075
rect 13771 8072 13783 8075
rect 14182 8072 14188 8084
rect 13771 8044 14188 8072
rect 13771 8041 13783 8044
rect 13725 8035 13783 8041
rect 14182 8032 14188 8044
rect 14240 8072 14246 8084
rect 15289 8075 15347 8081
rect 15289 8072 15301 8075
rect 14240 8044 15301 8072
rect 14240 8032 14246 8044
rect 15289 8041 15301 8044
rect 15335 8041 15347 8075
rect 15654 8072 15660 8084
rect 15567 8044 15660 8072
rect 15289 8035 15347 8041
rect 15654 8032 15660 8044
rect 15712 8072 15718 8084
rect 16390 8072 16396 8084
rect 15712 8044 16396 8072
rect 15712 8032 15718 8044
rect 16390 8032 16396 8044
rect 16448 8032 16454 8084
rect 16666 8072 16672 8084
rect 16627 8044 16672 8072
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 18322 8072 18328 8084
rect 18283 8044 18328 8072
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 18969 8075 19027 8081
rect 18969 8041 18981 8075
rect 19015 8072 19027 8075
rect 19242 8072 19248 8084
rect 19015 8044 19248 8072
rect 19015 8041 19027 8044
rect 18969 8035 19027 8041
rect 19242 8032 19248 8044
rect 19300 8072 19306 8084
rect 20901 8075 20959 8081
rect 20901 8072 20913 8075
rect 19300 8044 20913 8072
rect 19300 8032 19306 8044
rect 20901 8041 20913 8044
rect 20947 8041 20959 8075
rect 21266 8072 21272 8084
rect 21227 8044 21272 8072
rect 20901 8035 20959 8041
rect 21266 8032 21272 8044
rect 21324 8032 21330 8084
rect 25038 8032 25044 8084
rect 25096 8072 25102 8084
rect 25225 8075 25283 8081
rect 25225 8072 25237 8075
rect 25096 8044 25237 8072
rect 25096 8032 25102 8044
rect 25225 8041 25237 8044
rect 25271 8041 25283 8075
rect 25225 8035 25283 8041
rect 1486 7964 1492 8016
rect 1544 8004 1550 8016
rect 9582 8004 9588 8016
rect 1544 7976 9588 8004
rect 1544 7964 1550 7976
rect 9582 7964 9588 7976
rect 9640 7964 9646 8016
rect 11882 7964 11888 8016
rect 11940 8004 11946 8016
rect 13630 8004 13636 8016
rect 11940 7976 13636 8004
rect 11940 7964 11946 7976
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 15749 8007 15807 8013
rect 15749 7973 15761 8007
rect 15795 8004 15807 8007
rect 15930 8004 15936 8016
rect 15795 7976 15936 8004
rect 15795 7973 15807 7976
rect 15749 7967 15807 7973
rect 15930 7964 15936 7976
rect 15988 7964 15994 8016
rect 23201 8007 23259 8013
rect 23201 7973 23213 8007
rect 23247 8004 23259 8007
rect 24026 8004 24032 8016
rect 23247 7976 24032 8004
rect 23247 7973 23259 7976
rect 23201 7967 23259 7973
rect 24026 7964 24032 7976
rect 24084 7964 24090 8016
rect 17218 7945 17224 7948
rect 17212 7899 17224 7945
rect 17276 7936 17282 7948
rect 22833 7939 22891 7945
rect 17276 7908 17312 7936
rect 17218 7896 17224 7899
rect 17276 7896 17282 7908
rect 22833 7905 22845 7939
rect 22879 7936 22891 7939
rect 23290 7936 23296 7948
rect 22879 7908 23296 7936
rect 22879 7905 22891 7908
rect 22833 7899 22891 7905
rect 13814 7868 13820 7880
rect 13775 7840 13820 7868
rect 13814 7828 13820 7840
rect 13872 7828 13878 7880
rect 13909 7871 13967 7877
rect 13909 7837 13921 7871
rect 13955 7837 13967 7871
rect 13909 7831 13967 7837
rect 15933 7871 15991 7877
rect 15933 7837 15945 7871
rect 15979 7868 15991 7871
rect 16390 7868 16396 7880
rect 15979 7840 16396 7868
rect 15979 7837 15991 7840
rect 15933 7831 15991 7837
rect 13170 7760 13176 7812
rect 13228 7800 13234 7812
rect 13924 7800 13952 7831
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 16945 7871 17003 7877
rect 16945 7868 16957 7871
rect 16632 7840 16957 7868
rect 16632 7828 16638 7840
rect 16945 7837 16957 7840
rect 16991 7837 17003 7871
rect 19426 7868 19432 7880
rect 19387 7840 19432 7868
rect 16945 7831 17003 7837
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 20070 7828 20076 7880
rect 20128 7868 20134 7880
rect 21361 7871 21419 7877
rect 21361 7868 21373 7871
rect 20128 7840 21373 7868
rect 20128 7828 20134 7840
rect 21361 7837 21373 7840
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7868 21603 7871
rect 21634 7868 21640 7880
rect 21591 7840 21640 7868
rect 21591 7837 21603 7840
rect 21545 7831 21603 7837
rect 21634 7828 21640 7840
rect 21692 7828 21698 7880
rect 19334 7800 19340 7812
rect 13228 7772 13952 7800
rect 19295 7772 19340 7800
rect 13228 7760 13234 7772
rect 19334 7760 19340 7772
rect 19392 7760 19398 7812
rect 13354 7732 13360 7744
rect 13315 7704 13360 7732
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 14369 7735 14427 7741
rect 14369 7732 14381 7735
rect 13596 7704 14381 7732
rect 13596 7692 13602 7704
rect 14369 7701 14381 7704
rect 14415 7701 14427 7735
rect 14369 7695 14427 7701
rect 16393 7735 16451 7741
rect 16393 7701 16405 7735
rect 16439 7732 16451 7735
rect 16482 7732 16488 7744
rect 16439 7704 16488 7732
rect 16439 7701 16451 7704
rect 16393 7695 16451 7701
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 20717 7735 20775 7741
rect 20717 7701 20729 7735
rect 20763 7732 20775 7735
rect 21450 7732 21456 7744
rect 20763 7704 21456 7732
rect 20763 7701 20775 7704
rect 20717 7695 20775 7701
rect 21450 7692 21456 7704
rect 21508 7692 21514 7744
rect 21542 7692 21548 7744
rect 21600 7732 21606 7744
rect 21910 7732 21916 7744
rect 21600 7704 21916 7732
rect 21600 7692 21606 7704
rect 21910 7692 21916 7704
rect 21968 7732 21974 7744
rect 22005 7735 22063 7741
rect 22005 7732 22017 7735
rect 21968 7704 22017 7732
rect 21968 7692 21974 7704
rect 22005 7701 22017 7704
rect 22051 7732 22063 7735
rect 22848 7732 22876 7899
rect 23290 7896 23296 7908
rect 23348 7896 23354 7948
rect 23382 7896 23388 7948
rect 23440 7936 23446 7948
rect 23566 7945 23572 7948
rect 23560 7936 23572 7945
rect 23440 7908 23572 7936
rect 23440 7896 23446 7908
rect 23560 7899 23572 7908
rect 23624 7936 23630 7948
rect 24854 7936 24860 7948
rect 23624 7908 24860 7936
rect 23566 7896 23572 7899
rect 23624 7896 23630 7908
rect 24854 7896 24860 7908
rect 24912 7896 24918 7948
rect 22051 7704 22876 7732
rect 22051 7701 22063 7704
rect 22005 7695 22063 7701
rect 24210 7692 24216 7744
rect 24268 7732 24274 7744
rect 24673 7735 24731 7741
rect 24673 7732 24685 7735
rect 24268 7704 24685 7732
rect 24268 7692 24274 7704
rect 24673 7701 24685 7704
rect 24719 7701 24731 7735
rect 24673 7695 24731 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 13081 7531 13139 7537
rect 13081 7497 13093 7531
rect 13127 7528 13139 7531
rect 13170 7528 13176 7540
rect 13127 7500 13176 7528
rect 13127 7497 13139 7500
rect 13081 7491 13139 7497
rect 13170 7488 13176 7500
rect 13228 7488 13234 7540
rect 15565 7531 15623 7537
rect 15565 7497 15577 7531
rect 15611 7528 15623 7531
rect 15654 7528 15660 7540
rect 15611 7500 15660 7528
rect 15611 7497 15623 7500
rect 15565 7491 15623 7497
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 15930 7528 15936 7540
rect 15891 7500 15936 7528
rect 15930 7488 15936 7500
rect 15988 7488 15994 7540
rect 17129 7531 17187 7537
rect 17129 7497 17141 7531
rect 17175 7528 17187 7531
rect 17218 7528 17224 7540
rect 17175 7500 17224 7528
rect 17175 7497 17187 7500
rect 17129 7491 17187 7497
rect 17218 7488 17224 7500
rect 17276 7488 17282 7540
rect 19334 7488 19340 7540
rect 19392 7528 19398 7540
rect 20070 7528 20076 7540
rect 19392 7500 20076 7528
rect 19392 7488 19398 7500
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 21266 7488 21272 7540
rect 21324 7528 21330 7540
rect 22005 7531 22063 7537
rect 22005 7528 22017 7531
rect 21324 7500 22017 7528
rect 21324 7488 21330 7500
rect 22005 7497 22017 7500
rect 22051 7497 22063 7531
rect 25406 7528 25412 7540
rect 25367 7500 25412 7528
rect 22005 7491 22063 7497
rect 25406 7488 25412 7500
rect 25464 7488 25470 7540
rect 15102 7420 15108 7472
rect 15160 7460 15166 7472
rect 16025 7463 16083 7469
rect 16025 7460 16037 7463
rect 15160 7432 16037 7460
rect 15160 7420 15166 7432
rect 16025 7429 16037 7432
rect 16071 7429 16083 7463
rect 16025 7423 16083 7429
rect 19521 7463 19579 7469
rect 19521 7429 19533 7463
rect 19567 7460 19579 7463
rect 19978 7460 19984 7472
rect 19567 7432 19984 7460
rect 19567 7429 19579 7432
rect 19521 7423 19579 7429
rect 19978 7420 19984 7432
rect 20036 7420 20042 7472
rect 21634 7460 21640 7472
rect 21595 7432 21640 7460
rect 21634 7420 21640 7432
rect 21692 7420 21698 7472
rect 13449 7395 13507 7401
rect 13449 7361 13461 7395
rect 13495 7392 13507 7395
rect 16482 7392 16488 7404
rect 13495 7364 13676 7392
rect 16443 7364 16488 7392
rect 13495 7361 13507 7364
rect 13449 7355 13507 7361
rect 12618 7284 12624 7336
rect 12676 7324 12682 7336
rect 13538 7324 13544 7336
rect 12676 7296 13544 7324
rect 12676 7284 12682 7296
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 13648 7324 13676 7364
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 16577 7395 16635 7401
rect 16577 7361 16589 7395
rect 16623 7361 16635 7395
rect 16577 7355 16635 7361
rect 13808 7327 13866 7333
rect 13808 7324 13820 7327
rect 13648 7296 13820 7324
rect 13808 7293 13820 7296
rect 13854 7324 13866 7327
rect 14734 7324 14740 7336
rect 13854 7296 14740 7324
rect 13854 7293 13866 7296
rect 13808 7287 13866 7293
rect 14734 7284 14740 7296
rect 14792 7284 14798 7336
rect 16390 7284 16396 7336
rect 16448 7324 16454 7336
rect 16592 7324 16620 7355
rect 16666 7352 16672 7404
rect 16724 7392 16730 7404
rect 17862 7392 17868 7404
rect 16724 7364 17868 7392
rect 16724 7352 16730 7364
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 20898 7352 20904 7404
rect 20956 7392 20962 7404
rect 21085 7395 21143 7401
rect 21085 7392 21097 7395
rect 20956 7364 21097 7392
rect 20956 7352 20962 7364
rect 21085 7361 21097 7364
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 21269 7395 21327 7401
rect 21269 7361 21281 7395
rect 21315 7392 21327 7395
rect 21450 7392 21456 7404
rect 21315 7364 21456 7392
rect 21315 7361 21327 7364
rect 21269 7355 21327 7361
rect 21450 7352 21456 7364
rect 21508 7352 21514 7404
rect 24210 7352 24216 7404
rect 24268 7392 24274 7404
rect 24305 7395 24363 7401
rect 24305 7392 24317 7395
rect 24268 7364 24317 7392
rect 24268 7352 24274 7364
rect 24305 7361 24317 7364
rect 24351 7392 24363 7395
rect 24489 7395 24547 7401
rect 24489 7392 24501 7395
rect 24351 7364 24501 7392
rect 24351 7361 24363 7364
rect 24305 7355 24363 7361
rect 24489 7361 24501 7364
rect 24535 7361 24547 7395
rect 24489 7355 24547 7361
rect 16448 7296 16620 7324
rect 18141 7327 18199 7333
rect 16448 7284 16454 7296
rect 18141 7293 18153 7327
rect 18187 7324 18199 7327
rect 18230 7324 18236 7336
rect 18187 7296 18236 7324
rect 18187 7293 18199 7296
rect 18141 7287 18199 7293
rect 18230 7284 18236 7296
rect 18288 7284 18294 7336
rect 22186 7324 22192 7336
rect 22147 7296 22192 7324
rect 22186 7284 22192 7296
rect 22244 7324 22250 7336
rect 22741 7327 22799 7333
rect 22741 7324 22753 7327
rect 22244 7296 22753 7324
rect 22244 7284 22250 7296
rect 22741 7293 22753 7296
rect 22787 7293 22799 7327
rect 24026 7324 24032 7336
rect 23987 7296 24032 7324
rect 22741 7287 22799 7293
rect 24026 7284 24032 7296
rect 24084 7284 24090 7336
rect 25222 7324 25228 7336
rect 25183 7296 25228 7324
rect 25222 7284 25228 7296
rect 25280 7324 25286 7336
rect 25777 7327 25835 7333
rect 25777 7324 25789 7327
rect 25280 7296 25789 7324
rect 25280 7284 25286 7296
rect 25777 7293 25789 7296
rect 25823 7293 25835 7327
rect 25777 7287 25835 7293
rect 15562 7216 15568 7268
rect 15620 7256 15626 7268
rect 16206 7256 16212 7268
rect 15620 7228 16212 7256
rect 15620 7216 15626 7228
rect 16206 7216 16212 7228
rect 16264 7256 16270 7268
rect 17862 7256 17868 7268
rect 16264 7228 16436 7256
rect 17775 7228 17868 7256
rect 16264 7216 16270 7228
rect 12526 7188 12532 7200
rect 12487 7160 12532 7188
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 14918 7188 14924 7200
rect 14879 7160 14924 7188
rect 14918 7148 14924 7160
rect 14976 7148 14982 7200
rect 16408 7197 16436 7228
rect 17862 7216 17868 7228
rect 17920 7256 17926 7268
rect 18408 7259 18466 7265
rect 18408 7256 18420 7259
rect 17920 7228 18420 7256
rect 17920 7216 17926 7228
rect 18408 7225 18420 7228
rect 18454 7256 18466 7259
rect 19242 7256 19248 7268
rect 18454 7228 19248 7256
rect 18454 7225 18466 7228
rect 18408 7219 18466 7225
rect 19242 7216 19248 7228
rect 19300 7216 19306 7268
rect 20993 7259 21051 7265
rect 20993 7256 21005 7259
rect 20456 7228 21005 7256
rect 16393 7191 16451 7197
rect 16393 7157 16405 7191
rect 16439 7157 16451 7191
rect 16393 7151 16451 7157
rect 16574 7148 16580 7200
rect 16632 7188 16638 7200
rect 17405 7191 17463 7197
rect 17405 7188 17417 7191
rect 16632 7160 17417 7188
rect 16632 7148 16638 7160
rect 17405 7157 17417 7160
rect 17451 7157 17463 7191
rect 17405 7151 17463 7157
rect 19334 7148 19340 7200
rect 19392 7188 19398 7200
rect 20456 7197 20484 7228
rect 20993 7225 21005 7228
rect 21039 7225 21051 7259
rect 20993 7219 21051 7225
rect 23382 7216 23388 7268
rect 23440 7256 23446 7268
rect 24121 7259 24179 7265
rect 24121 7256 24133 7259
rect 23440 7228 24133 7256
rect 23440 7216 23446 7228
rect 24121 7225 24133 7228
rect 24167 7256 24179 7259
rect 25041 7259 25099 7265
rect 25041 7256 25053 7259
rect 24167 7228 25053 7256
rect 24167 7225 24179 7228
rect 24121 7219 24179 7225
rect 25041 7225 25053 7228
rect 25087 7225 25099 7259
rect 25041 7219 25099 7225
rect 20441 7191 20499 7197
rect 20441 7188 20453 7191
rect 19392 7160 20453 7188
rect 19392 7148 19398 7160
rect 20441 7157 20453 7160
rect 20487 7157 20499 7191
rect 20622 7188 20628 7200
rect 20583 7160 20628 7188
rect 20441 7151 20499 7157
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 22370 7188 22376 7200
rect 22331 7160 22376 7188
rect 22370 7148 22376 7160
rect 22428 7148 22434 7200
rect 23014 7148 23020 7200
rect 23072 7188 23078 7200
rect 23293 7191 23351 7197
rect 23293 7188 23305 7191
rect 23072 7160 23305 7188
rect 23072 7148 23078 7160
rect 23293 7157 23305 7160
rect 23339 7188 23351 7191
rect 23566 7188 23572 7200
rect 23339 7160 23572 7188
rect 23339 7157 23351 7160
rect 23293 7151 23351 7157
rect 23566 7148 23572 7160
rect 23624 7148 23630 7200
rect 23661 7191 23719 7197
rect 23661 7157 23673 7191
rect 23707 7188 23719 7191
rect 24026 7188 24032 7200
rect 23707 7160 24032 7188
rect 23707 7157 23719 7160
rect 23661 7151 23719 7157
rect 24026 7148 24032 7160
rect 24084 7148 24090 7200
rect 24489 7191 24547 7197
rect 24489 7157 24501 7191
rect 24535 7188 24547 7191
rect 24765 7191 24823 7197
rect 24765 7188 24777 7191
rect 24535 7160 24777 7188
rect 24535 7157 24547 7160
rect 24489 7151 24547 7157
rect 24765 7157 24777 7160
rect 24811 7188 24823 7191
rect 25406 7188 25412 7200
rect 24811 7160 25412 7188
rect 24811 7157 24823 7160
rect 24765 7151 24823 7157
rect 25406 7148 25412 7160
rect 25464 7148 25470 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 13170 6984 13176 6996
rect 13131 6956 13176 6984
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 16206 6984 16212 6996
rect 16167 6956 16212 6984
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 17770 6944 17776 6996
rect 17828 6984 17834 6996
rect 18414 6984 18420 6996
rect 17828 6956 18420 6984
rect 17828 6944 17834 6956
rect 18414 6944 18420 6956
rect 18472 6984 18478 6996
rect 18601 6987 18659 6993
rect 18601 6984 18613 6987
rect 18472 6956 18613 6984
rect 18472 6944 18478 6956
rect 18601 6953 18613 6956
rect 18647 6953 18659 6987
rect 18601 6947 18659 6953
rect 20717 6987 20775 6993
rect 20717 6953 20729 6987
rect 20763 6984 20775 6987
rect 20898 6984 20904 6996
rect 20763 6956 20904 6984
rect 20763 6953 20775 6956
rect 20717 6947 20775 6953
rect 20898 6944 20904 6956
rect 20956 6944 20962 6996
rect 23290 6944 23296 6996
rect 23348 6984 23354 6996
rect 23661 6987 23719 6993
rect 23661 6984 23673 6987
rect 23348 6956 23673 6984
rect 23348 6944 23354 6956
rect 23661 6953 23673 6956
rect 23707 6953 23719 6987
rect 25130 6984 25136 6996
rect 25091 6956 25136 6984
rect 23661 6947 23719 6953
rect 25130 6944 25136 6956
rect 25188 6944 25194 6996
rect 14918 6876 14924 6928
rect 14976 6916 14982 6928
rect 15473 6919 15531 6925
rect 15473 6916 15485 6919
rect 14976 6888 15485 6916
rect 14976 6876 14982 6888
rect 15473 6885 15485 6888
rect 15519 6916 15531 6919
rect 16390 6916 16396 6928
rect 15519 6888 16396 6916
rect 15519 6885 15531 6888
rect 15473 6879 15531 6885
rect 16390 6876 16396 6888
rect 16448 6916 16454 6928
rect 16485 6919 16543 6925
rect 16485 6916 16497 6919
rect 16448 6888 16497 6916
rect 16448 6876 16454 6888
rect 16485 6885 16497 6888
rect 16531 6885 16543 6919
rect 21266 6916 21272 6928
rect 16485 6879 16543 6885
rect 20640 6888 21272 6916
rect 12066 6857 12072 6860
rect 12060 6848 12072 6857
rect 12027 6820 12072 6848
rect 12060 6811 12072 6820
rect 12066 6808 12072 6811
rect 12124 6808 12130 6860
rect 14182 6848 14188 6860
rect 14143 6820 14188 6848
rect 14182 6808 14188 6820
rect 14240 6808 14246 6860
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 15105 6851 15163 6857
rect 15105 6848 15117 6851
rect 14884 6820 15117 6848
rect 14884 6808 14890 6820
rect 15105 6817 15117 6820
rect 15151 6817 15163 6851
rect 15105 6811 15163 6817
rect 17037 6851 17095 6857
rect 17037 6817 17049 6851
rect 17083 6848 17095 6851
rect 17681 6851 17739 6857
rect 17681 6848 17693 6851
rect 17083 6820 17693 6848
rect 17083 6817 17095 6820
rect 17037 6811 17095 6817
rect 17681 6817 17693 6820
rect 17727 6817 17739 6851
rect 17681 6811 17739 6817
rect 11790 6780 11796 6792
rect 11751 6752 11796 6780
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 15654 6780 15660 6792
rect 15615 6752 15660 6780
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 17126 6780 17132 6792
rect 17087 6752 17132 6780
rect 17126 6740 17132 6752
rect 17184 6740 17190 6792
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17276 6752 17321 6780
rect 17276 6740 17282 6752
rect 13814 6712 13820 6724
rect 13727 6684 13820 6712
rect 13814 6672 13820 6684
rect 13872 6712 13878 6724
rect 15102 6712 15108 6724
rect 13872 6684 15108 6712
rect 13872 6672 13878 6684
rect 15102 6672 15108 6684
rect 15160 6672 15166 6724
rect 17696 6712 17724 6811
rect 18690 6808 18696 6860
rect 18748 6848 18754 6860
rect 19150 6848 19156 6860
rect 18748 6820 19156 6848
rect 18748 6808 18754 6820
rect 19150 6808 19156 6820
rect 19208 6808 19214 6860
rect 20349 6851 20407 6857
rect 20349 6817 20361 6851
rect 20395 6848 20407 6851
rect 20640 6848 20668 6888
rect 21266 6876 21272 6888
rect 21324 6876 21330 6928
rect 23569 6919 23627 6925
rect 23569 6916 23581 6919
rect 23400 6888 23581 6916
rect 20395 6820 20668 6848
rect 20395 6817 20407 6820
rect 20349 6811 20407 6817
rect 22646 6808 22652 6860
rect 22704 6848 22710 6860
rect 23400 6848 23428 6888
rect 23569 6885 23581 6888
rect 23615 6916 23627 6919
rect 23615 6888 25360 6916
rect 23615 6885 23627 6888
rect 23569 6879 23627 6885
rect 25332 6860 25360 6888
rect 22704 6820 23428 6848
rect 22704 6808 22710 6820
rect 25314 6808 25320 6860
rect 25372 6808 25378 6860
rect 18785 6783 18843 6789
rect 18785 6780 18797 6783
rect 18708 6752 18797 6780
rect 18233 6715 18291 6721
rect 18233 6712 18245 6715
rect 17696 6684 18245 6712
rect 18233 6681 18245 6684
rect 18279 6681 18291 6715
rect 18233 6675 18291 6681
rect 18708 6656 18736 6752
rect 18785 6749 18797 6752
rect 18831 6749 18843 6783
rect 18785 6743 18843 6749
rect 19797 6783 19855 6789
rect 19797 6749 19809 6783
rect 19843 6780 19855 6783
rect 20162 6780 20168 6792
rect 19843 6752 20168 6780
rect 19843 6749 19855 6752
rect 19797 6743 19855 6749
rect 20162 6740 20168 6752
rect 20220 6740 20226 6792
rect 20438 6740 20444 6792
rect 20496 6780 20502 6792
rect 21361 6783 21419 6789
rect 21361 6780 21373 6783
rect 20496 6752 21373 6780
rect 20496 6740 20502 6752
rect 21361 6749 21373 6752
rect 21407 6749 21419 6783
rect 21542 6780 21548 6792
rect 21503 6752 21548 6780
rect 21361 6743 21419 6749
rect 21542 6740 21548 6752
rect 21600 6740 21606 6792
rect 23014 6740 23020 6792
rect 23072 6780 23078 6792
rect 23753 6783 23811 6789
rect 23072 6752 23612 6780
rect 23072 6740 23078 6752
rect 22002 6672 22008 6724
rect 22060 6712 22066 6724
rect 23201 6715 23259 6721
rect 22060 6684 22968 6712
rect 22060 6672 22066 6684
rect 22940 6656 22968 6684
rect 23201 6681 23213 6715
rect 23247 6712 23259 6715
rect 23382 6712 23388 6724
rect 23247 6684 23388 6712
rect 23247 6681 23259 6684
rect 23201 6675 23259 6681
rect 23382 6672 23388 6684
rect 23440 6672 23446 6724
rect 23584 6712 23612 6752
rect 23753 6749 23765 6783
rect 23799 6749 23811 6783
rect 23753 6743 23811 6749
rect 23768 6712 23796 6743
rect 24946 6740 24952 6792
rect 25004 6780 25010 6792
rect 25225 6783 25283 6789
rect 25225 6780 25237 6783
rect 25004 6752 25237 6780
rect 25004 6740 25010 6752
rect 25225 6749 25237 6752
rect 25271 6749 25283 6783
rect 25406 6780 25412 6792
rect 25367 6752 25412 6780
rect 25225 6743 25283 6749
rect 25406 6740 25412 6752
rect 25464 6740 25470 6792
rect 24210 6712 24216 6724
rect 23584 6684 23796 6712
rect 24171 6684 24216 6712
rect 24210 6672 24216 6684
rect 24268 6672 24274 6724
rect 14734 6604 14740 6656
rect 14792 6644 14798 6656
rect 14921 6647 14979 6653
rect 14921 6644 14933 6647
rect 14792 6616 14933 6644
rect 14792 6604 14798 6616
rect 14921 6613 14933 6616
rect 14967 6644 14979 6647
rect 16482 6644 16488 6656
rect 14967 6616 16488 6644
rect 14967 6613 14979 6616
rect 14921 6607 14979 6613
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 16669 6647 16727 6653
rect 16669 6613 16681 6647
rect 16715 6644 16727 6647
rect 16850 6644 16856 6656
rect 16715 6616 16856 6644
rect 16715 6613 16727 6616
rect 16669 6607 16727 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 18141 6647 18199 6653
rect 18141 6613 18153 6647
rect 18187 6644 18199 6647
rect 18690 6644 18696 6656
rect 18187 6616 18696 6644
rect 18187 6613 18199 6616
rect 18141 6607 18199 6613
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 19337 6647 19395 6653
rect 19337 6613 19349 6647
rect 19383 6644 19395 6647
rect 19518 6644 19524 6656
rect 19383 6616 19524 6644
rect 19383 6613 19395 6616
rect 19337 6607 19395 6613
rect 19518 6604 19524 6616
rect 19576 6604 19582 6656
rect 19610 6604 19616 6656
rect 19668 6644 19674 6656
rect 20898 6644 20904 6656
rect 19668 6616 19713 6644
rect 20859 6616 20904 6644
rect 19668 6604 19674 6616
rect 20898 6604 20904 6616
rect 20956 6604 20962 6656
rect 22922 6604 22928 6656
rect 22980 6644 22986 6656
rect 23017 6647 23075 6653
rect 23017 6644 23029 6647
rect 22980 6616 23029 6644
rect 22980 6604 22986 6616
rect 23017 6613 23029 6616
rect 23063 6644 23075 6647
rect 23290 6644 23296 6656
rect 23063 6616 23296 6644
rect 23063 6613 23075 6616
rect 23017 6607 23075 6613
rect 23290 6604 23296 6616
rect 23348 6604 23354 6656
rect 24118 6604 24124 6656
rect 24176 6644 24182 6656
rect 24765 6647 24823 6653
rect 24765 6644 24777 6647
rect 24176 6616 24777 6644
rect 24176 6604 24182 6616
rect 24765 6613 24777 6616
rect 24811 6613 24823 6647
rect 24765 6607 24823 6613
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 11885 6443 11943 6449
rect 11885 6409 11897 6443
rect 11931 6440 11943 6443
rect 12066 6440 12072 6452
rect 11931 6412 12072 6440
rect 11931 6409 11943 6412
rect 11885 6403 11943 6409
rect 12066 6400 12072 6412
rect 12124 6400 12130 6452
rect 17497 6443 17555 6449
rect 17497 6409 17509 6443
rect 17543 6440 17555 6443
rect 17770 6440 17776 6452
rect 17543 6412 17776 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 21542 6400 21548 6452
rect 21600 6440 21606 6452
rect 21913 6443 21971 6449
rect 21913 6440 21925 6443
rect 21600 6412 21925 6440
rect 21600 6400 21606 6412
rect 21913 6409 21925 6412
rect 21959 6409 21971 6443
rect 22646 6440 22652 6452
rect 22607 6412 22652 6440
rect 21913 6403 21971 6409
rect 22646 6400 22652 6412
rect 22704 6400 22710 6452
rect 23106 6440 23112 6452
rect 23067 6412 23112 6440
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 23658 6440 23664 6452
rect 23619 6412 23664 6440
rect 23658 6400 23664 6412
rect 23716 6400 23722 6452
rect 24857 6443 24915 6449
rect 24857 6409 24869 6443
rect 24903 6440 24915 6443
rect 24946 6440 24952 6452
rect 24903 6412 24952 6440
rect 24903 6409 24915 6412
rect 24857 6403 24915 6409
rect 24946 6400 24952 6412
rect 25004 6400 25010 6452
rect 16301 6375 16359 6381
rect 16301 6341 16313 6375
rect 16347 6372 16359 6375
rect 19150 6372 19156 6384
rect 16347 6344 17080 6372
rect 19111 6344 19156 6372
rect 16347 6341 16359 6344
rect 16301 6335 16359 6341
rect 17052 6313 17080 6344
rect 19150 6332 19156 6344
rect 19208 6332 19214 6384
rect 23477 6375 23535 6381
rect 23477 6341 23489 6375
rect 23523 6372 23535 6375
rect 23566 6372 23572 6384
rect 23523 6344 23572 6372
rect 23523 6341 23535 6344
rect 23477 6335 23535 6341
rect 23566 6332 23572 6344
rect 23624 6332 23630 6384
rect 14829 6307 14887 6313
rect 14829 6273 14841 6307
rect 14875 6304 14887 6307
rect 17037 6307 17095 6313
rect 14875 6276 16804 6304
rect 14875 6273 14887 6276
rect 14829 6267 14887 6273
rect 16776 6248 16804 6276
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17862 6304 17868 6316
rect 17083 6276 17868 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17862 6264 17868 6276
rect 17920 6264 17926 6316
rect 18690 6304 18696 6316
rect 18651 6276 18696 6304
rect 18690 6264 18696 6276
rect 18748 6304 18754 6316
rect 19429 6307 19487 6313
rect 19429 6304 19441 6307
rect 18748 6276 19441 6304
rect 18748 6264 18754 6276
rect 19429 6273 19441 6276
rect 19475 6273 19487 6307
rect 24210 6304 24216 6316
rect 24171 6276 24216 6304
rect 19429 6267 19487 6273
rect 24210 6264 24216 6276
rect 24268 6264 24274 6316
rect 11517 6239 11575 6245
rect 11517 6205 11529 6239
rect 11563 6236 11575 6239
rect 11790 6236 11796 6248
rect 11563 6208 11796 6236
rect 11563 6205 11575 6208
rect 11517 6199 11575 6205
rect 11790 6196 11796 6208
rect 11848 6236 11854 6248
rect 12618 6236 12624 6248
rect 11848 6208 12624 6236
rect 11848 6196 11854 6208
rect 12618 6196 12624 6208
rect 12676 6236 12682 6248
rect 12713 6239 12771 6245
rect 12713 6236 12725 6239
rect 12676 6208 12725 6236
rect 12676 6196 12682 6208
rect 12713 6205 12725 6208
rect 12759 6205 12771 6239
rect 12713 6199 12771 6205
rect 15289 6239 15347 6245
rect 15289 6205 15301 6239
rect 15335 6236 15347 6239
rect 16758 6236 16764 6248
rect 15335 6208 15369 6236
rect 16671 6208 16764 6236
rect 15335 6205 15347 6208
rect 15289 6199 15347 6205
rect 12253 6171 12311 6177
rect 12253 6137 12265 6171
rect 12299 6168 12311 6171
rect 12980 6171 13038 6177
rect 12980 6168 12992 6171
rect 12299 6140 12992 6168
rect 12299 6137 12311 6140
rect 12253 6131 12311 6137
rect 12980 6137 12992 6140
rect 13026 6168 13038 6171
rect 13170 6168 13176 6180
rect 13026 6140 13176 6168
rect 13026 6137 13038 6140
rect 12980 6131 13038 6137
rect 13170 6128 13176 6140
rect 13228 6128 13234 6180
rect 15197 6171 15255 6177
rect 15197 6137 15209 6171
rect 15243 6168 15255 6171
rect 15304 6168 15332 6199
rect 16758 6196 16764 6208
rect 16816 6196 16822 6248
rect 18506 6236 18512 6248
rect 18467 6208 18512 6236
rect 18506 6196 18512 6208
rect 18564 6196 18570 6248
rect 19610 6196 19616 6248
rect 19668 6236 19674 6248
rect 19797 6239 19855 6245
rect 19797 6236 19809 6239
rect 19668 6208 19809 6236
rect 19668 6196 19674 6208
rect 19797 6205 19809 6208
rect 19843 6205 19855 6239
rect 20530 6236 20536 6248
rect 20491 6208 20536 6236
rect 19797 6199 19855 6205
rect 20530 6196 20536 6208
rect 20588 6196 20594 6248
rect 23106 6196 23112 6248
rect 23164 6236 23170 6248
rect 24121 6239 24179 6245
rect 24121 6236 24133 6239
rect 23164 6208 24133 6236
rect 23164 6196 23170 6208
rect 24121 6205 24133 6208
rect 24167 6205 24179 6239
rect 24121 6199 24179 6205
rect 24854 6196 24860 6248
rect 24912 6236 24918 6248
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 24912 6208 25237 6236
rect 24912 6196 24918 6208
rect 25225 6205 25237 6208
rect 25271 6236 25283 6239
rect 25961 6239 26019 6245
rect 25961 6236 25973 6239
rect 25271 6208 25973 6236
rect 25271 6205 25283 6208
rect 25225 6199 25283 6205
rect 25961 6205 25973 6208
rect 26007 6205 26019 6239
rect 25961 6199 26019 6205
rect 16298 6168 16304 6180
rect 15243 6140 16304 6168
rect 15243 6137 15255 6140
rect 15197 6131 15255 6137
rect 16298 6128 16304 6140
rect 16356 6128 16362 6180
rect 18417 6171 18475 6177
rect 18417 6168 18429 6171
rect 17788 6140 18429 6168
rect 14093 6103 14151 6109
rect 14093 6069 14105 6103
rect 14139 6100 14151 6103
rect 14182 6100 14188 6112
rect 14139 6072 14188 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 15470 6100 15476 6112
rect 15431 6072 15476 6100
rect 15470 6060 15476 6072
rect 15528 6060 15534 6112
rect 15930 6100 15936 6112
rect 15891 6072 15936 6100
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16390 6100 16396 6112
rect 16351 6072 16396 6100
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 16908 6072 16953 6100
rect 16908 6060 16914 6072
rect 17494 6060 17500 6112
rect 17552 6100 17558 6112
rect 17788 6109 17816 6140
rect 18417 6137 18429 6140
rect 18463 6168 18475 6171
rect 19334 6168 19340 6180
rect 18463 6140 19340 6168
rect 18463 6137 18475 6140
rect 18417 6131 18475 6137
rect 19334 6128 19340 6140
rect 19392 6128 19398 6180
rect 20441 6171 20499 6177
rect 20441 6137 20453 6171
rect 20487 6168 20499 6171
rect 20800 6171 20858 6177
rect 20800 6168 20812 6171
rect 20487 6140 20812 6168
rect 20487 6137 20499 6140
rect 20441 6131 20499 6137
rect 20800 6137 20812 6140
rect 20846 6168 20858 6171
rect 21450 6168 21456 6180
rect 20846 6140 21456 6168
rect 20846 6137 20858 6140
rect 20800 6131 20858 6137
rect 21450 6128 21456 6140
rect 21508 6128 21514 6180
rect 23566 6128 23572 6180
rect 23624 6168 23630 6180
rect 24029 6171 24087 6177
rect 24029 6168 24041 6171
rect 23624 6140 24041 6168
rect 23624 6128 23630 6140
rect 24029 6137 24041 6140
rect 24075 6137 24087 6171
rect 25498 6168 25504 6180
rect 25459 6140 25504 6168
rect 24029 6131 24087 6137
rect 25498 6128 25504 6140
rect 25556 6128 25562 6180
rect 17773 6103 17831 6109
rect 17773 6100 17785 6103
rect 17552 6072 17785 6100
rect 17552 6060 17558 6072
rect 17773 6069 17785 6072
rect 17819 6069 17831 6103
rect 17773 6063 17831 6069
rect 17862 6060 17868 6112
rect 17920 6100 17926 6112
rect 18049 6103 18107 6109
rect 18049 6100 18061 6103
rect 17920 6072 18061 6100
rect 17920 6060 17926 6072
rect 18049 6069 18061 6072
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 19518 6060 19524 6112
rect 19576 6100 19582 6112
rect 19613 6103 19671 6109
rect 19613 6100 19625 6103
rect 19576 6072 19625 6100
rect 19576 6060 19582 6072
rect 19613 6069 19625 6072
rect 19659 6069 19671 6103
rect 19613 6063 19671 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 12897 5899 12955 5905
rect 12897 5865 12909 5899
rect 12943 5896 12955 5899
rect 13354 5896 13360 5908
rect 12943 5868 13360 5896
rect 12943 5865 12955 5868
rect 12897 5859 12955 5865
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 14826 5856 14832 5908
rect 14884 5896 14890 5908
rect 14921 5899 14979 5905
rect 14921 5896 14933 5899
rect 14884 5868 14933 5896
rect 14884 5856 14890 5868
rect 14921 5865 14933 5868
rect 14967 5865 14979 5899
rect 14921 5859 14979 5865
rect 15657 5899 15715 5905
rect 15657 5865 15669 5899
rect 15703 5896 15715 5899
rect 16850 5896 16856 5908
rect 15703 5868 16856 5896
rect 15703 5865 15715 5868
rect 15657 5859 15715 5865
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 17126 5856 17132 5908
rect 17184 5896 17190 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17184 5868 17693 5896
rect 17184 5856 17190 5868
rect 17681 5865 17693 5868
rect 17727 5896 17739 5899
rect 17862 5896 17868 5908
rect 17727 5868 17868 5896
rect 17727 5865 17739 5868
rect 17681 5859 17739 5865
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 19242 5856 19248 5908
rect 19300 5896 19306 5908
rect 19613 5899 19671 5905
rect 19613 5896 19625 5899
rect 19300 5868 19625 5896
rect 19300 5856 19306 5868
rect 19613 5865 19625 5868
rect 19659 5865 19671 5899
rect 19613 5859 19671 5865
rect 20349 5899 20407 5905
rect 20349 5865 20361 5899
rect 20395 5896 20407 5899
rect 20438 5896 20444 5908
rect 20395 5868 20444 5896
rect 20395 5865 20407 5868
rect 20349 5859 20407 5865
rect 20438 5856 20444 5868
rect 20496 5896 20502 5908
rect 20806 5896 20812 5908
rect 20496 5868 20812 5896
rect 20496 5856 20502 5868
rect 20806 5856 20812 5868
rect 20864 5856 20870 5908
rect 20898 5856 20904 5908
rect 20956 5896 20962 5908
rect 21361 5899 21419 5905
rect 21361 5896 21373 5899
rect 20956 5868 21373 5896
rect 20956 5856 20962 5868
rect 21361 5865 21373 5868
rect 21407 5896 21419 5899
rect 22002 5896 22008 5908
rect 21407 5868 22008 5896
rect 21407 5865 21419 5868
rect 21361 5859 21419 5865
rect 22002 5856 22008 5868
rect 22060 5856 22066 5908
rect 23014 5896 23020 5908
rect 22975 5868 23020 5896
rect 23014 5856 23020 5868
rect 23072 5856 23078 5908
rect 24210 5856 24216 5908
rect 24268 5896 24274 5908
rect 24489 5899 24547 5905
rect 24489 5896 24501 5899
rect 24268 5868 24501 5896
rect 24268 5856 24274 5868
rect 24489 5865 24501 5868
rect 24535 5865 24547 5899
rect 25130 5896 25136 5908
rect 25091 5868 25136 5896
rect 24489 5859 24547 5865
rect 25130 5856 25136 5868
rect 25188 5856 25194 5908
rect 25406 5896 25412 5908
rect 25367 5868 25412 5896
rect 25406 5856 25412 5868
rect 25464 5856 25470 5908
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 13725 5831 13783 5837
rect 13725 5828 13737 5831
rect 12584 5800 13737 5828
rect 12584 5788 12590 5800
rect 13725 5797 13737 5800
rect 13771 5828 13783 5831
rect 13814 5828 13820 5840
rect 13771 5800 13820 5828
rect 13771 5797 13783 5800
rect 13725 5791 13783 5797
rect 13814 5788 13820 5800
rect 13872 5788 13878 5840
rect 17218 5788 17224 5840
rect 17276 5828 17282 5840
rect 18478 5831 18536 5837
rect 18478 5828 18490 5831
rect 17276 5800 18490 5828
rect 17276 5788 17282 5800
rect 18478 5797 18490 5800
rect 18524 5828 18536 5831
rect 19058 5828 19064 5840
rect 18524 5800 19064 5828
rect 18524 5797 18536 5800
rect 18478 5791 18536 5797
rect 19058 5788 19064 5800
rect 19116 5788 19122 5840
rect 19518 5788 19524 5840
rect 19576 5828 19582 5840
rect 20530 5828 20536 5840
rect 19576 5800 20536 5828
rect 19576 5788 19582 5800
rect 20530 5788 20536 5800
rect 20588 5828 20594 5840
rect 21910 5828 21916 5840
rect 20588 5800 21916 5828
rect 20588 5788 20594 5800
rect 21910 5788 21916 5800
rect 21968 5828 21974 5840
rect 22830 5828 22836 5840
rect 21968 5800 22836 5828
rect 21968 5788 21974 5800
rect 22830 5788 22836 5800
rect 22888 5828 22894 5840
rect 23376 5831 23434 5837
rect 22888 5800 23152 5828
rect 22888 5788 22894 5800
rect 13170 5720 13176 5772
rect 13228 5760 13234 5772
rect 16022 5769 16028 5772
rect 16016 5760 16028 5769
rect 13228 5732 13952 5760
rect 15983 5732 16028 5760
rect 13228 5720 13234 5732
rect 11330 5692 11336 5704
rect 11291 5664 11336 5692
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 12345 5695 12403 5701
rect 12345 5661 12357 5695
rect 12391 5692 12403 5695
rect 12434 5692 12440 5704
rect 12391 5664 12440 5692
rect 12391 5661 12403 5664
rect 12345 5655 12403 5661
rect 12434 5652 12440 5664
rect 12492 5652 12498 5704
rect 13265 5695 13323 5701
rect 13265 5661 13277 5695
rect 13311 5692 13323 5695
rect 13630 5692 13636 5704
rect 13311 5664 13636 5692
rect 13311 5661 13323 5664
rect 13265 5655 13323 5661
rect 13630 5652 13636 5664
rect 13688 5692 13694 5704
rect 13924 5701 13952 5732
rect 16016 5723 16028 5732
rect 16022 5720 16028 5723
rect 16080 5720 16086 5772
rect 18230 5760 18236 5772
rect 18143 5732 18236 5760
rect 18230 5720 18236 5732
rect 18288 5760 18294 5772
rect 19536 5760 19564 5788
rect 18288 5732 19564 5760
rect 18288 5720 18294 5732
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 23124 5769 23152 5800
rect 23376 5797 23388 5831
rect 23422 5828 23434 5831
rect 23566 5828 23572 5840
rect 23422 5800 23572 5828
rect 23422 5797 23434 5800
rect 23376 5791 23434 5797
rect 23566 5788 23572 5800
rect 23624 5788 23630 5840
rect 21269 5763 21327 5769
rect 21269 5760 21281 5763
rect 20772 5732 21281 5760
rect 20772 5720 20778 5732
rect 21269 5729 21281 5732
rect 21315 5729 21327 5763
rect 21269 5723 21327 5729
rect 23109 5763 23167 5769
rect 23109 5729 23121 5763
rect 23155 5729 23167 5763
rect 23109 5723 23167 5729
rect 13817 5695 13875 5701
rect 13817 5692 13829 5695
rect 13688 5664 13829 5692
rect 13688 5652 13694 5664
rect 13817 5661 13829 5664
rect 13863 5661 13875 5695
rect 13817 5655 13875 5661
rect 13909 5695 13967 5701
rect 13909 5661 13921 5695
rect 13955 5661 13967 5695
rect 15749 5695 15807 5701
rect 15749 5692 15761 5695
rect 13909 5655 13967 5661
rect 14752 5664 15761 5692
rect 12253 5627 12311 5633
rect 12253 5593 12265 5627
rect 12299 5624 12311 5627
rect 12618 5624 12624 5636
rect 12299 5596 12624 5624
rect 12299 5593 12311 5596
rect 12253 5587 12311 5593
rect 12618 5584 12624 5596
rect 12676 5624 12682 5636
rect 12676 5596 14504 5624
rect 12676 5584 12682 5596
rect 13078 5516 13084 5568
rect 13136 5556 13142 5568
rect 14476 5565 14504 5596
rect 14752 5568 14780 5664
rect 15749 5661 15761 5664
rect 15795 5661 15807 5695
rect 15749 5655 15807 5661
rect 21358 5652 21364 5704
rect 21416 5692 21422 5704
rect 21453 5695 21511 5701
rect 21453 5692 21465 5695
rect 21416 5664 21465 5692
rect 21416 5652 21422 5664
rect 21453 5661 21465 5664
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 20530 5584 20536 5636
rect 20588 5624 20594 5636
rect 20717 5627 20775 5633
rect 20717 5624 20729 5627
rect 20588 5596 20729 5624
rect 20588 5584 20594 5596
rect 20717 5593 20729 5596
rect 20763 5624 20775 5627
rect 21542 5624 21548 5636
rect 20763 5596 21548 5624
rect 20763 5593 20775 5596
rect 20717 5587 20775 5593
rect 21542 5584 21548 5596
rect 21600 5584 21606 5636
rect 13357 5559 13415 5565
rect 13357 5556 13369 5559
rect 13136 5528 13369 5556
rect 13136 5516 13142 5528
rect 13357 5525 13369 5528
rect 13403 5525 13415 5559
rect 13357 5519 13415 5525
rect 14461 5559 14519 5565
rect 14461 5525 14473 5559
rect 14507 5556 14519 5559
rect 14734 5556 14740 5568
rect 14507 5528 14740 5556
rect 14507 5525 14519 5528
rect 14461 5519 14519 5525
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 15930 5516 15936 5568
rect 15988 5556 15994 5568
rect 17129 5559 17187 5565
rect 17129 5556 17141 5559
rect 15988 5528 17141 5556
rect 15988 5516 15994 5528
rect 17129 5525 17141 5528
rect 17175 5556 17187 5559
rect 17218 5556 17224 5568
rect 17175 5528 17224 5556
rect 17175 5525 17187 5528
rect 17129 5519 17187 5525
rect 17218 5516 17224 5528
rect 17276 5516 17282 5568
rect 18141 5559 18199 5565
rect 18141 5525 18153 5559
rect 18187 5556 18199 5559
rect 18506 5556 18512 5568
rect 18187 5528 18512 5556
rect 18187 5525 18199 5528
rect 18141 5519 18199 5525
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 20898 5556 20904 5568
rect 20859 5528 20904 5556
rect 20898 5516 20904 5528
rect 20956 5516 20962 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 13814 5352 13820 5364
rect 13775 5324 13820 5352
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 14182 5352 14188 5364
rect 14143 5324 14188 5352
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 15657 5355 15715 5361
rect 15657 5321 15669 5355
rect 15703 5352 15715 5355
rect 16022 5352 16028 5364
rect 15703 5324 16028 5352
rect 15703 5321 15715 5324
rect 15657 5315 15715 5321
rect 16022 5312 16028 5324
rect 16080 5352 16086 5364
rect 16209 5355 16267 5361
rect 16209 5352 16221 5355
rect 16080 5324 16221 5352
rect 16080 5312 16086 5324
rect 16209 5321 16221 5324
rect 16255 5321 16267 5355
rect 16209 5315 16267 5321
rect 16761 5355 16819 5361
rect 16761 5321 16773 5355
rect 16807 5352 16819 5355
rect 16850 5352 16856 5364
rect 16807 5324 16856 5352
rect 16807 5321 16819 5324
rect 16761 5315 16819 5321
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 13265 5219 13323 5225
rect 13265 5216 13277 5219
rect 12299 5188 13277 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 13265 5185 13277 5188
rect 13311 5216 13323 5219
rect 14200 5216 14228 5312
rect 16224 5284 16252 5315
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 18049 5355 18107 5361
rect 18049 5352 18061 5355
rect 18012 5324 18061 5352
rect 18012 5312 18018 5324
rect 18049 5321 18061 5324
rect 18095 5321 18107 5355
rect 19058 5352 19064 5364
rect 19019 5324 19064 5352
rect 18049 5315 18107 5321
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 21269 5355 21327 5361
rect 21269 5321 21281 5355
rect 21315 5352 21327 5355
rect 21358 5352 21364 5364
rect 21315 5324 21364 5352
rect 21315 5321 21327 5324
rect 21269 5315 21327 5321
rect 21358 5312 21364 5324
rect 21416 5352 21422 5364
rect 21821 5355 21879 5361
rect 21821 5352 21833 5355
rect 21416 5324 21833 5352
rect 21416 5312 21422 5324
rect 21821 5321 21833 5324
rect 21867 5321 21879 5355
rect 21821 5315 21879 5321
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 22189 5355 22247 5361
rect 22189 5352 22201 5355
rect 22152 5324 22201 5352
rect 22152 5312 22158 5324
rect 22189 5321 22201 5324
rect 22235 5321 22247 5355
rect 22189 5315 22247 5321
rect 22738 5312 22744 5364
rect 22796 5352 22802 5364
rect 23017 5355 23075 5361
rect 23017 5352 23029 5355
rect 22796 5324 23029 5352
rect 22796 5312 22802 5324
rect 23017 5321 23029 5324
rect 23063 5321 23075 5355
rect 23017 5315 23075 5321
rect 23477 5355 23535 5361
rect 23477 5321 23489 5355
rect 23523 5352 23535 5355
rect 23566 5352 23572 5364
rect 23523 5324 23572 5352
rect 23523 5321 23535 5324
rect 23477 5315 23535 5321
rect 23566 5312 23572 5324
rect 23624 5312 23630 5364
rect 23661 5355 23719 5361
rect 23661 5321 23673 5355
rect 23707 5352 23719 5355
rect 24762 5352 24768 5364
rect 23707 5324 24768 5352
rect 23707 5321 23719 5324
rect 23661 5315 23719 5321
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 17405 5287 17463 5293
rect 17405 5284 17417 5287
rect 16224 5256 17417 5284
rect 17405 5253 17417 5256
rect 17451 5284 17463 5287
rect 25041 5287 25099 5293
rect 25041 5284 25053 5287
rect 17451 5256 18552 5284
rect 17451 5253 17463 5256
rect 17405 5247 17463 5253
rect 13311 5188 14412 5216
rect 13311 5185 13323 5188
rect 13265 5179 13323 5185
rect 11885 5151 11943 5157
rect 11885 5117 11897 5151
rect 11931 5148 11943 5151
rect 13078 5148 13084 5160
rect 11931 5120 13084 5148
rect 11931 5117 11943 5120
rect 11885 5111 11943 5117
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13173 5151 13231 5157
rect 13173 5117 13185 5151
rect 13219 5148 13231 5151
rect 13354 5148 13360 5160
rect 13219 5120 13360 5148
rect 13219 5117 13231 5120
rect 13173 5111 13231 5117
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 14277 5151 14335 5157
rect 14277 5117 14289 5151
rect 14323 5117 14335 5151
rect 14384 5148 14412 5188
rect 14533 5151 14591 5157
rect 14533 5148 14545 5151
rect 14384 5120 14545 5148
rect 14277 5111 14335 5117
rect 14533 5117 14545 5120
rect 14579 5117 14591 5151
rect 16850 5148 16856 5160
rect 16811 5120 16856 5148
rect 14533 5111 14591 5117
rect 14292 5080 14320 5111
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 17865 5151 17923 5157
rect 17865 5117 17877 5151
rect 17911 5148 17923 5151
rect 18414 5148 18420 5160
rect 17911 5120 18420 5148
rect 17911 5117 17923 5120
rect 17865 5111 17923 5117
rect 18414 5108 18420 5120
rect 18472 5108 18478 5160
rect 18524 5148 18552 5256
rect 24136 5256 25053 5284
rect 18690 5176 18696 5228
rect 18748 5216 18754 5228
rect 19797 5219 19855 5225
rect 18748 5188 18841 5216
rect 18748 5176 18754 5188
rect 19797 5185 19809 5219
rect 19843 5216 19855 5219
rect 19843 5188 20024 5216
rect 19843 5185 19855 5188
rect 19797 5179 19855 5185
rect 18708 5148 18736 5176
rect 18524 5120 18736 5148
rect 19518 5108 19524 5160
rect 19576 5148 19582 5160
rect 19889 5151 19947 5157
rect 19889 5148 19901 5151
rect 19576 5120 19901 5148
rect 19576 5108 19582 5120
rect 19889 5117 19901 5120
rect 19935 5117 19947 5151
rect 19996 5148 20024 5188
rect 24026 5176 24032 5228
rect 24084 5216 24090 5228
rect 24136 5225 24164 5256
rect 25041 5253 25053 5256
rect 25087 5253 25099 5287
rect 25041 5247 25099 5253
rect 25409 5287 25467 5293
rect 25409 5253 25421 5287
rect 25455 5284 25467 5287
rect 26878 5284 26884 5296
rect 25455 5256 26884 5284
rect 25455 5253 25467 5256
rect 25409 5247 25467 5253
rect 26878 5244 26884 5256
rect 26936 5244 26942 5296
rect 24121 5219 24179 5225
rect 24121 5216 24133 5219
rect 24084 5188 24133 5216
rect 24084 5176 24090 5188
rect 24121 5185 24133 5188
rect 24167 5185 24179 5219
rect 24121 5179 24179 5185
rect 24305 5219 24363 5225
rect 24305 5185 24317 5219
rect 24351 5216 24363 5219
rect 24670 5216 24676 5228
rect 24351 5188 24676 5216
rect 24351 5185 24363 5188
rect 24305 5179 24363 5185
rect 24670 5176 24676 5188
rect 24728 5176 24734 5228
rect 20156 5151 20214 5157
rect 20156 5148 20168 5151
rect 19996 5120 20168 5148
rect 19889 5111 19947 5117
rect 20156 5117 20168 5120
rect 20202 5148 20214 5151
rect 20530 5148 20536 5160
rect 20202 5120 20536 5148
rect 20202 5117 20214 5120
rect 20156 5111 20214 5117
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 22465 5151 22523 5157
rect 22465 5117 22477 5151
rect 22511 5148 22523 5151
rect 22738 5148 22744 5160
rect 22511 5120 22744 5148
rect 22511 5117 22523 5120
rect 22465 5111 22523 5117
rect 22738 5108 22744 5120
rect 22796 5108 22802 5160
rect 25222 5148 25228 5160
rect 25183 5120 25228 5148
rect 25222 5108 25228 5120
rect 25280 5148 25286 5160
rect 25777 5151 25835 5157
rect 25777 5148 25789 5151
rect 25280 5120 25789 5148
rect 25280 5108 25286 5120
rect 25777 5117 25789 5120
rect 25823 5117 25835 5151
rect 25777 5111 25835 5117
rect 14734 5080 14740 5092
rect 14292 5052 14740 5080
rect 14734 5040 14740 5052
rect 14792 5040 14798 5092
rect 24029 5083 24087 5089
rect 24029 5049 24041 5083
rect 24075 5080 24087 5083
rect 24118 5080 24124 5092
rect 24075 5052 24124 5080
rect 24075 5049 24087 5052
rect 24029 5043 24087 5049
rect 24118 5040 24124 5052
rect 24176 5040 24182 5092
rect 11330 5012 11336 5024
rect 11291 4984 11336 5012
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 12713 5015 12771 5021
rect 12713 4981 12725 5015
rect 12759 5012 12771 5015
rect 12802 5012 12808 5024
rect 12759 4984 12808 5012
rect 12759 4981 12771 4984
rect 12713 4975 12771 4981
rect 12802 4972 12808 4984
rect 12860 4972 12866 5024
rect 17034 5012 17040 5024
rect 16995 4984 17040 5012
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 18046 4972 18052 5024
rect 18104 5012 18110 5024
rect 18509 5015 18567 5021
rect 18509 5012 18521 5015
rect 18104 4984 18521 5012
rect 18104 4972 18110 4984
rect 18509 4981 18521 4984
rect 18555 4981 18567 5015
rect 22646 5012 22652 5024
rect 22607 4984 22652 5012
rect 18509 4975 18567 4981
rect 22646 4972 22652 4984
rect 22704 4972 22710 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 12894 4808 12900 4820
rect 12492 4780 12900 4808
rect 12492 4768 12498 4780
rect 12894 4768 12900 4780
rect 12952 4808 12958 4820
rect 13081 4811 13139 4817
rect 13081 4808 13093 4811
rect 12952 4780 13093 4808
rect 12952 4768 12958 4780
rect 13081 4777 13093 4780
rect 13127 4777 13139 4811
rect 13081 4771 13139 4777
rect 13170 4768 13176 4820
rect 13228 4808 13234 4820
rect 13449 4811 13507 4817
rect 13449 4808 13461 4811
rect 13228 4780 13461 4808
rect 13228 4768 13234 4780
rect 13449 4777 13461 4780
rect 13495 4777 13507 4811
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 13449 4771 13507 4777
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 13998 4768 14004 4820
rect 14056 4808 14062 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 14056 4780 14105 4808
rect 14056 4768 14062 4780
rect 14093 4777 14105 4780
rect 14139 4808 14151 4811
rect 14366 4808 14372 4820
rect 14139 4780 14372 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 16390 4808 16396 4820
rect 16351 4780 16396 4808
rect 16390 4768 16396 4780
rect 16448 4768 16454 4820
rect 16761 4811 16819 4817
rect 16761 4777 16773 4811
rect 16807 4808 16819 4811
rect 17313 4811 17371 4817
rect 17313 4808 17325 4811
rect 16807 4780 17325 4808
rect 16807 4777 16819 4780
rect 16761 4771 16819 4777
rect 17313 4777 17325 4780
rect 17359 4808 17371 4811
rect 17770 4808 17776 4820
rect 17359 4780 17776 4808
rect 17359 4777 17371 4780
rect 17313 4771 17371 4777
rect 17770 4768 17776 4780
rect 17828 4768 17834 4820
rect 18046 4808 18052 4820
rect 18007 4780 18052 4808
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 19242 4808 19248 4820
rect 19203 4780 19248 4808
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 20530 4768 20536 4820
rect 20588 4808 20594 4820
rect 20714 4808 20720 4820
rect 20588 4780 20720 4808
rect 20588 4768 20594 4780
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 20806 4768 20812 4820
rect 20864 4808 20870 4820
rect 20901 4811 20959 4817
rect 20901 4808 20913 4811
rect 20864 4780 20913 4808
rect 20864 4768 20870 4780
rect 20901 4777 20913 4780
rect 20947 4777 20959 4811
rect 20901 4771 20959 4777
rect 21082 4768 21088 4820
rect 21140 4808 21146 4820
rect 21361 4811 21419 4817
rect 21361 4808 21373 4811
rect 21140 4780 21373 4808
rect 21140 4768 21146 4780
rect 21361 4777 21373 4780
rect 21407 4777 21419 4811
rect 21361 4771 21419 4777
rect 22097 4811 22155 4817
rect 22097 4777 22109 4811
rect 22143 4808 22155 4811
rect 22554 4808 22560 4820
rect 22143 4780 22560 4808
rect 22143 4777 22155 4780
rect 22097 4771 22155 4777
rect 22554 4768 22560 4780
rect 22612 4768 22618 4820
rect 22830 4808 22836 4820
rect 22791 4780 22836 4808
rect 22830 4768 22836 4780
rect 22888 4768 22894 4820
rect 23566 4768 23572 4820
rect 23624 4808 23630 4820
rect 24210 4808 24216 4820
rect 23624 4780 24216 4808
rect 23624 4768 23630 4780
rect 24210 4768 24216 4780
rect 24268 4808 24274 4820
rect 24673 4811 24731 4817
rect 24673 4808 24685 4811
rect 24268 4780 24685 4808
rect 24268 4768 24274 4780
rect 24673 4777 24685 4780
rect 24719 4777 24731 4811
rect 24673 4771 24731 4777
rect 12529 4743 12587 4749
rect 12529 4709 12541 4743
rect 12575 4740 12587 4743
rect 13262 4740 13268 4752
rect 12575 4712 13268 4740
rect 12575 4709 12587 4712
rect 12529 4703 12587 4709
rect 13262 4700 13268 4712
rect 13320 4700 13326 4752
rect 15838 4700 15844 4752
rect 15896 4740 15902 4752
rect 17221 4743 17279 4749
rect 17221 4740 17233 4743
rect 15896 4712 17233 4740
rect 15896 4700 15902 4712
rect 17221 4709 17233 4712
rect 17267 4709 17279 4743
rect 17221 4703 17279 4709
rect 12158 4632 12164 4684
rect 12216 4672 12222 4684
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 12216 4644 12449 4672
rect 12216 4632 12222 4644
rect 12437 4641 12449 4644
rect 12483 4641 12495 4675
rect 12437 4635 12495 4641
rect 13814 4632 13820 4684
rect 13872 4672 13878 4684
rect 14001 4675 14059 4681
rect 14001 4672 14013 4675
rect 13872 4644 14013 4672
rect 13872 4632 13878 4644
rect 14001 4641 14013 4644
rect 14047 4641 14059 4675
rect 14001 4635 14059 4641
rect 15378 4632 15384 4684
rect 15436 4672 15442 4684
rect 15749 4675 15807 4681
rect 15749 4672 15761 4675
rect 15436 4644 15761 4672
rect 15436 4632 15442 4644
rect 15749 4641 15761 4644
rect 15795 4672 15807 4675
rect 16022 4672 16028 4684
rect 15795 4644 16028 4672
rect 15795 4641 15807 4644
rect 15749 4635 15807 4641
rect 16022 4632 16028 4644
rect 16080 4632 16086 4684
rect 18417 4675 18475 4681
rect 18417 4641 18429 4675
rect 18463 4672 18475 4675
rect 19260 4672 19288 4768
rect 18463 4644 19288 4672
rect 19705 4675 19763 4681
rect 18463 4641 18475 4644
rect 18417 4635 18475 4641
rect 19705 4641 19717 4675
rect 19751 4672 19763 4675
rect 19978 4672 19984 4684
rect 19751 4644 19984 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 20806 4632 20812 4684
rect 20864 4672 20870 4684
rect 21269 4675 21327 4681
rect 21269 4672 21281 4675
rect 20864 4644 21281 4672
rect 20864 4632 20870 4644
rect 21269 4641 21281 4644
rect 21315 4641 21327 4675
rect 22848 4672 22876 4768
rect 23201 4743 23259 4749
rect 23201 4709 23213 4743
rect 23247 4740 23259 4743
rect 24118 4740 24124 4752
rect 23247 4712 24124 4740
rect 23247 4709 23259 4712
rect 23201 4703 23259 4709
rect 24118 4700 24124 4712
rect 24176 4700 24182 4752
rect 23290 4672 23296 4684
rect 22848 4644 23296 4672
rect 21269 4635 21327 4641
rect 23290 4632 23296 4644
rect 23348 4632 23354 4684
rect 23382 4632 23388 4684
rect 23440 4672 23446 4684
rect 23549 4675 23607 4681
rect 23549 4672 23561 4675
rect 23440 4644 23561 4672
rect 23440 4632 23446 4644
rect 23549 4641 23561 4644
rect 23595 4641 23607 4675
rect 23549 4635 23607 4641
rect 12710 4604 12716 4616
rect 12671 4576 12716 4604
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 17218 4564 17224 4616
rect 17276 4604 17282 4616
rect 17405 4607 17463 4613
rect 17405 4604 17417 4607
rect 17276 4576 17417 4604
rect 17276 4564 17282 4576
rect 17405 4573 17417 4576
rect 17451 4573 17463 4607
rect 18598 4604 18604 4616
rect 18559 4576 18604 4604
rect 17405 4567 17463 4573
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 21450 4564 21456 4616
rect 21508 4604 21514 4616
rect 21508 4576 21553 4604
rect 21508 4564 21514 4576
rect 11977 4539 12035 4545
rect 11977 4505 11989 4539
rect 12023 4536 12035 4539
rect 13078 4536 13084 4548
rect 12023 4508 13084 4536
rect 12023 4505 12035 4508
rect 11977 4499 12035 4505
rect 13078 4496 13084 4508
rect 13136 4496 13142 4548
rect 15930 4536 15936 4548
rect 15891 4508 15936 4536
rect 15930 4496 15936 4508
rect 15988 4496 15994 4548
rect 16758 4496 16764 4548
rect 16816 4536 16822 4548
rect 16853 4539 16911 4545
rect 16853 4536 16865 4539
rect 16816 4508 16865 4536
rect 16816 4496 16822 4508
rect 16853 4505 16865 4508
rect 16899 4505 16911 4539
rect 20257 4539 20315 4545
rect 20257 4536 20269 4539
rect 16853 4499 16911 4505
rect 19536 4508 20269 4536
rect 19536 4480 19564 4508
rect 20257 4505 20269 4508
rect 20303 4505 20315 4539
rect 20257 4499 20315 4505
rect 11333 4471 11391 4477
rect 11333 4437 11345 4471
rect 11379 4468 11391 4471
rect 11422 4468 11428 4480
rect 11379 4440 11428 4468
rect 11379 4437 11391 4440
rect 11333 4431 11391 4437
rect 11422 4428 11428 4440
rect 11480 4428 11486 4480
rect 12066 4468 12072 4480
rect 12027 4440 12072 4468
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 14734 4468 14740 4480
rect 14647 4440 14740 4468
rect 14734 4428 14740 4440
rect 14792 4468 14798 4480
rect 15013 4471 15071 4477
rect 15013 4468 15025 4471
rect 14792 4440 15025 4468
rect 14792 4428 14798 4440
rect 15013 4437 15025 4440
rect 15059 4468 15071 4471
rect 15378 4468 15384 4480
rect 15059 4440 15384 4468
rect 15059 4437 15071 4440
rect 15013 4431 15071 4437
rect 15378 4428 15384 4440
rect 15436 4468 15442 4480
rect 15565 4471 15623 4477
rect 15565 4468 15577 4471
rect 15436 4440 15577 4468
rect 15436 4428 15442 4440
rect 15565 4437 15577 4440
rect 15611 4437 15623 4471
rect 19518 4468 19524 4480
rect 19479 4440 19524 4468
rect 15565 4431 15623 4437
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 19889 4471 19947 4477
rect 19889 4437 19901 4471
rect 19935 4468 19947 4471
rect 20070 4468 20076 4480
rect 19935 4440 20076 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 22462 4468 22468 4480
rect 22423 4440 22468 4468
rect 22462 4428 22468 4440
rect 22520 4428 22526 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 14274 4224 14280 4276
rect 14332 4264 14338 4276
rect 14737 4267 14795 4273
rect 14737 4264 14749 4267
rect 14332 4236 14749 4264
rect 14332 4224 14338 4236
rect 14737 4233 14749 4236
rect 14783 4233 14795 4267
rect 16022 4264 16028 4276
rect 15983 4236 16028 4264
rect 14737 4227 14795 4233
rect 16022 4224 16028 4236
rect 16080 4224 16086 4276
rect 19705 4267 19763 4273
rect 19705 4233 19717 4267
rect 19751 4264 19763 4267
rect 19978 4264 19984 4276
rect 19751 4236 19984 4264
rect 19751 4233 19763 4236
rect 19705 4227 19763 4233
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 20806 4224 20812 4276
rect 20864 4264 20870 4276
rect 20901 4267 20959 4273
rect 20901 4264 20913 4267
rect 20864 4236 20913 4264
rect 20864 4224 20870 4236
rect 20901 4233 20913 4236
rect 20947 4233 20959 4267
rect 20901 4227 20959 4233
rect 21082 4224 21088 4276
rect 21140 4264 21146 4276
rect 21269 4267 21327 4273
rect 21269 4264 21281 4267
rect 21140 4236 21281 4264
rect 21140 4224 21146 4236
rect 21269 4233 21281 4236
rect 21315 4233 21327 4267
rect 21269 4227 21327 4233
rect 23474 4224 23480 4276
rect 23532 4264 23538 4276
rect 23661 4267 23719 4273
rect 23661 4264 23673 4267
rect 23532 4236 23673 4264
rect 23532 4224 23538 4236
rect 23661 4233 23673 4236
rect 23707 4233 23719 4267
rect 23661 4227 23719 4233
rect 21634 4156 21640 4208
rect 21692 4196 21698 4208
rect 21821 4199 21879 4205
rect 21821 4196 21833 4199
rect 21692 4168 21833 4196
rect 21692 4156 21698 4168
rect 21821 4165 21833 4168
rect 21867 4196 21879 4199
rect 22278 4196 22284 4208
rect 21867 4168 22284 4196
rect 21867 4165 21879 4168
rect 21821 4159 21879 4165
rect 22278 4156 22284 4168
rect 22336 4156 22342 4208
rect 22462 4156 22468 4208
rect 22520 4196 22526 4208
rect 23109 4199 23167 4205
rect 23109 4196 23121 4199
rect 22520 4168 23121 4196
rect 22520 4156 22526 4168
rect 9122 4088 9128 4140
rect 9180 4128 9186 4140
rect 9674 4128 9680 4140
rect 9180 4100 9680 4128
rect 9180 4088 9186 4100
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 12066 4088 12072 4140
rect 12124 4128 12130 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12124 4100 12909 4128
rect 12124 4088 12130 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 13078 4128 13084 4140
rect 13039 4100 13084 4128
rect 12897 4091 12955 4097
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 13630 4128 13636 4140
rect 13591 4100 13636 4128
rect 13630 4088 13636 4100
rect 13688 4088 13694 4140
rect 14277 4131 14335 4137
rect 14277 4097 14289 4131
rect 14323 4128 14335 4131
rect 14458 4128 14464 4140
rect 14323 4100 14464 4128
rect 14323 4097 14335 4100
rect 14277 4091 14335 4097
rect 14458 4088 14464 4100
rect 14516 4088 14522 4140
rect 15286 4128 15292 4140
rect 15247 4100 15292 4128
rect 15286 4088 15292 4100
rect 15344 4128 15350 4140
rect 15344 4100 15424 4128
rect 15344 4088 15350 4100
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4060 11299 4063
rect 11422 4060 11428 4072
rect 11287 4032 11428 4060
rect 11287 4029 11299 4032
rect 11241 4023 11299 4029
rect 11422 4020 11428 4032
rect 11480 4060 11486 4072
rect 12342 4060 12348 4072
rect 11480 4032 12348 4060
rect 11480 4020 11486 4032
rect 12342 4020 12348 4032
rect 12400 4020 12406 4072
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 12452 4032 14013 4060
rect 11149 3927 11207 3933
rect 11149 3893 11161 3927
rect 11195 3924 11207 3927
rect 11238 3924 11244 3936
rect 11195 3896 11244 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 11422 3924 11428 3936
rect 11383 3896 11428 3924
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 11790 3884 11796 3936
rect 11848 3924 11854 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 11848 3896 12081 3924
rect 11848 3884 11854 3896
rect 12069 3893 12081 3896
rect 12115 3924 12127 3927
rect 12158 3924 12164 3936
rect 12115 3896 12164 3924
rect 12115 3893 12127 3896
rect 12069 3887 12127 3893
rect 12158 3884 12164 3896
rect 12216 3884 12222 3936
rect 12452 3933 12480 4032
rect 14001 4029 14013 4032
rect 14047 4060 14059 4063
rect 14366 4060 14372 4072
rect 14047 4032 14372 4060
rect 14047 4029 14059 4032
rect 14001 4023 14059 4029
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 15396 4069 15424 4100
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16356 4100 16681 4128
rect 16356 4088 16362 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 17678 4088 17684 4140
rect 17736 4128 17742 4140
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 17736 4100 17785 4128
rect 17736 4088 17742 4100
rect 17773 4097 17785 4100
rect 17819 4128 17831 4131
rect 18782 4128 18788 4140
rect 17819 4100 18644 4128
rect 18743 4100 18788 4128
rect 17819 4097 17831 4100
rect 17773 4091 17831 4097
rect 15381 4063 15439 4069
rect 15381 4029 15393 4063
rect 15427 4029 15439 4063
rect 15381 4023 15439 4029
rect 16390 4020 16396 4072
rect 16448 4060 16454 4072
rect 18616 4069 18644 4100
rect 18782 4088 18788 4100
rect 18840 4088 18846 4140
rect 19337 4131 19395 4137
rect 19337 4097 19349 4131
rect 19383 4128 19395 4131
rect 20438 4128 20444 4140
rect 19383 4100 20444 4128
rect 19383 4097 19395 4100
rect 19337 4091 19395 4097
rect 20438 4088 20444 4100
rect 20496 4088 20502 4140
rect 22664 4137 22692 4168
rect 23109 4165 23121 4168
rect 23155 4196 23167 4199
rect 23382 4196 23388 4208
rect 23155 4168 23388 4196
rect 23155 4165 23167 4168
rect 23109 4159 23167 4165
rect 23382 4156 23388 4168
rect 23440 4196 23446 4208
rect 23440 4168 24900 4196
rect 23440 4156 23446 4168
rect 22649 4131 22707 4137
rect 22649 4097 22661 4131
rect 22695 4097 22707 4131
rect 22649 4091 22707 4097
rect 23290 4088 23296 4140
rect 23348 4128 23354 4140
rect 24302 4128 24308 4140
rect 23348 4100 24164 4128
rect 24263 4100 24308 4128
rect 23348 4088 23354 4100
rect 16485 4063 16543 4069
rect 16485 4060 16497 4063
rect 16448 4032 16497 4060
rect 16448 4020 16454 4032
rect 16485 4029 16497 4032
rect 16531 4029 16543 4063
rect 16485 4023 16543 4029
rect 18601 4063 18659 4069
rect 18601 4029 18613 4063
rect 18647 4029 18659 4063
rect 20254 4060 20260 4072
rect 20167 4032 20260 4060
rect 18601 4023 18659 4029
rect 20254 4020 20260 4032
rect 20312 4060 20318 4072
rect 20622 4060 20628 4072
rect 20312 4032 20628 4060
rect 20312 4020 20318 4032
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 22465 4063 22523 4069
rect 22465 4029 22477 4063
rect 22511 4060 22523 4063
rect 22554 4060 22560 4072
rect 22511 4032 22560 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 22554 4020 22560 4032
rect 22612 4060 22618 4072
rect 23382 4060 23388 4072
rect 22612 4032 23388 4060
rect 22612 4020 22618 4032
rect 23382 4020 23388 4032
rect 23440 4020 23446 4072
rect 23477 4063 23535 4069
rect 23477 4029 23489 4063
rect 23523 4060 23535 4063
rect 24026 4060 24032 4072
rect 23523 4032 24032 4060
rect 23523 4029 23535 4032
rect 23477 4023 23535 4029
rect 24026 4020 24032 4032
rect 24084 4020 24090 4072
rect 24136 4060 24164 4100
rect 24302 4088 24308 4100
rect 24360 4088 24366 4140
rect 24872 4128 24900 4168
rect 24946 4128 24952 4140
rect 24872 4100 24952 4128
rect 24946 4088 24952 4100
rect 25004 4088 25010 4140
rect 25038 4060 25044 4072
rect 24136 4032 25044 4060
rect 25038 4020 25044 4032
rect 25096 4020 25102 4072
rect 25225 4063 25283 4069
rect 25225 4029 25237 4063
rect 25271 4060 25283 4063
rect 25314 4060 25320 4072
rect 25271 4032 25320 4060
rect 25271 4029 25283 4032
rect 25225 4023 25283 4029
rect 25314 4020 25320 4032
rect 25372 4060 25378 4072
rect 25777 4063 25835 4069
rect 25777 4060 25789 4063
rect 25372 4032 25789 4060
rect 25372 4020 25378 4032
rect 25777 4029 25789 4032
rect 25823 4029 25835 4063
rect 25777 4023 25835 4029
rect 12805 3995 12863 4001
rect 12805 3961 12817 3995
rect 12851 3992 12863 3995
rect 12894 3992 12900 4004
rect 12851 3964 12900 3992
rect 12851 3961 12863 3964
rect 12805 3955 12863 3961
rect 12894 3952 12900 3964
rect 12952 3952 12958 4004
rect 15838 3952 15844 4004
rect 15896 3992 15902 4004
rect 16301 3995 16359 4001
rect 16301 3992 16313 3995
rect 15896 3964 16313 3992
rect 15896 3952 15902 3964
rect 16301 3961 16313 3964
rect 16347 3961 16359 3995
rect 16301 3955 16359 3961
rect 17497 3995 17555 4001
rect 17497 3961 17509 3995
rect 17543 3992 17555 3995
rect 20530 3992 20536 4004
rect 17543 3964 18736 3992
rect 17543 3961 17555 3964
rect 17497 3955 17555 3961
rect 18708 3936 18736 3964
rect 19812 3964 20536 3992
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3893 12495 3927
rect 12437 3887 12495 3893
rect 12526 3884 12532 3936
rect 12584 3924 12590 3936
rect 13446 3924 13452 3936
rect 12584 3896 13452 3924
rect 12584 3884 12590 3896
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 15562 3924 15568 3936
rect 15523 3896 15568 3924
rect 15562 3884 15568 3896
rect 15620 3884 15626 3936
rect 18230 3924 18236 3936
rect 18191 3896 18236 3924
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 18690 3924 18696 3936
rect 18651 3896 18696 3924
rect 18690 3884 18696 3896
rect 18748 3884 18754 3936
rect 19812 3933 19840 3964
rect 20530 3952 20536 3964
rect 20588 3952 20594 4004
rect 24121 3995 24179 4001
rect 24121 3992 24133 3995
rect 22020 3964 24133 3992
rect 19797 3927 19855 3933
rect 19797 3893 19809 3927
rect 19843 3893 19855 3927
rect 19797 3887 19855 3893
rect 19978 3884 19984 3936
rect 20036 3924 20042 3936
rect 22020 3933 22048 3964
rect 24121 3961 24133 3964
rect 24167 3992 24179 3995
rect 24673 3995 24731 4001
rect 24673 3992 24685 3995
rect 24167 3964 24685 3992
rect 24167 3961 24179 3964
rect 24121 3955 24179 3961
rect 24673 3961 24685 3964
rect 24719 3961 24731 3995
rect 24673 3955 24731 3961
rect 20165 3927 20223 3933
rect 20165 3924 20177 3927
rect 20036 3896 20177 3924
rect 20036 3884 20042 3896
rect 20165 3893 20177 3896
rect 20211 3893 20223 3927
rect 20165 3887 20223 3893
rect 22005 3927 22063 3933
rect 22005 3893 22017 3927
rect 22051 3893 22063 3927
rect 22005 3887 22063 3893
rect 22278 3884 22284 3936
rect 22336 3924 22342 3936
rect 22373 3927 22431 3933
rect 22373 3924 22385 3927
rect 22336 3896 22385 3924
rect 22336 3884 22342 3896
rect 22373 3893 22385 3896
rect 22419 3893 22431 3927
rect 24026 3924 24032 3936
rect 23939 3896 24032 3924
rect 22373 3887 22431 3893
rect 24026 3884 24032 3896
rect 24084 3924 24090 3936
rect 24762 3924 24768 3936
rect 24084 3896 24768 3924
rect 24084 3884 24090 3896
rect 24762 3884 24768 3896
rect 24820 3884 24826 3936
rect 25406 3924 25412 3936
rect 25367 3896 25412 3924
rect 25406 3884 25412 3896
rect 25464 3884 25470 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 11146 3720 11152 3732
rect 11107 3692 11152 3720
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 11609 3723 11667 3729
rect 11609 3689 11621 3723
rect 11655 3720 11667 3723
rect 12066 3720 12072 3732
rect 11655 3692 12072 3720
rect 11655 3689 11667 3692
rect 11609 3683 11667 3689
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 13078 3680 13084 3732
rect 13136 3720 13142 3732
rect 13446 3720 13452 3732
rect 13136 3692 13452 3720
rect 13136 3680 13142 3692
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 13998 3720 14004 3732
rect 13959 3692 14004 3720
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 14366 3720 14372 3732
rect 14327 3692 14372 3720
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 17218 3720 17224 3732
rect 17179 3692 17224 3720
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 19334 3680 19340 3732
rect 19392 3720 19398 3732
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 19392 3692 19809 3720
rect 19392 3680 19398 3692
rect 19797 3689 19809 3692
rect 19843 3720 19855 3723
rect 19978 3720 19984 3732
rect 19843 3692 19984 3720
rect 19843 3689 19855 3692
rect 19797 3683 19855 3689
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 20254 3720 20260 3732
rect 20215 3692 20260 3720
rect 20254 3680 20260 3692
rect 20312 3680 20318 3732
rect 21177 3723 21235 3729
rect 21177 3689 21189 3723
rect 21223 3720 21235 3723
rect 21450 3720 21456 3732
rect 21223 3692 21456 3720
rect 21223 3689 21235 3692
rect 21177 3683 21235 3689
rect 21450 3680 21456 3692
rect 21508 3680 21514 3732
rect 23290 3720 23296 3732
rect 23251 3692 23296 3720
rect 23290 3680 23296 3692
rect 23348 3680 23354 3732
rect 23753 3723 23811 3729
rect 23753 3689 23765 3723
rect 23799 3720 23811 3723
rect 24210 3720 24216 3732
rect 23799 3692 24216 3720
rect 23799 3689 23811 3692
rect 23753 3683 23811 3689
rect 24210 3680 24216 3692
rect 24268 3680 24274 3732
rect 24946 3680 24952 3732
rect 25004 3720 25010 3732
rect 25225 3723 25283 3729
rect 25225 3720 25237 3723
rect 25004 3692 25237 3720
rect 25004 3680 25010 3692
rect 25225 3689 25237 3692
rect 25271 3689 25283 3723
rect 25225 3683 25283 3689
rect 11238 3612 11244 3664
rect 11296 3652 11302 3664
rect 12250 3652 12256 3664
rect 11296 3624 12256 3652
rect 11296 3612 11302 3624
rect 12250 3612 12256 3624
rect 12308 3661 12314 3664
rect 12308 3655 12372 3661
rect 12308 3621 12326 3655
rect 12360 3621 12372 3655
rect 12308 3615 12372 3621
rect 12308 3612 12314 3615
rect 12710 3612 12716 3664
rect 12768 3652 12774 3664
rect 13538 3652 13544 3664
rect 12768 3624 13544 3652
rect 12768 3612 12774 3624
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 15286 3612 15292 3664
rect 15344 3652 15350 3664
rect 15534 3655 15592 3661
rect 15534 3652 15546 3655
rect 15344 3624 15546 3652
rect 15344 3612 15350 3624
rect 15534 3621 15546 3624
rect 15580 3621 15592 3655
rect 15534 3615 15592 3621
rect 9861 3587 9919 3593
rect 9861 3553 9873 3587
rect 9907 3584 9919 3587
rect 9950 3584 9956 3596
rect 9907 3556 9956 3584
rect 9907 3553 9919 3556
rect 9861 3547 9919 3553
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3584 11023 3587
rect 11514 3584 11520 3596
rect 11011 3556 11520 3584
rect 11011 3553 11023 3556
rect 10965 3547 11023 3553
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 12069 3587 12127 3593
rect 12069 3553 12081 3587
rect 12115 3584 12127 3587
rect 12618 3584 12624 3596
rect 12115 3556 12624 3584
rect 12115 3553 12127 3556
rect 12069 3547 12127 3553
rect 12618 3544 12624 3556
rect 12676 3584 12682 3596
rect 15378 3584 15384 3596
rect 12676 3556 15384 3584
rect 12676 3544 12682 3556
rect 15304 3525 15332 3556
rect 15378 3544 15384 3556
rect 15436 3544 15442 3596
rect 17494 3544 17500 3596
rect 17552 3584 17558 3596
rect 18029 3587 18087 3593
rect 18029 3584 18041 3587
rect 17552 3556 18041 3584
rect 17552 3544 17558 3556
rect 18029 3553 18041 3556
rect 18075 3553 18087 3587
rect 18029 3547 18087 3553
rect 21628 3587 21686 3593
rect 21628 3553 21640 3587
rect 21674 3584 21686 3587
rect 21910 3584 21916 3596
rect 21674 3556 21916 3584
rect 21674 3553 21686 3556
rect 21628 3547 21686 3553
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 22738 3544 22744 3596
rect 22796 3584 22802 3596
rect 24118 3593 24124 3596
rect 24101 3587 24124 3593
rect 24101 3584 24113 3587
rect 22796 3556 24113 3584
rect 22796 3544 22802 3556
rect 24101 3553 24113 3556
rect 24176 3584 24182 3596
rect 24176 3556 24249 3584
rect 24101 3547 24124 3553
rect 24118 3544 24124 3547
rect 24176 3544 24182 3556
rect 15289 3519 15347 3525
rect 15289 3485 15301 3519
rect 15335 3485 15347 3519
rect 17770 3516 17776 3528
rect 17731 3488 17776 3516
rect 15289 3479 15347 3485
rect 17770 3476 17776 3488
rect 17828 3476 17834 3528
rect 21361 3519 21419 3525
rect 21361 3516 21373 3519
rect 20732 3488 21373 3516
rect 20732 3460 20760 3488
rect 21361 3485 21373 3488
rect 21407 3485 21419 3519
rect 21361 3479 21419 3485
rect 23290 3476 23296 3528
rect 23348 3516 23354 3528
rect 23845 3519 23903 3525
rect 23845 3516 23857 3519
rect 23348 3488 23857 3516
rect 23348 3476 23354 3488
rect 23845 3485 23857 3488
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 10042 3448 10048 3460
rect 10003 3420 10048 3448
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 16669 3451 16727 3457
rect 16669 3417 16681 3451
rect 16715 3448 16727 3451
rect 16758 3448 16764 3460
rect 16715 3420 16764 3448
rect 16715 3417 16727 3420
rect 16669 3411 16727 3417
rect 16758 3408 16764 3420
rect 16816 3448 16822 3460
rect 17494 3448 17500 3460
rect 16816 3420 17500 3448
rect 16816 3408 16822 3420
rect 17494 3408 17500 3420
rect 17552 3408 17558 3460
rect 19886 3408 19892 3460
rect 19944 3448 19950 3460
rect 20533 3451 20591 3457
rect 20533 3448 20545 3451
rect 19944 3420 20545 3448
rect 19944 3408 19950 3420
rect 20533 3417 20545 3420
rect 20579 3448 20591 3451
rect 20714 3448 20720 3460
rect 20579 3420 20720 3448
rect 20579 3417 20591 3420
rect 20533 3411 20591 3417
rect 20714 3408 20720 3420
rect 20772 3408 20778 3460
rect 11974 3380 11980 3392
rect 11935 3352 11980 3380
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 15105 3383 15163 3389
rect 15105 3349 15117 3383
rect 15151 3380 15163 3383
rect 15286 3380 15292 3392
rect 15151 3352 15292 3380
rect 15151 3349 15163 3352
rect 15105 3343 15163 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 17681 3383 17739 3389
rect 17681 3349 17693 3383
rect 17727 3380 17739 3383
rect 18046 3380 18052 3392
rect 17727 3352 18052 3380
rect 17727 3349 17739 3352
rect 17681 3343 17739 3349
rect 18046 3340 18052 3352
rect 18104 3380 18110 3392
rect 18782 3380 18788 3392
rect 18104 3352 18788 3380
rect 18104 3340 18110 3352
rect 18782 3340 18788 3352
rect 18840 3380 18846 3392
rect 19153 3383 19211 3389
rect 19153 3380 19165 3383
rect 18840 3352 19165 3380
rect 18840 3340 18846 3352
rect 19153 3349 19165 3352
rect 19199 3349 19211 3383
rect 22738 3380 22744 3392
rect 22699 3352 22744 3380
rect 19153 3343 19211 3349
rect 22738 3340 22744 3352
rect 22796 3340 22802 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 10689 3179 10747 3185
rect 10689 3176 10701 3179
rect 9916 3148 10701 3176
rect 9916 3136 9922 3148
rect 10152 2981 10180 3148
rect 10689 3145 10701 3148
rect 10735 3145 10747 3179
rect 11422 3176 11428 3188
rect 11383 3148 11428 3176
rect 10689 3139 10747 3145
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 11882 3176 11888 3188
rect 11843 3148 11888 3176
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 12250 3176 12256 3188
rect 12211 3148 12256 3176
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 13446 3176 13452 3188
rect 13407 3148 13452 3176
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 15654 3136 15660 3188
rect 15712 3176 15718 3188
rect 15933 3179 15991 3185
rect 15933 3176 15945 3179
rect 15712 3148 15945 3176
rect 15712 3136 15718 3148
rect 15933 3145 15945 3148
rect 15979 3176 15991 3179
rect 16298 3176 16304 3188
rect 15979 3148 16304 3176
rect 15979 3145 15991 3148
rect 15933 3139 15991 3145
rect 16298 3136 16304 3148
rect 16356 3136 16362 3188
rect 17494 3176 17500 3188
rect 17455 3148 17500 3176
rect 17494 3136 17500 3148
rect 17552 3136 17558 3188
rect 18325 3179 18383 3185
rect 18325 3145 18337 3179
rect 18371 3176 18383 3179
rect 18966 3176 18972 3188
rect 18371 3148 18972 3176
rect 18371 3145 18383 3148
rect 18325 3139 18383 3145
rect 18966 3136 18972 3148
rect 19024 3136 19030 3188
rect 23477 3179 23535 3185
rect 23477 3145 23489 3179
rect 23523 3176 23535 3179
rect 23566 3176 23572 3188
rect 23523 3148 23572 3176
rect 23523 3145 23535 3148
rect 23477 3139 23535 3145
rect 23566 3136 23572 3148
rect 23624 3136 23630 3188
rect 24118 3136 24124 3188
rect 24176 3176 24182 3188
rect 24397 3179 24455 3185
rect 24397 3176 24409 3179
rect 24176 3148 24409 3176
rect 24176 3136 24182 3148
rect 24397 3145 24409 3148
rect 24443 3145 24455 3179
rect 24397 3139 24455 3145
rect 24857 3179 24915 3185
rect 24857 3145 24869 3179
rect 24903 3176 24915 3179
rect 25038 3176 25044 3188
rect 24903 3148 25044 3176
rect 24903 3145 24915 3148
rect 24857 3139 24915 3145
rect 25038 3136 25044 3148
rect 25096 3136 25102 3188
rect 10318 3108 10324 3120
rect 10279 3080 10324 3108
rect 10318 3068 10324 3080
rect 10376 3068 10382 3120
rect 11149 3111 11207 3117
rect 11149 3077 11161 3111
rect 11195 3108 11207 3111
rect 11514 3108 11520 3120
rect 11195 3080 11520 3108
rect 11195 3077 11207 3080
rect 11149 3071 11207 3077
rect 11514 3068 11520 3080
rect 11572 3068 11578 3120
rect 13464 3040 13492 3136
rect 15013 3111 15071 3117
rect 15013 3077 15025 3111
rect 15059 3108 15071 3111
rect 15286 3108 15292 3120
rect 15059 3080 15292 3108
rect 15059 3077 15071 3080
rect 15013 3071 15071 3077
rect 15286 3068 15292 3080
rect 15344 3108 15350 3120
rect 16114 3108 16120 3120
rect 15344 3080 16120 3108
rect 15344 3068 15350 3080
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 21358 3068 21364 3120
rect 21416 3108 21422 3120
rect 22557 3111 22615 3117
rect 22557 3108 22569 3111
rect 21416 3080 22569 3108
rect 21416 3068 21422 3080
rect 22557 3077 22569 3080
rect 22603 3077 22615 3111
rect 22557 3071 22615 3077
rect 15657 3043 15715 3049
rect 13464 3012 13768 3040
rect 10137 2975 10195 2981
rect 10137 2941 10149 2975
rect 10183 2941 10195 2975
rect 10137 2935 10195 2941
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11882 2972 11888 2984
rect 11287 2944 11888 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11882 2932 11888 2944
rect 11940 2932 11946 2984
rect 12529 2975 12587 2981
rect 12529 2941 12541 2975
rect 12575 2941 12587 2975
rect 12529 2935 12587 2941
rect 12544 2904 12572 2935
rect 12618 2932 12624 2984
rect 12676 2972 12682 2984
rect 13633 2975 13691 2981
rect 13633 2972 13645 2975
rect 12676 2944 13645 2972
rect 12676 2932 12682 2944
rect 13633 2941 13645 2944
rect 13679 2941 13691 2975
rect 13740 2972 13768 3012
rect 15657 3009 15669 3043
rect 15703 3040 15715 3043
rect 16758 3040 16764 3052
rect 15703 3012 16764 3040
rect 15703 3009 15715 3012
rect 15657 3003 15715 3009
rect 16758 3000 16764 3012
rect 16816 3000 16822 3052
rect 18230 3000 18236 3052
rect 18288 3040 18294 3052
rect 18785 3043 18843 3049
rect 18785 3040 18797 3043
rect 18288 3012 18797 3040
rect 18288 3000 18294 3012
rect 18785 3009 18797 3012
rect 18831 3009 18843 3043
rect 18785 3003 18843 3009
rect 18969 3043 19027 3049
rect 18969 3009 18981 3043
rect 19015 3040 19027 3043
rect 19337 3043 19395 3049
rect 19337 3040 19349 3043
rect 19015 3012 19349 3040
rect 19015 3009 19027 3012
rect 18969 3003 19027 3009
rect 19337 3009 19349 3012
rect 19383 3040 19395 3043
rect 19518 3040 19524 3052
rect 19383 3012 19524 3040
rect 19383 3009 19395 3012
rect 19337 3003 19395 3009
rect 13889 2975 13947 2981
rect 13889 2972 13901 2975
rect 13740 2944 13901 2972
rect 13633 2935 13691 2941
rect 13889 2941 13901 2944
rect 13935 2941 13947 2975
rect 13889 2935 13947 2941
rect 16482 2932 16488 2984
rect 16540 2972 16546 2984
rect 16577 2975 16635 2981
rect 16577 2972 16589 2975
rect 16540 2944 16589 2972
rect 16540 2932 16546 2944
rect 16577 2941 16589 2944
rect 16623 2941 16635 2975
rect 18800 2972 18828 3003
rect 19518 3000 19524 3012
rect 19576 3040 19582 3052
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 19576 3012 19717 3040
rect 19576 3000 19582 3012
rect 19705 3009 19717 3012
rect 19751 3040 19763 3043
rect 23842 3040 23848 3052
rect 19751 3012 20024 3040
rect 23803 3012 23848 3040
rect 19751 3009 19763 3012
rect 19705 3003 19763 3009
rect 19242 2972 19248 2984
rect 18800 2944 19248 2972
rect 16577 2935 16635 2941
rect 19242 2932 19248 2944
rect 19300 2932 19306 2984
rect 19886 2972 19892 2984
rect 19847 2944 19892 2972
rect 19886 2932 19892 2944
rect 19944 2932 19950 2984
rect 19996 2972 20024 3012
rect 23842 3000 23848 3012
rect 23900 3000 23906 3052
rect 20145 2975 20203 2981
rect 20145 2972 20157 2975
rect 19996 2944 20157 2972
rect 20145 2941 20157 2944
rect 20191 2941 20203 2975
rect 20145 2935 20203 2941
rect 20714 2932 20720 2984
rect 20772 2972 20778 2984
rect 22189 2975 22247 2981
rect 22189 2972 22201 2975
rect 20772 2944 22201 2972
rect 20772 2932 20778 2944
rect 22189 2941 22201 2944
rect 22235 2941 22247 2975
rect 22189 2935 22247 2941
rect 22373 2975 22431 2981
rect 22373 2941 22385 2975
rect 22419 2972 22431 2975
rect 22922 2972 22928 2984
rect 22419 2944 22928 2972
rect 22419 2941 22431 2944
rect 22373 2935 22431 2941
rect 22922 2932 22928 2944
rect 22980 2932 22986 2984
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23624 2944 23673 2972
rect 23624 2932 23630 2944
rect 23661 2941 23673 2944
rect 23707 2941 23719 2975
rect 23661 2935 23719 2941
rect 24949 2975 25007 2981
rect 24949 2941 24961 2975
rect 24995 2972 25007 2975
rect 25130 2972 25136 2984
rect 24995 2944 25136 2972
rect 24995 2941 25007 2944
rect 24949 2935 25007 2941
rect 25130 2932 25136 2944
rect 25188 2972 25194 2984
rect 25685 2975 25743 2981
rect 25685 2972 25697 2975
rect 25188 2944 25697 2972
rect 25188 2932 25194 2944
rect 25685 2941 25697 2944
rect 25731 2941 25743 2975
rect 25685 2935 25743 2941
rect 13170 2904 13176 2916
rect 12544 2876 13176 2904
rect 13170 2864 13176 2876
rect 13228 2864 13234 2916
rect 16666 2904 16672 2916
rect 16132 2876 16672 2904
rect 9950 2836 9956 2848
rect 9911 2808 9956 2836
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 12710 2836 12716 2848
rect 12671 2808 12716 2836
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 16132 2845 16160 2876
rect 16666 2864 16672 2876
rect 16724 2864 16730 2916
rect 17865 2907 17923 2913
rect 17865 2873 17877 2907
rect 17911 2904 17923 2907
rect 18693 2907 18751 2913
rect 18693 2904 18705 2907
rect 17911 2876 18705 2904
rect 17911 2873 17923 2876
rect 17865 2867 17923 2873
rect 18693 2873 18705 2876
rect 18739 2904 18751 2907
rect 19426 2904 19432 2916
rect 18739 2876 19432 2904
rect 18739 2873 18751 2876
rect 18693 2867 18751 2873
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 25222 2904 25228 2916
rect 25183 2876 25228 2904
rect 25222 2864 25228 2876
rect 25280 2864 25286 2916
rect 16117 2839 16175 2845
rect 16117 2805 16129 2839
rect 16163 2805 16175 2839
rect 16117 2799 16175 2805
rect 16298 2796 16304 2848
rect 16356 2836 16362 2848
rect 16485 2839 16543 2845
rect 16485 2836 16497 2839
rect 16356 2808 16497 2836
rect 16356 2796 16362 2808
rect 16485 2805 16497 2808
rect 16531 2805 16543 2839
rect 16485 2799 16543 2805
rect 21269 2839 21327 2845
rect 21269 2805 21281 2839
rect 21315 2836 21327 2839
rect 21910 2836 21916 2848
rect 21315 2808 21916 2836
rect 21315 2805 21327 2808
rect 21269 2799 21327 2805
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 10965 2635 11023 2641
rect 10965 2601 10977 2635
rect 11011 2632 11023 2635
rect 11238 2632 11244 2644
rect 11011 2604 11244 2632
rect 11011 2601 11023 2604
rect 10965 2595 11023 2601
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 10321 2499 10379 2505
rect 8619 2468 9260 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 9232 2372 9260 2468
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 10980 2496 11008 2595
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 12066 2632 12072 2644
rect 12027 2604 12072 2632
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 12618 2632 12624 2644
rect 12483 2604 12624 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 14001 2635 14059 2641
rect 14001 2601 14013 2635
rect 14047 2632 14059 2635
rect 14642 2632 14648 2644
rect 14047 2604 14648 2632
rect 14047 2601 14059 2604
rect 14001 2595 14059 2601
rect 10367 2468 11008 2496
rect 11425 2499 11483 2505
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 12084 2496 12112 2592
rect 12802 2496 12808 2508
rect 11471 2468 12112 2496
rect 12715 2468 12808 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 12802 2456 12808 2468
rect 12860 2496 12866 2508
rect 14108 2505 14136 2604
rect 14642 2592 14648 2604
rect 14700 2592 14706 2644
rect 18046 2632 18052 2644
rect 18007 2604 18052 2632
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 19797 2635 19855 2641
rect 19797 2632 19809 2635
rect 19576 2604 19809 2632
rect 19576 2592 19582 2604
rect 19797 2601 19809 2604
rect 19843 2601 19855 2635
rect 20714 2632 20720 2644
rect 20675 2604 20720 2632
rect 19797 2595 19855 2601
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 22002 2632 22008 2644
rect 21963 2604 22008 2632
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 23477 2635 23535 2641
rect 23477 2601 23489 2635
rect 23523 2632 23535 2635
rect 24489 2635 24547 2641
rect 24489 2632 24501 2635
rect 23523 2604 24501 2632
rect 23523 2601 23535 2604
rect 23477 2595 23535 2601
rect 24489 2601 24501 2604
rect 24535 2632 24547 2635
rect 24578 2632 24584 2644
rect 24535 2604 24584 2632
rect 24535 2601 24547 2604
rect 24489 2595 24547 2601
rect 24578 2592 24584 2604
rect 24636 2592 24642 2644
rect 24854 2592 24860 2644
rect 24912 2632 24918 2644
rect 25593 2635 25651 2641
rect 25593 2632 25605 2635
rect 24912 2604 25605 2632
rect 24912 2592 24918 2604
rect 25593 2601 25605 2604
rect 25639 2601 25651 2635
rect 25593 2595 25651 2601
rect 18064 2564 18092 2592
rect 18662 2567 18720 2573
rect 18662 2564 18674 2567
rect 18064 2536 18674 2564
rect 18662 2533 18674 2536
rect 18708 2533 18720 2567
rect 18662 2527 18720 2533
rect 19242 2524 19248 2576
rect 19300 2564 19306 2576
rect 20349 2567 20407 2573
rect 20349 2564 20361 2567
rect 19300 2536 20361 2564
rect 19300 2524 19306 2536
rect 20349 2533 20361 2536
rect 20395 2533 20407 2567
rect 20349 2527 20407 2533
rect 21545 2567 21603 2573
rect 21545 2533 21557 2567
rect 21591 2564 21603 2567
rect 21591 2536 22692 2564
rect 21591 2533 21603 2536
rect 21545 2527 21603 2533
rect 13541 2499 13599 2505
rect 13541 2496 13553 2499
rect 12860 2468 13553 2496
rect 12860 2456 12866 2468
rect 13541 2465 13553 2468
rect 13587 2465 13599 2499
rect 13541 2459 13599 2465
rect 14093 2499 14151 2505
rect 14093 2465 14105 2499
rect 14139 2465 14151 2499
rect 14093 2459 14151 2465
rect 15378 2456 15384 2508
rect 15436 2496 15442 2508
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 15436 2468 15853 2496
rect 15436 2456 15442 2468
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 15841 2459 15899 2465
rect 15933 2499 15991 2505
rect 15933 2465 15945 2499
rect 15979 2496 15991 2499
rect 16390 2496 16396 2508
rect 15979 2468 16396 2496
rect 15979 2465 15991 2468
rect 15933 2459 15991 2465
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12492 2400 13001 2428
rect 12492 2388 12498 2400
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 14274 2428 14280 2440
rect 14235 2400 14280 2428
rect 12989 2391 13047 2397
rect 14274 2388 14280 2400
rect 14332 2388 14338 2440
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15948 2428 15976 2459
rect 16390 2456 16396 2468
rect 16448 2456 16454 2508
rect 17129 2499 17187 2505
rect 17129 2465 17141 2499
rect 17175 2496 17187 2499
rect 17770 2496 17776 2508
rect 17175 2468 17776 2496
rect 17175 2465 17187 2468
rect 17129 2459 17187 2465
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 18414 2496 18420 2508
rect 18375 2468 18420 2496
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 21821 2499 21879 2505
rect 21821 2496 21833 2499
rect 20220 2468 21833 2496
rect 20220 2456 20226 2468
rect 21821 2465 21833 2468
rect 21867 2496 21879 2499
rect 22373 2499 22431 2505
rect 22373 2496 22385 2499
rect 21867 2468 22385 2496
rect 21867 2465 21879 2468
rect 21821 2459 21879 2465
rect 22373 2465 22385 2468
rect 22419 2465 22431 2499
rect 22373 2459 22431 2465
rect 16114 2428 16120 2440
rect 14967 2400 15976 2428
rect 16075 2400 16120 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 16114 2388 16120 2400
rect 16172 2428 16178 2440
rect 22664 2437 22692 2536
rect 23750 2456 23756 2508
rect 23808 2496 23814 2508
rect 24397 2499 24455 2505
rect 24397 2496 24409 2499
rect 23808 2468 24409 2496
rect 23808 2456 23814 2468
rect 24397 2465 24409 2468
rect 24443 2465 24455 2499
rect 24397 2459 24455 2465
rect 16485 2431 16543 2437
rect 16485 2428 16497 2431
rect 16172 2400 16497 2428
rect 16172 2388 16178 2400
rect 16485 2397 16497 2400
rect 16531 2397 16543 2431
rect 16485 2391 16543 2397
rect 22465 2431 22523 2437
rect 22465 2397 22477 2431
rect 22511 2397 22523 2431
rect 22465 2391 22523 2397
rect 22649 2431 22707 2437
rect 22649 2397 22661 2431
rect 22695 2428 22707 2431
rect 22738 2428 22744 2440
rect 22695 2400 22744 2428
rect 22695 2397 22707 2400
rect 22649 2391 22707 2397
rect 9214 2360 9220 2372
rect 9175 2332 9220 2360
rect 9214 2320 9220 2332
rect 9272 2320 9278 2372
rect 15473 2363 15531 2369
rect 15473 2329 15485 2363
rect 15519 2360 15531 2363
rect 16853 2363 16911 2369
rect 16853 2360 16865 2363
rect 15519 2332 16865 2360
rect 15519 2329 15531 2332
rect 15473 2323 15531 2329
rect 16500 2304 16528 2332
rect 16853 2329 16865 2332
rect 16899 2329 16911 2363
rect 22480 2360 22508 2391
rect 22738 2388 22744 2400
rect 22796 2388 22802 2440
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 24544 2400 24593 2428
rect 24544 2388 24550 2400
rect 24581 2397 24593 2400
rect 24627 2428 24639 2431
rect 25041 2431 25099 2437
rect 25041 2428 25053 2431
rect 24627 2400 25053 2428
rect 24627 2397 24639 2400
rect 24581 2391 24639 2397
rect 25041 2397 25053 2400
rect 25087 2397 25099 2431
rect 25041 2391 25099 2397
rect 23109 2363 23167 2369
rect 23109 2360 23121 2363
rect 22480 2332 23121 2360
rect 16853 2323 16911 2329
rect 23109 2329 23121 2332
rect 23155 2360 23167 2363
rect 24029 2363 24087 2369
rect 24029 2360 24041 2363
rect 23155 2332 24041 2360
rect 23155 2329 23167 2332
rect 23109 2323 23167 2329
rect 24029 2329 24041 2332
rect 24075 2329 24087 2363
rect 24029 2323 24087 2329
rect 8754 2292 8760 2304
rect 8715 2264 8760 2292
rect 8754 2252 8760 2264
rect 8812 2252 8818 2304
rect 10505 2295 10563 2301
rect 10505 2261 10517 2295
rect 10551 2292 10563 2295
rect 10962 2292 10968 2304
rect 10551 2264 10968 2292
rect 10551 2261 10563 2264
rect 10505 2255 10563 2261
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 15289 2295 15347 2301
rect 15289 2261 15301 2295
rect 15335 2292 15347 2295
rect 15378 2292 15384 2304
rect 15335 2264 15384 2292
rect 15335 2261 15347 2264
rect 15289 2255 15347 2261
rect 15378 2252 15384 2264
rect 15436 2252 15442 2304
rect 16482 2252 16488 2304
rect 16540 2252 16546 2304
rect 17313 2295 17371 2301
rect 17313 2261 17325 2295
rect 17359 2292 17371 2295
rect 17586 2292 17592 2304
rect 17359 2264 17592 2292
rect 17359 2261 17371 2264
rect 17313 2255 17371 2261
rect 17586 2252 17592 2264
rect 17644 2252 17650 2304
rect 23750 2292 23756 2304
rect 23711 2264 23756 2292
rect 23750 2252 23756 2264
rect 23808 2252 23814 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 21266 552 21272 604
rect 21324 592 21330 604
rect 23474 592 23480 604
rect 21324 564 23480 592
rect 21324 552 21330 564
rect 23474 552 23480 564
rect 23532 552 23538 604
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 17316 25440 17368 25492
rect 22744 25440 22796 25492
rect 24584 25440 24636 25492
rect 24768 25483 24820 25492
rect 24768 25449 24777 25483
rect 24777 25449 24811 25483
rect 24811 25449 24820 25483
rect 24768 25440 24820 25449
rect 24124 25372 24176 25424
rect 16304 25304 16356 25356
rect 18972 25304 19024 25356
rect 20168 25304 20220 25356
rect 22376 25304 22428 25356
rect 22560 25304 22612 25356
rect 23940 25304 23992 25356
rect 26884 25168 26936 25220
rect 19432 25143 19484 25152
rect 19432 25109 19441 25143
rect 19441 25109 19475 25143
rect 19475 25109 19484 25143
rect 19432 25100 19484 25109
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 24768 24896 24820 24948
rect 22560 24828 22612 24880
rect 17040 24760 17092 24812
rect 16856 24735 16908 24744
rect 16856 24701 16865 24735
rect 16865 24701 16899 24735
rect 16899 24701 16908 24735
rect 16856 24692 16908 24701
rect 14372 24599 14424 24608
rect 14372 24565 14381 24599
rect 14381 24565 14415 24599
rect 14415 24565 14424 24599
rect 14372 24556 14424 24565
rect 14556 24556 14608 24608
rect 16488 24624 16540 24676
rect 19248 24692 19300 24744
rect 20260 24735 20312 24744
rect 20260 24701 20269 24735
rect 20269 24701 20303 24735
rect 20303 24701 20312 24735
rect 20260 24692 20312 24701
rect 21916 24692 21968 24744
rect 22468 24735 22520 24744
rect 22468 24701 22477 24735
rect 22477 24701 22511 24735
rect 22511 24701 22520 24735
rect 22468 24692 22520 24701
rect 23848 24692 23900 24744
rect 16304 24556 16356 24608
rect 17776 24599 17828 24608
rect 17776 24565 17785 24599
rect 17785 24565 17819 24599
rect 17819 24565 17828 24599
rect 17776 24556 17828 24565
rect 17960 24556 18012 24608
rect 18972 24599 19024 24608
rect 18972 24565 18981 24599
rect 18981 24565 19015 24599
rect 19015 24565 19024 24599
rect 18972 24556 19024 24565
rect 20076 24624 20128 24676
rect 20168 24556 20220 24608
rect 20628 24556 20680 24608
rect 22008 24624 22060 24676
rect 21916 24599 21968 24608
rect 21916 24565 21925 24599
rect 21925 24565 21959 24599
rect 21959 24565 21968 24599
rect 21916 24556 21968 24565
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 23296 24556 23348 24608
rect 23940 24556 23992 24608
rect 24768 24599 24820 24608
rect 24768 24565 24777 24599
rect 24777 24565 24811 24599
rect 24811 24565 24820 24599
rect 24768 24556 24820 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 13728 24352 13780 24404
rect 15108 24352 15160 24404
rect 17960 24395 18012 24404
rect 17960 24361 17969 24395
rect 17969 24361 18003 24395
rect 18003 24361 18012 24395
rect 17960 24352 18012 24361
rect 18696 24352 18748 24404
rect 21364 24352 21416 24404
rect 23112 24352 23164 24404
rect 23664 24395 23716 24404
rect 23664 24361 23673 24395
rect 23673 24361 23707 24395
rect 23707 24361 23716 24395
rect 23664 24352 23716 24361
rect 13912 24284 13964 24336
rect 16396 24284 16448 24336
rect 14096 24259 14148 24268
rect 14096 24225 14105 24259
rect 14105 24225 14139 24259
rect 14139 24225 14148 24259
rect 14096 24216 14148 24225
rect 14188 24216 14240 24268
rect 15752 24259 15804 24268
rect 15752 24225 15761 24259
rect 15761 24225 15795 24259
rect 15795 24225 15804 24259
rect 15752 24216 15804 24225
rect 17684 24216 17736 24268
rect 20076 24284 20128 24336
rect 19156 24259 19208 24268
rect 19156 24225 19165 24259
rect 19165 24225 19199 24259
rect 19199 24225 19208 24259
rect 19156 24216 19208 24225
rect 21732 24216 21784 24268
rect 23020 24216 23072 24268
rect 23480 24259 23532 24268
rect 23480 24225 23489 24259
rect 23489 24225 23523 24259
rect 23523 24225 23532 24259
rect 23480 24216 23532 24225
rect 24032 24216 24084 24268
rect 16028 24148 16080 24200
rect 18328 24080 18380 24132
rect 16488 24012 16540 24064
rect 16672 24055 16724 24064
rect 16672 24021 16681 24055
rect 16681 24021 16715 24055
rect 16715 24021 16724 24055
rect 16672 24012 16724 24021
rect 17408 24055 17460 24064
rect 17408 24021 17417 24055
rect 17417 24021 17451 24055
rect 17451 24021 17460 24055
rect 17408 24012 17460 24021
rect 17592 24055 17644 24064
rect 17592 24021 17601 24055
rect 17601 24021 17635 24055
rect 17635 24021 17644 24055
rect 17592 24012 17644 24021
rect 24676 24012 24728 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 12808 23851 12860 23860
rect 12808 23817 12817 23851
rect 12817 23817 12851 23851
rect 12851 23817 12860 23851
rect 12808 23808 12860 23817
rect 15752 23808 15804 23860
rect 16396 23851 16448 23860
rect 16396 23817 16405 23851
rect 16405 23817 16439 23851
rect 16439 23817 16448 23851
rect 16396 23808 16448 23817
rect 17132 23808 17184 23860
rect 17684 23851 17736 23860
rect 17684 23817 17693 23851
rect 17693 23817 17727 23851
rect 17727 23817 17736 23851
rect 17684 23808 17736 23817
rect 19524 23808 19576 23860
rect 23204 23808 23256 23860
rect 16856 23715 16908 23724
rect 16856 23681 16865 23715
rect 16865 23681 16899 23715
rect 16899 23681 16908 23715
rect 16856 23672 16908 23681
rect 13452 23536 13504 23588
rect 16672 23604 16724 23656
rect 17500 23604 17552 23656
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 18328 23647 18380 23656
rect 18328 23613 18362 23647
rect 18362 23613 18380 23647
rect 18328 23604 18380 23613
rect 20076 23604 20128 23656
rect 19156 23536 19208 23588
rect 24216 23604 24268 23656
rect 23572 23536 23624 23588
rect 13544 23511 13596 23520
rect 13544 23477 13553 23511
rect 13553 23477 13587 23511
rect 13587 23477 13596 23511
rect 13544 23468 13596 23477
rect 14004 23511 14056 23520
rect 14004 23477 14013 23511
rect 14013 23477 14047 23511
rect 14047 23477 14056 23511
rect 14004 23468 14056 23477
rect 15384 23468 15436 23520
rect 19340 23468 19392 23520
rect 21732 23468 21784 23520
rect 23020 23511 23072 23520
rect 23020 23477 23029 23511
rect 23029 23477 23063 23511
rect 23063 23477 23072 23511
rect 23020 23468 23072 23477
rect 23480 23468 23532 23520
rect 24032 23468 24084 23520
rect 24768 23511 24820 23520
rect 24768 23477 24777 23511
rect 24777 23477 24811 23511
rect 24811 23477 24820 23511
rect 24768 23468 24820 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 12624 23264 12676 23316
rect 13544 23264 13596 23316
rect 14648 23307 14700 23316
rect 14648 23273 14657 23307
rect 14657 23273 14691 23307
rect 14691 23273 14700 23307
rect 14648 23264 14700 23273
rect 17868 23264 17920 23316
rect 18052 23264 18104 23316
rect 19064 23264 19116 23316
rect 17592 23196 17644 23248
rect 23480 23196 23532 23248
rect 23572 23196 23624 23248
rect 10692 23171 10744 23180
rect 10692 23137 10726 23171
rect 10726 23137 10744 23171
rect 13268 23171 13320 23180
rect 10692 23128 10744 23137
rect 13268 23137 13277 23171
rect 13277 23137 13311 23171
rect 13311 23137 13320 23171
rect 13268 23128 13320 23137
rect 15384 23128 15436 23180
rect 16028 23128 16080 23180
rect 10048 22924 10100 22976
rect 13544 23103 13596 23112
rect 13544 23069 13553 23103
rect 13553 23069 13587 23103
rect 13587 23069 13596 23103
rect 13544 23060 13596 23069
rect 14648 23060 14700 23112
rect 20260 23128 20312 23180
rect 20812 23128 20864 23180
rect 22928 23128 22980 23180
rect 23756 23171 23808 23180
rect 23756 23137 23765 23171
rect 23765 23137 23799 23171
rect 23799 23137 23808 23171
rect 23756 23128 23808 23137
rect 25044 23171 25096 23180
rect 25044 23137 25053 23171
rect 25053 23137 25087 23171
rect 25087 23137 25096 23171
rect 25044 23128 25096 23137
rect 18420 23103 18472 23112
rect 18420 23069 18429 23103
rect 18429 23069 18463 23103
rect 18463 23069 18472 23103
rect 18420 23060 18472 23069
rect 19340 23060 19392 23112
rect 19800 23103 19852 23112
rect 19800 23069 19809 23103
rect 19809 23069 19843 23103
rect 19843 23069 19852 23103
rect 19800 23060 19852 23069
rect 20996 23060 21048 23112
rect 21456 23103 21508 23112
rect 21456 23069 21465 23103
rect 21465 23069 21499 23103
rect 21499 23069 21508 23103
rect 21456 23060 21508 23069
rect 22100 23060 22152 23112
rect 11796 22967 11848 22976
rect 11796 22933 11805 22967
rect 11805 22933 11839 22967
rect 11839 22933 11848 22967
rect 11796 22924 11848 22933
rect 12716 22967 12768 22976
rect 12716 22933 12725 22967
rect 12725 22933 12759 22967
rect 12759 22933 12768 22967
rect 12716 22924 12768 22933
rect 12900 22967 12952 22976
rect 12900 22933 12909 22967
rect 12909 22933 12943 22967
rect 12943 22933 12952 22967
rect 12900 22924 12952 22933
rect 14096 22967 14148 22976
rect 14096 22933 14105 22967
rect 14105 22933 14139 22967
rect 14139 22933 14148 22967
rect 14096 22924 14148 22933
rect 17408 22924 17460 22976
rect 20904 22967 20956 22976
rect 20904 22933 20913 22967
rect 20913 22933 20947 22967
rect 20947 22933 20956 22967
rect 20904 22924 20956 22933
rect 21916 22967 21968 22976
rect 21916 22933 21925 22967
rect 21925 22933 21959 22967
rect 21959 22933 21968 22967
rect 21916 22924 21968 22933
rect 25320 22924 25372 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 10600 22763 10652 22772
rect 10600 22729 10609 22763
rect 10609 22729 10643 22763
rect 10643 22729 10652 22763
rect 10600 22720 10652 22729
rect 10784 22763 10836 22772
rect 10784 22729 10793 22763
rect 10793 22729 10827 22763
rect 10827 22729 10836 22763
rect 10784 22720 10836 22729
rect 11796 22720 11848 22772
rect 12716 22720 12768 22772
rect 16580 22720 16632 22772
rect 17592 22720 17644 22772
rect 17868 22763 17920 22772
rect 17868 22729 17877 22763
rect 17877 22729 17911 22763
rect 17911 22729 17920 22763
rect 17868 22720 17920 22729
rect 18420 22720 18472 22772
rect 20996 22763 21048 22772
rect 20996 22729 21005 22763
rect 21005 22729 21039 22763
rect 21039 22729 21048 22763
rect 20996 22720 21048 22729
rect 23572 22720 23624 22772
rect 23756 22720 23808 22772
rect 25044 22720 25096 22772
rect 25504 22720 25556 22772
rect 11152 22559 11204 22568
rect 11152 22525 11161 22559
rect 11161 22525 11195 22559
rect 11195 22525 11204 22559
rect 11152 22516 11204 22525
rect 14648 22584 14700 22636
rect 11888 22516 11940 22568
rect 9864 22448 9916 22500
rect 12716 22559 12768 22568
rect 12716 22525 12750 22559
rect 12750 22525 12768 22559
rect 19064 22559 19116 22568
rect 12716 22516 12768 22525
rect 19064 22525 19073 22559
rect 19073 22525 19107 22559
rect 19107 22525 19116 22559
rect 19064 22516 19116 22525
rect 19340 22559 19392 22568
rect 19340 22525 19374 22559
rect 19374 22525 19392 22559
rect 19340 22516 19392 22525
rect 19892 22516 19944 22568
rect 20168 22516 20220 22568
rect 22100 22627 22152 22636
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 23940 22627 23992 22636
rect 22100 22584 22152 22593
rect 23940 22593 23949 22627
rect 23949 22593 23983 22627
rect 23983 22593 23992 22627
rect 23940 22584 23992 22593
rect 21088 22516 21140 22568
rect 21916 22559 21968 22568
rect 21916 22525 21925 22559
rect 21925 22525 21959 22559
rect 21959 22525 21968 22559
rect 21916 22516 21968 22525
rect 12624 22448 12676 22500
rect 10140 22380 10192 22432
rect 13544 22380 13596 22432
rect 20812 22448 20864 22500
rect 23664 22559 23716 22568
rect 23664 22525 23673 22559
rect 23673 22525 23707 22559
rect 23707 22525 23716 22559
rect 23664 22516 23716 22525
rect 24952 22559 25004 22568
rect 24952 22525 24961 22559
rect 24961 22525 24995 22559
rect 24995 22525 25004 22559
rect 24952 22516 25004 22525
rect 14832 22380 14884 22432
rect 18052 22423 18104 22432
rect 18052 22389 18061 22423
rect 18061 22389 18095 22423
rect 18095 22389 18104 22423
rect 18052 22380 18104 22389
rect 20720 22380 20772 22432
rect 21548 22423 21600 22432
rect 21548 22389 21557 22423
rect 21557 22389 21591 22423
rect 21591 22389 21600 22423
rect 21548 22380 21600 22389
rect 22928 22423 22980 22432
rect 22928 22389 22937 22423
rect 22937 22389 22971 22423
rect 22971 22389 22980 22423
rect 22928 22380 22980 22389
rect 24676 22380 24728 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 9864 22176 9916 22228
rect 10692 22176 10744 22228
rect 12256 22219 12308 22228
rect 12256 22185 12265 22219
rect 12265 22185 12299 22219
rect 12299 22185 12308 22219
rect 12256 22176 12308 22185
rect 12992 22219 13044 22228
rect 12992 22185 13001 22219
rect 13001 22185 13035 22219
rect 13035 22185 13044 22219
rect 12992 22176 13044 22185
rect 13268 22176 13320 22228
rect 16028 22219 16080 22228
rect 16028 22185 16037 22219
rect 16037 22185 16071 22219
rect 16071 22185 16080 22219
rect 16028 22176 16080 22185
rect 16580 22176 16632 22228
rect 19524 22176 19576 22228
rect 20904 22176 20956 22228
rect 12900 22108 12952 22160
rect 20260 22151 20312 22160
rect 20260 22117 20269 22151
rect 20269 22117 20303 22151
rect 20303 22117 20312 22151
rect 20260 22108 20312 22117
rect 9772 22040 9824 22092
rect 10232 22040 10284 22092
rect 13268 22040 13320 22092
rect 14004 22040 14056 22092
rect 14832 22040 14884 22092
rect 8208 21879 8260 21888
rect 8208 21845 8217 21879
rect 8217 21845 8251 21879
rect 8251 21845 8260 21879
rect 17316 22040 17368 22092
rect 19708 22083 19760 22092
rect 19708 22049 19717 22083
rect 19717 22049 19751 22083
rect 19751 22049 19760 22083
rect 21548 22108 21600 22160
rect 19708 22040 19760 22049
rect 20720 22040 20772 22092
rect 21456 22040 21508 22092
rect 23756 22083 23808 22092
rect 23756 22049 23765 22083
rect 23765 22049 23799 22083
rect 23799 22049 23808 22083
rect 23756 22040 23808 22049
rect 24032 22083 24084 22092
rect 24032 22049 24041 22083
rect 24041 22049 24075 22083
rect 24075 22049 24084 22083
rect 24032 22040 24084 22049
rect 25044 22083 25096 22092
rect 25044 22049 25053 22083
rect 25053 22049 25087 22083
rect 25087 22049 25096 22083
rect 25044 22040 25096 22049
rect 15568 22015 15620 22024
rect 15568 21981 15577 22015
rect 15577 21981 15611 22015
rect 15611 21981 15620 22015
rect 15568 21972 15620 21981
rect 17408 22015 17460 22024
rect 17408 21981 17417 22015
rect 17417 21981 17451 22015
rect 17451 21981 17460 22015
rect 17408 21972 17460 21981
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 19892 21972 19944 21981
rect 20076 21972 20128 22024
rect 20904 22015 20956 22024
rect 20904 21981 20913 22015
rect 20913 21981 20947 22015
rect 20947 21981 20956 22015
rect 20904 21972 20956 21981
rect 15476 21904 15528 21956
rect 17868 21904 17920 21956
rect 18512 21904 18564 21956
rect 8208 21836 8260 21845
rect 10048 21836 10100 21888
rect 14464 21879 14516 21888
rect 14464 21845 14473 21879
rect 14473 21845 14507 21879
rect 14507 21845 14516 21879
rect 14464 21836 14516 21845
rect 14648 21836 14700 21888
rect 14740 21836 14792 21888
rect 16948 21836 17000 21888
rect 18144 21879 18196 21888
rect 18144 21845 18153 21879
rect 18153 21845 18187 21879
rect 18187 21845 18196 21879
rect 18144 21836 18196 21845
rect 19064 21879 19116 21888
rect 19064 21845 19073 21879
rect 19073 21845 19107 21879
rect 19107 21845 19116 21879
rect 19064 21836 19116 21845
rect 19248 21879 19300 21888
rect 19248 21845 19257 21879
rect 19257 21845 19291 21879
rect 19291 21845 19300 21879
rect 19248 21836 19300 21845
rect 20076 21836 20128 21888
rect 20720 21836 20772 21888
rect 22284 21879 22336 21888
rect 22284 21845 22293 21879
rect 22293 21845 22327 21879
rect 22327 21845 22336 21879
rect 22284 21836 22336 21845
rect 24860 21836 24912 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 12716 21675 12768 21684
rect 12716 21641 12725 21675
rect 12725 21641 12759 21675
rect 12759 21641 12768 21675
rect 12716 21632 12768 21641
rect 13268 21675 13320 21684
rect 13268 21641 13277 21675
rect 13277 21641 13311 21675
rect 13311 21641 13320 21675
rect 13268 21632 13320 21641
rect 14004 21632 14056 21684
rect 17408 21632 17460 21684
rect 19708 21675 19760 21684
rect 19708 21641 19717 21675
rect 19717 21641 19751 21675
rect 19751 21641 19760 21675
rect 19708 21632 19760 21641
rect 20076 21675 20128 21684
rect 20076 21641 20085 21675
rect 20085 21641 20119 21675
rect 20119 21641 20128 21675
rect 20076 21632 20128 21641
rect 20904 21632 20956 21684
rect 21272 21632 21324 21684
rect 25044 21675 25096 21684
rect 25044 21641 25053 21675
rect 25053 21641 25087 21675
rect 25087 21641 25096 21675
rect 25044 21632 25096 21641
rect 11152 21539 11204 21548
rect 11152 21505 11161 21539
rect 11161 21505 11195 21539
rect 11195 21505 11204 21539
rect 11152 21496 11204 21505
rect 7656 21428 7708 21480
rect 8208 21471 8260 21480
rect 8208 21437 8217 21471
rect 8217 21437 8251 21471
rect 8251 21437 8260 21471
rect 8208 21428 8260 21437
rect 10140 21428 10192 21480
rect 13084 21496 13136 21548
rect 13268 21496 13320 21548
rect 13544 21496 13596 21548
rect 16948 21539 17000 21548
rect 12716 21428 12768 21480
rect 14740 21428 14792 21480
rect 16948 21505 16957 21539
rect 16957 21505 16991 21539
rect 16991 21505 17000 21539
rect 16948 21496 17000 21505
rect 18144 21496 18196 21548
rect 19156 21496 19208 21548
rect 19892 21496 19944 21548
rect 24216 21539 24268 21548
rect 16396 21428 16448 21480
rect 18052 21428 18104 21480
rect 19064 21428 19116 21480
rect 20536 21471 20588 21480
rect 20536 21437 20545 21471
rect 20545 21437 20579 21471
rect 20579 21437 20588 21471
rect 20536 21428 20588 21437
rect 24216 21505 24225 21539
rect 24225 21505 24259 21539
rect 24259 21505 24268 21539
rect 24216 21496 24268 21505
rect 25504 21539 25556 21548
rect 25504 21505 25513 21539
rect 25513 21505 25547 21539
rect 25547 21505 25556 21539
rect 25504 21496 25556 21505
rect 22284 21428 22336 21480
rect 23940 21471 23992 21480
rect 23940 21437 23949 21471
rect 23949 21437 23983 21471
rect 23983 21437 23992 21471
rect 23940 21428 23992 21437
rect 25228 21471 25280 21480
rect 25228 21437 25237 21471
rect 25237 21437 25271 21471
rect 25271 21437 25280 21471
rect 25228 21428 25280 21437
rect 8484 21403 8536 21412
rect 8484 21369 8518 21403
rect 8518 21369 8536 21403
rect 8484 21360 8536 21369
rect 12808 21360 12860 21412
rect 12992 21360 13044 21412
rect 14648 21403 14700 21412
rect 14648 21369 14657 21403
rect 14657 21369 14691 21403
rect 14691 21369 14700 21403
rect 14648 21360 14700 21369
rect 17224 21360 17276 21412
rect 18512 21403 18564 21412
rect 18512 21369 18521 21403
rect 18521 21369 18555 21403
rect 18555 21369 18564 21403
rect 18512 21360 18564 21369
rect 10140 21292 10192 21344
rect 10692 21335 10744 21344
rect 10692 21301 10701 21335
rect 10701 21301 10735 21335
rect 10735 21301 10744 21335
rect 10692 21292 10744 21301
rect 11060 21335 11112 21344
rect 11060 21301 11069 21335
rect 11069 21301 11103 21335
rect 11103 21301 11112 21335
rect 11060 21292 11112 21301
rect 12624 21292 12676 21344
rect 14832 21335 14884 21344
rect 14832 21301 14841 21335
rect 14841 21301 14875 21335
rect 14875 21301 14884 21335
rect 14832 21292 14884 21301
rect 16488 21292 16540 21344
rect 16764 21335 16816 21344
rect 16764 21301 16773 21335
rect 16773 21301 16807 21335
rect 16807 21301 16816 21335
rect 16764 21292 16816 21301
rect 16856 21335 16908 21344
rect 16856 21301 16865 21335
rect 16865 21301 16899 21335
rect 16899 21301 16908 21335
rect 16856 21292 16908 21301
rect 17316 21292 17368 21344
rect 18420 21292 18472 21344
rect 21916 21335 21968 21344
rect 21916 21301 21925 21335
rect 21925 21301 21959 21335
rect 21959 21301 21968 21335
rect 21916 21292 21968 21301
rect 23756 21292 23808 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 8208 21131 8260 21140
rect 8208 21097 8217 21131
rect 8217 21097 8251 21131
rect 8251 21097 8260 21131
rect 8208 21088 8260 21097
rect 9772 21088 9824 21140
rect 11060 21088 11112 21140
rect 12900 21131 12952 21140
rect 12900 21097 12909 21131
rect 12909 21097 12943 21131
rect 12943 21097 12952 21131
rect 12900 21088 12952 21097
rect 12992 21088 13044 21140
rect 13452 21088 13504 21140
rect 13544 21088 13596 21140
rect 14832 21088 14884 21140
rect 16856 21088 16908 21140
rect 16948 21088 17000 21140
rect 17408 21088 17460 21140
rect 18052 21131 18104 21140
rect 18052 21097 18061 21131
rect 18061 21097 18095 21131
rect 18095 21097 18104 21131
rect 18052 21088 18104 21097
rect 18144 21088 18196 21140
rect 19064 21088 19116 21140
rect 19524 21088 19576 21140
rect 20536 21088 20588 21140
rect 22652 21131 22704 21140
rect 22652 21097 22661 21131
rect 22661 21097 22695 21131
rect 22695 21097 22704 21131
rect 22652 21088 22704 21097
rect 23940 21088 23992 21140
rect 9864 21020 9916 21072
rect 10140 21020 10192 21072
rect 15476 21063 15528 21072
rect 15476 21029 15485 21063
rect 15485 21029 15519 21063
rect 15519 21029 15528 21063
rect 15476 21020 15528 21029
rect 9772 20952 9824 21004
rect 11244 20995 11296 21004
rect 7104 20884 7156 20936
rect 8300 20927 8352 20936
rect 8300 20893 8309 20927
rect 8309 20893 8343 20927
rect 8343 20893 8352 20927
rect 8300 20884 8352 20893
rect 8484 20927 8536 20936
rect 8484 20893 8493 20927
rect 8493 20893 8527 20927
rect 8527 20893 8536 20927
rect 8484 20884 8536 20893
rect 11244 20961 11253 20995
rect 11253 20961 11287 20995
rect 11287 20961 11296 20995
rect 11244 20952 11296 20961
rect 12256 20952 12308 21004
rect 14740 20952 14792 21004
rect 16396 20995 16448 21004
rect 16396 20961 16430 20995
rect 16430 20961 16448 20995
rect 16396 20952 16448 20961
rect 17960 20952 18012 21004
rect 19064 20995 19116 21004
rect 19064 20961 19073 20995
rect 19073 20961 19107 20995
rect 19107 20961 19116 20995
rect 19064 20952 19116 20961
rect 11520 20927 11572 20936
rect 11520 20893 11529 20927
rect 11529 20893 11563 20927
rect 11563 20893 11572 20927
rect 11520 20884 11572 20893
rect 13176 20884 13228 20936
rect 13360 20884 13412 20936
rect 13728 20927 13780 20936
rect 13728 20893 13737 20927
rect 13737 20893 13771 20927
rect 13771 20893 13780 20927
rect 13728 20884 13780 20893
rect 10784 20816 10836 20868
rect 19156 20927 19208 20936
rect 19156 20893 19165 20927
rect 19165 20893 19199 20927
rect 19199 20893 19208 20927
rect 19156 20884 19208 20893
rect 22468 20995 22520 21004
rect 22468 20961 22477 20995
rect 22477 20961 22511 20995
rect 22511 20961 22520 20995
rect 22468 20952 22520 20961
rect 23940 20995 23992 21004
rect 23940 20961 23949 20995
rect 23949 20961 23983 20995
rect 23983 20961 23992 20995
rect 23940 20952 23992 20961
rect 25136 20995 25188 21004
rect 25136 20961 25145 20995
rect 25145 20961 25179 20995
rect 25179 20961 25188 20995
rect 25136 20952 25188 20961
rect 21364 20927 21416 20936
rect 21364 20893 21373 20927
rect 21373 20893 21407 20927
rect 21407 20893 21416 20927
rect 21364 20884 21416 20893
rect 20812 20816 20864 20868
rect 20996 20816 21048 20868
rect 22008 20884 22060 20936
rect 23664 20884 23716 20936
rect 24860 20884 24912 20936
rect 9680 20791 9732 20800
rect 9680 20757 9689 20791
rect 9689 20757 9723 20791
rect 9723 20757 9732 20791
rect 9680 20748 9732 20757
rect 12532 20791 12584 20800
rect 12532 20757 12541 20791
rect 12541 20757 12575 20791
rect 12575 20757 12584 20791
rect 12532 20748 12584 20757
rect 13084 20791 13136 20800
rect 13084 20757 13093 20791
rect 13093 20757 13127 20791
rect 13127 20757 13136 20791
rect 13084 20748 13136 20757
rect 14464 20748 14516 20800
rect 14832 20748 14884 20800
rect 18512 20748 18564 20800
rect 20904 20791 20956 20800
rect 20904 20757 20913 20791
rect 20913 20757 20947 20791
rect 20947 20757 20956 20791
rect 20904 20748 20956 20757
rect 23480 20791 23532 20800
rect 23480 20757 23489 20791
rect 23489 20757 23523 20791
rect 23523 20757 23532 20791
rect 23480 20748 23532 20757
rect 25320 20791 25372 20800
rect 25320 20757 25329 20791
rect 25329 20757 25363 20791
rect 25363 20757 25372 20791
rect 25320 20748 25372 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 8208 20544 8260 20596
rect 10692 20544 10744 20596
rect 17408 20587 17460 20596
rect 17408 20553 17417 20587
rect 17417 20553 17451 20587
rect 17451 20553 17460 20587
rect 17408 20544 17460 20553
rect 20720 20544 20772 20596
rect 21364 20544 21416 20596
rect 21916 20587 21968 20596
rect 21916 20553 21925 20587
rect 21925 20553 21959 20587
rect 21959 20553 21968 20587
rect 21916 20544 21968 20553
rect 22652 20587 22704 20596
rect 22652 20553 22661 20587
rect 22661 20553 22695 20587
rect 22695 20553 22704 20587
rect 22652 20544 22704 20553
rect 23940 20544 23992 20596
rect 24860 20544 24912 20596
rect 25136 20544 25188 20596
rect 11244 20476 11296 20528
rect 9680 20408 9732 20460
rect 10140 20451 10192 20460
rect 10140 20417 10149 20451
rect 10149 20417 10183 20451
rect 10183 20417 10192 20451
rect 10140 20408 10192 20417
rect 10232 20451 10284 20460
rect 10232 20417 10241 20451
rect 10241 20417 10275 20451
rect 10275 20417 10284 20451
rect 10784 20451 10836 20460
rect 10232 20408 10284 20417
rect 10784 20417 10793 20451
rect 10793 20417 10827 20451
rect 10827 20417 10836 20451
rect 10784 20408 10836 20417
rect 20996 20476 21048 20528
rect 21548 20451 21600 20460
rect 9588 20383 9640 20392
rect 9588 20349 9597 20383
rect 9597 20349 9631 20383
rect 9631 20349 9640 20383
rect 9588 20340 9640 20349
rect 10692 20340 10744 20392
rect 10232 20272 10284 20324
rect 12532 20340 12584 20392
rect 13820 20340 13872 20392
rect 14924 20383 14976 20392
rect 14924 20349 14933 20383
rect 14933 20349 14967 20383
rect 14967 20349 14976 20383
rect 14924 20340 14976 20349
rect 18052 20383 18104 20392
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 21548 20417 21557 20451
rect 21557 20417 21591 20451
rect 21591 20417 21600 20451
rect 22468 20476 22520 20528
rect 21548 20408 21600 20417
rect 23480 20408 23532 20460
rect 18696 20340 18748 20392
rect 19064 20340 19116 20392
rect 22836 20340 22888 20392
rect 12808 20272 12860 20324
rect 15844 20272 15896 20324
rect 16672 20272 16724 20324
rect 8300 20247 8352 20256
rect 8300 20213 8309 20247
rect 8309 20213 8343 20247
rect 8343 20213 8352 20247
rect 8300 20204 8352 20213
rect 8484 20204 8536 20256
rect 9036 20204 9088 20256
rect 11428 20204 11480 20256
rect 12256 20204 12308 20256
rect 13820 20247 13872 20256
rect 13820 20213 13829 20247
rect 13829 20213 13863 20247
rect 13863 20213 13872 20247
rect 13820 20204 13872 20213
rect 16396 20204 16448 20256
rect 17040 20272 17092 20324
rect 19156 20272 19208 20324
rect 20904 20272 20956 20324
rect 25228 20383 25280 20392
rect 25228 20349 25237 20383
rect 25237 20349 25271 20383
rect 25271 20349 25280 20383
rect 25228 20340 25280 20349
rect 17868 20247 17920 20256
rect 17868 20213 17877 20247
rect 17877 20213 17911 20247
rect 17911 20213 17920 20247
rect 17868 20204 17920 20213
rect 18328 20204 18380 20256
rect 23848 20204 23900 20256
rect 24032 20247 24084 20256
rect 24032 20213 24041 20247
rect 24041 20213 24075 20247
rect 24075 20213 24084 20247
rect 24032 20204 24084 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 9864 20043 9916 20052
rect 9864 20009 9873 20043
rect 9873 20009 9907 20043
rect 9907 20009 9916 20043
rect 9864 20000 9916 20009
rect 10140 20000 10192 20052
rect 13176 20043 13228 20052
rect 13176 20009 13185 20043
rect 13185 20009 13219 20043
rect 13219 20009 13228 20043
rect 13176 20000 13228 20009
rect 16672 20043 16724 20052
rect 16672 20009 16681 20043
rect 16681 20009 16715 20043
rect 16715 20009 16724 20043
rect 16672 20000 16724 20009
rect 16764 20000 16816 20052
rect 20720 20043 20772 20052
rect 10876 19975 10928 19984
rect 10876 19941 10910 19975
rect 10910 19941 10928 19975
rect 10876 19932 10928 19941
rect 13084 19932 13136 19984
rect 16580 19932 16632 19984
rect 19156 19975 19208 19984
rect 19156 19941 19165 19975
rect 19165 19941 19199 19975
rect 19199 19941 19208 19975
rect 19156 19932 19208 19941
rect 20720 20009 20729 20043
rect 20729 20009 20763 20043
rect 20763 20009 20772 20043
rect 20720 20000 20772 20009
rect 20904 20000 20956 20052
rect 21272 20000 21324 20052
rect 22008 20000 22060 20052
rect 22100 20000 22152 20052
rect 21548 19932 21600 19984
rect 13728 19907 13780 19916
rect 13728 19873 13737 19907
rect 13737 19873 13771 19907
rect 13771 19873 13780 19907
rect 13728 19864 13780 19873
rect 9680 19796 9732 19848
rect 13452 19796 13504 19848
rect 15384 19864 15436 19916
rect 18052 19864 18104 19916
rect 19340 19907 19392 19916
rect 19340 19873 19349 19907
rect 19349 19873 19383 19907
rect 19383 19873 19392 19907
rect 19340 19864 19392 19873
rect 20536 19864 20588 19916
rect 20904 19907 20956 19916
rect 20904 19873 20913 19907
rect 20913 19873 20947 19907
rect 20947 19873 20956 19907
rect 20904 19864 20956 19873
rect 23940 20000 23992 20052
rect 23480 19932 23532 19984
rect 25228 20000 25280 20052
rect 23204 19864 23256 19916
rect 13912 19728 13964 19780
rect 14924 19728 14976 19780
rect 17684 19796 17736 19848
rect 18328 19839 18380 19848
rect 18328 19805 18337 19839
rect 18337 19805 18371 19839
rect 18371 19805 18380 19839
rect 18328 19796 18380 19805
rect 19616 19839 19668 19848
rect 19616 19805 19625 19839
rect 19625 19805 19659 19839
rect 19659 19805 19668 19839
rect 19616 19796 19668 19805
rect 23296 19728 23348 19780
rect 11888 19660 11940 19712
rect 12808 19703 12860 19712
rect 12808 19669 12817 19703
rect 12817 19669 12851 19703
rect 12851 19669 12860 19703
rect 12808 19660 12860 19669
rect 13360 19703 13412 19712
rect 13360 19669 13369 19703
rect 13369 19669 13403 19703
rect 13403 19669 13412 19703
rect 13360 19660 13412 19669
rect 14832 19660 14884 19712
rect 18696 19660 18748 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 9036 19499 9088 19508
rect 9036 19465 9045 19499
rect 9045 19465 9079 19499
rect 9079 19465 9088 19499
rect 9036 19456 9088 19465
rect 10876 19456 10928 19508
rect 13084 19456 13136 19508
rect 15384 19499 15436 19508
rect 15384 19465 15393 19499
rect 15393 19465 15427 19499
rect 15427 19465 15436 19499
rect 15384 19456 15436 19465
rect 15752 19456 15804 19508
rect 16212 19456 16264 19508
rect 16764 19456 16816 19508
rect 17408 19499 17460 19508
rect 17408 19465 17417 19499
rect 17417 19465 17451 19499
rect 17451 19465 17460 19499
rect 17408 19456 17460 19465
rect 20812 19499 20864 19508
rect 20812 19465 20821 19499
rect 20821 19465 20855 19499
rect 20855 19465 20864 19499
rect 20812 19456 20864 19465
rect 21548 19456 21600 19508
rect 23204 19456 23256 19508
rect 24860 19456 24912 19508
rect 10968 19320 11020 19372
rect 17040 19363 17092 19372
rect 17040 19329 17049 19363
rect 17049 19329 17083 19363
rect 17083 19329 17092 19363
rect 17040 19320 17092 19329
rect 22008 19388 22060 19440
rect 23296 19388 23348 19440
rect 21824 19320 21876 19372
rect 22928 19320 22980 19372
rect 7656 19295 7708 19304
rect 7656 19261 7665 19295
rect 7665 19261 7699 19295
rect 7699 19261 7708 19295
rect 7656 19252 7708 19261
rect 12808 19252 12860 19304
rect 13912 19252 13964 19304
rect 17316 19252 17368 19304
rect 17684 19252 17736 19304
rect 18512 19295 18564 19304
rect 18512 19261 18521 19295
rect 18521 19261 18555 19295
rect 18555 19261 18564 19295
rect 18512 19252 18564 19261
rect 19800 19295 19852 19304
rect 19800 19261 19809 19295
rect 19809 19261 19843 19295
rect 19843 19261 19852 19295
rect 19800 19252 19852 19261
rect 10140 19159 10192 19168
rect 10140 19125 10149 19159
rect 10149 19125 10183 19159
rect 10183 19125 10192 19159
rect 10140 19116 10192 19125
rect 10692 19184 10744 19236
rect 13636 19227 13688 19236
rect 13636 19193 13670 19227
rect 13670 19193 13688 19227
rect 13636 19184 13688 19193
rect 16120 19184 16172 19236
rect 18420 19227 18472 19236
rect 18420 19193 18429 19227
rect 18429 19193 18463 19227
rect 18463 19193 18472 19227
rect 18420 19184 18472 19193
rect 10784 19116 10836 19168
rect 12164 19116 12216 19168
rect 16396 19116 16448 19168
rect 18052 19159 18104 19168
rect 18052 19125 18061 19159
rect 18061 19125 18095 19159
rect 18095 19125 18104 19159
rect 18052 19116 18104 19125
rect 20904 19116 20956 19168
rect 22192 19252 22244 19304
rect 23204 19252 23256 19304
rect 23296 19252 23348 19304
rect 24952 19252 25004 19304
rect 22560 19184 22612 19236
rect 23480 19184 23532 19236
rect 21824 19116 21876 19168
rect 22008 19116 22060 19168
rect 22652 19159 22704 19168
rect 22652 19125 22661 19159
rect 22661 19125 22695 19159
rect 22695 19125 22704 19159
rect 22652 19116 22704 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 10784 18912 10836 18964
rect 13452 18955 13504 18964
rect 13452 18921 13461 18955
rect 13461 18921 13495 18955
rect 13495 18921 13504 18955
rect 13452 18912 13504 18921
rect 14464 18912 14516 18964
rect 15292 18912 15344 18964
rect 15752 18955 15804 18964
rect 15752 18921 15761 18955
rect 15761 18921 15795 18955
rect 15795 18921 15804 18955
rect 15752 18912 15804 18921
rect 18052 18912 18104 18964
rect 19340 18912 19392 18964
rect 21640 18955 21692 18964
rect 21640 18921 21649 18955
rect 21649 18921 21683 18955
rect 21683 18921 21692 18955
rect 21640 18912 21692 18921
rect 22744 18955 22796 18964
rect 22744 18921 22753 18955
rect 22753 18921 22787 18955
rect 22787 18921 22796 18955
rect 22744 18912 22796 18921
rect 23480 18955 23532 18964
rect 23480 18921 23489 18955
rect 23489 18921 23523 18955
rect 23523 18921 23532 18955
rect 23480 18912 23532 18921
rect 23664 18955 23716 18964
rect 23664 18921 23673 18955
rect 23673 18921 23707 18955
rect 23707 18921 23716 18955
rect 23664 18912 23716 18921
rect 21548 18844 21600 18896
rect 9496 18819 9548 18828
rect 9496 18785 9505 18819
rect 9505 18785 9539 18819
rect 9539 18785 9548 18819
rect 9496 18776 9548 18785
rect 9956 18819 10008 18828
rect 9956 18785 9990 18819
rect 9990 18785 10008 18819
rect 9956 18776 10008 18785
rect 12256 18776 12308 18828
rect 9680 18751 9732 18760
rect 7656 18640 7708 18692
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 10968 18640 11020 18692
rect 11152 18572 11204 18624
rect 12716 18751 12768 18760
rect 12716 18717 12725 18751
rect 12725 18717 12759 18751
rect 12759 18717 12768 18751
rect 12716 18708 12768 18717
rect 14280 18708 14332 18760
rect 13820 18615 13872 18624
rect 13820 18581 13829 18615
rect 13829 18581 13863 18615
rect 13863 18581 13872 18615
rect 13820 18572 13872 18581
rect 13912 18572 13964 18624
rect 14832 18572 14884 18624
rect 16764 18776 16816 18828
rect 17592 18819 17644 18828
rect 17592 18785 17601 18819
rect 17601 18785 17635 18819
rect 17635 18785 17644 18819
rect 17592 18776 17644 18785
rect 18144 18776 18196 18828
rect 19248 18819 19300 18828
rect 19248 18785 19257 18819
rect 19257 18785 19291 18819
rect 19291 18785 19300 18819
rect 19248 18776 19300 18785
rect 15844 18751 15896 18760
rect 15844 18717 15853 18751
rect 15853 18717 15887 18751
rect 15887 18717 15896 18751
rect 15844 18708 15896 18717
rect 17684 18751 17736 18760
rect 17684 18717 17693 18751
rect 17693 18717 17727 18751
rect 17727 18717 17736 18751
rect 17684 18708 17736 18717
rect 18788 18751 18840 18760
rect 15292 18683 15344 18692
rect 15292 18649 15301 18683
rect 15301 18649 15335 18683
rect 15335 18649 15344 18683
rect 15292 18640 15344 18649
rect 16672 18640 16724 18692
rect 18236 18640 18288 18692
rect 18788 18717 18797 18751
rect 18797 18717 18831 18751
rect 18831 18717 18840 18751
rect 19524 18751 19576 18760
rect 18788 18708 18840 18717
rect 19524 18717 19533 18751
rect 19533 18717 19567 18751
rect 19567 18717 19576 18751
rect 19524 18708 19576 18717
rect 21088 18776 21140 18828
rect 22560 18819 22612 18828
rect 22560 18785 22569 18819
rect 22569 18785 22603 18819
rect 22603 18785 22612 18819
rect 22560 18776 22612 18785
rect 23296 18776 23348 18828
rect 21180 18708 21232 18760
rect 23480 18708 23532 18760
rect 25228 18819 25280 18828
rect 25228 18785 25237 18819
rect 25237 18785 25271 18819
rect 25271 18785 25280 18819
rect 25228 18776 25280 18785
rect 16120 18572 16172 18624
rect 17224 18615 17276 18624
rect 17224 18581 17233 18615
rect 17233 18581 17267 18615
rect 17267 18581 17276 18615
rect 17224 18572 17276 18581
rect 18420 18615 18472 18624
rect 18420 18581 18429 18615
rect 18429 18581 18463 18615
rect 18463 18581 18472 18615
rect 18420 18572 18472 18581
rect 18880 18615 18932 18624
rect 18880 18581 18889 18615
rect 18889 18581 18923 18615
rect 18923 18581 18932 18615
rect 18880 18572 18932 18581
rect 20076 18572 20128 18624
rect 20536 18572 20588 18624
rect 24952 18572 25004 18624
rect 25412 18615 25464 18624
rect 25412 18581 25421 18615
rect 25421 18581 25455 18615
rect 25455 18581 25464 18615
rect 25412 18572 25464 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 10692 18368 10744 18420
rect 11888 18411 11940 18420
rect 9956 18232 10008 18284
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 12256 18411 12308 18420
rect 12256 18377 12265 18411
rect 12265 18377 12299 18411
rect 12299 18377 12308 18411
rect 12256 18368 12308 18377
rect 13452 18368 13504 18420
rect 12716 18232 12768 18284
rect 14832 18368 14884 18420
rect 15476 18368 15528 18420
rect 15844 18368 15896 18420
rect 19524 18368 19576 18420
rect 20720 18411 20772 18420
rect 20720 18377 20729 18411
rect 20729 18377 20763 18411
rect 20763 18377 20772 18411
rect 20720 18368 20772 18377
rect 22100 18411 22152 18420
rect 22100 18377 22109 18411
rect 22109 18377 22143 18411
rect 22143 18377 22152 18411
rect 22100 18368 22152 18377
rect 25228 18368 25280 18420
rect 14004 18300 14056 18352
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 14464 18164 14516 18216
rect 12716 18139 12768 18148
rect 12716 18105 12725 18139
rect 12725 18105 12759 18139
rect 12759 18105 12768 18139
rect 12716 18096 12768 18105
rect 11336 18028 11388 18080
rect 11520 18028 11572 18080
rect 14188 18071 14240 18080
rect 14188 18037 14197 18071
rect 14197 18037 14231 18071
rect 14231 18037 14240 18071
rect 14188 18028 14240 18037
rect 14464 18028 14516 18080
rect 16948 18232 17000 18284
rect 17408 18232 17460 18284
rect 18236 18232 18288 18284
rect 21364 18343 21416 18352
rect 21364 18309 21373 18343
rect 21373 18309 21407 18343
rect 21407 18309 21416 18343
rect 21364 18300 21416 18309
rect 22468 18232 22520 18284
rect 23296 18232 23348 18284
rect 16580 18164 16632 18216
rect 17684 18164 17736 18216
rect 15844 18096 15896 18148
rect 15384 18071 15436 18080
rect 15384 18037 15393 18071
rect 15393 18037 15427 18071
rect 15427 18037 15436 18071
rect 15384 18028 15436 18037
rect 16948 18071 17000 18080
rect 16948 18037 16957 18071
rect 16957 18037 16991 18071
rect 16991 18037 17000 18071
rect 16948 18028 17000 18037
rect 18420 18096 18472 18148
rect 20996 18096 21048 18148
rect 17684 18028 17736 18080
rect 19248 18028 19300 18080
rect 21088 18071 21140 18080
rect 21088 18037 21097 18071
rect 21097 18037 21131 18071
rect 21131 18037 21140 18071
rect 21088 18028 21140 18037
rect 21180 18028 21232 18080
rect 22100 18164 22152 18216
rect 23296 18096 23348 18148
rect 24492 18164 24544 18216
rect 24860 18164 24912 18216
rect 24952 18096 25004 18148
rect 21916 18028 21968 18080
rect 23480 18071 23532 18080
rect 23480 18037 23489 18071
rect 23489 18037 23523 18071
rect 23523 18037 23532 18071
rect 23480 18028 23532 18037
rect 25136 18028 25188 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 9496 17824 9548 17876
rect 10968 17824 11020 17876
rect 12072 17867 12124 17876
rect 12072 17833 12081 17867
rect 12081 17833 12115 17867
rect 12115 17833 12124 17867
rect 12072 17824 12124 17833
rect 12440 17824 12492 17876
rect 14188 17824 14240 17876
rect 14740 17824 14792 17876
rect 18236 17824 18288 17876
rect 19340 17824 19392 17876
rect 24492 17867 24544 17876
rect 24492 17833 24501 17867
rect 24501 17833 24535 17867
rect 24535 17833 24544 17867
rect 24492 17824 24544 17833
rect 25228 17867 25280 17876
rect 25228 17833 25237 17867
rect 25237 17833 25271 17867
rect 25271 17833 25280 17867
rect 25228 17824 25280 17833
rect 10140 17756 10192 17808
rect 14372 17756 14424 17808
rect 9864 17688 9916 17740
rect 10784 17731 10836 17740
rect 10784 17697 10793 17731
rect 10793 17697 10827 17731
rect 10827 17697 10836 17731
rect 10784 17688 10836 17697
rect 12900 17688 12952 17740
rect 13084 17688 13136 17740
rect 14280 17688 14332 17740
rect 14740 17688 14792 17740
rect 15292 17688 15344 17740
rect 16672 17756 16724 17808
rect 15844 17688 15896 17740
rect 17132 17688 17184 17740
rect 18328 17688 18380 17740
rect 21180 17731 21232 17740
rect 21180 17697 21214 17731
rect 21214 17697 21232 17731
rect 21180 17688 21232 17697
rect 22652 17688 22704 17740
rect 24860 17688 24912 17740
rect 25044 17731 25096 17740
rect 25044 17697 25053 17731
rect 25053 17697 25087 17731
rect 25087 17697 25096 17731
rect 25044 17688 25096 17697
rect 10968 17663 11020 17672
rect 10968 17629 10977 17663
rect 10977 17629 11011 17663
rect 11011 17629 11020 17663
rect 10968 17620 11020 17629
rect 12256 17620 12308 17672
rect 13636 17620 13688 17672
rect 14832 17620 14884 17672
rect 18236 17663 18288 17672
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 9680 17484 9732 17536
rect 10876 17484 10928 17536
rect 12164 17484 12216 17536
rect 16764 17552 16816 17604
rect 17868 17552 17920 17604
rect 15752 17484 15804 17536
rect 16028 17484 16080 17536
rect 16396 17484 16448 17536
rect 17132 17527 17184 17536
rect 17132 17493 17141 17527
rect 17141 17493 17175 17527
rect 17175 17493 17184 17527
rect 17132 17484 17184 17493
rect 20076 17484 20128 17536
rect 23664 17620 23716 17672
rect 24676 17620 24728 17672
rect 25136 17620 25188 17672
rect 23480 17595 23532 17604
rect 23480 17561 23489 17595
rect 23489 17561 23523 17595
rect 23523 17561 23532 17595
rect 23480 17552 23532 17561
rect 22284 17527 22336 17536
rect 22284 17493 22293 17527
rect 22293 17493 22327 17527
rect 22327 17493 22336 17527
rect 22284 17484 22336 17493
rect 23388 17527 23440 17536
rect 23388 17493 23397 17527
rect 23397 17493 23431 17527
rect 23431 17493 23440 17527
rect 23388 17484 23440 17493
rect 24952 17527 25004 17536
rect 24952 17493 24961 17527
rect 24961 17493 24995 17527
rect 24995 17493 25004 17527
rect 24952 17484 25004 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 10968 17280 11020 17332
rect 12256 17280 12308 17332
rect 14740 17323 14792 17332
rect 14740 17289 14749 17323
rect 14749 17289 14783 17323
rect 14783 17289 14792 17323
rect 14740 17280 14792 17289
rect 16488 17280 16540 17332
rect 21180 17280 21232 17332
rect 21456 17280 21508 17332
rect 22652 17323 22704 17332
rect 22652 17289 22661 17323
rect 22661 17289 22695 17323
rect 22695 17289 22704 17323
rect 22652 17280 22704 17289
rect 23664 17280 23716 17332
rect 25136 17323 25188 17332
rect 25136 17289 25145 17323
rect 25145 17289 25179 17323
rect 25179 17289 25188 17323
rect 25136 17280 25188 17289
rect 10784 17255 10836 17264
rect 10784 17221 10793 17255
rect 10793 17221 10827 17255
rect 10827 17221 10836 17255
rect 10784 17212 10836 17221
rect 10140 17144 10192 17196
rect 11336 17187 11388 17196
rect 11336 17153 11345 17187
rect 11345 17153 11379 17187
rect 11379 17153 11388 17187
rect 11336 17144 11388 17153
rect 12164 17144 12216 17196
rect 15384 17144 15436 17196
rect 17868 17212 17920 17264
rect 11060 17119 11112 17128
rect 11060 17085 11069 17119
rect 11069 17085 11103 17119
rect 11103 17085 11112 17119
rect 11060 17076 11112 17085
rect 17132 17144 17184 17196
rect 18052 17144 18104 17196
rect 18880 17187 18932 17196
rect 18880 17153 18889 17187
rect 18889 17153 18923 17187
rect 18923 17153 18932 17187
rect 18880 17144 18932 17153
rect 17960 17076 18012 17128
rect 18236 17076 18288 17128
rect 18604 17119 18656 17128
rect 18604 17085 18613 17119
rect 18613 17085 18647 17119
rect 18647 17085 18656 17119
rect 18604 17076 18656 17085
rect 19340 17076 19392 17128
rect 20076 17076 20128 17128
rect 23388 17144 23440 17196
rect 23664 17144 23716 17196
rect 24216 17187 24268 17196
rect 24216 17153 24225 17187
rect 24225 17153 24259 17187
rect 24259 17153 24268 17187
rect 24216 17144 24268 17153
rect 23480 17076 23532 17128
rect 25228 17119 25280 17128
rect 25228 17085 25237 17119
rect 25237 17085 25271 17119
rect 25271 17085 25280 17119
rect 25228 17076 25280 17085
rect 13176 17008 13228 17060
rect 19156 17008 19208 17060
rect 20352 17008 20404 17060
rect 25504 17051 25556 17060
rect 25504 17017 25513 17051
rect 25513 17017 25547 17051
rect 25547 17017 25556 17051
rect 25504 17008 25556 17017
rect 14188 16940 14240 16992
rect 14280 16940 14332 16992
rect 15844 16983 15896 16992
rect 15844 16949 15853 16983
rect 15853 16949 15887 16983
rect 15887 16949 15896 16983
rect 15844 16940 15896 16949
rect 16396 16983 16448 16992
rect 16396 16949 16405 16983
rect 16405 16949 16439 16983
rect 16439 16949 16448 16983
rect 16396 16940 16448 16949
rect 18512 16940 18564 16992
rect 18696 16983 18748 16992
rect 18696 16949 18705 16983
rect 18705 16949 18739 16983
rect 18739 16949 18748 16983
rect 18696 16940 18748 16949
rect 19248 16983 19300 16992
rect 19248 16949 19257 16983
rect 19257 16949 19291 16983
rect 19291 16949 19300 16983
rect 19248 16940 19300 16949
rect 22744 16983 22796 16992
rect 22744 16949 22753 16983
rect 22753 16949 22787 16983
rect 22787 16949 22796 16983
rect 22744 16940 22796 16949
rect 23756 16940 23808 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 10784 16736 10836 16788
rect 11060 16736 11112 16788
rect 13176 16779 13228 16788
rect 13176 16745 13185 16779
rect 13185 16745 13219 16779
rect 13219 16745 13228 16779
rect 13176 16736 13228 16745
rect 13636 16736 13688 16788
rect 12256 16668 12308 16720
rect 14004 16736 14056 16788
rect 15292 16736 15344 16788
rect 16396 16736 16448 16788
rect 17868 16736 17920 16788
rect 18236 16779 18288 16788
rect 18236 16745 18245 16779
rect 18245 16745 18279 16779
rect 18279 16745 18288 16779
rect 18236 16736 18288 16745
rect 18328 16736 18380 16788
rect 18604 16779 18656 16788
rect 18604 16745 18613 16779
rect 18613 16745 18647 16779
rect 18647 16745 18656 16779
rect 18604 16736 18656 16745
rect 19248 16779 19300 16788
rect 19248 16745 19257 16779
rect 19257 16745 19291 16779
rect 19291 16745 19300 16779
rect 19248 16736 19300 16745
rect 20352 16779 20404 16788
rect 20352 16745 20361 16779
rect 20361 16745 20395 16779
rect 20395 16745 20404 16779
rect 20352 16736 20404 16745
rect 22284 16779 22336 16788
rect 22284 16745 22293 16779
rect 22293 16745 22327 16779
rect 22327 16745 22336 16779
rect 22284 16736 22336 16745
rect 22744 16736 22796 16788
rect 24216 16736 24268 16788
rect 25044 16779 25096 16788
rect 25044 16745 25053 16779
rect 25053 16745 25087 16779
rect 25087 16745 25096 16779
rect 25044 16736 25096 16745
rect 25412 16779 25464 16788
rect 25412 16745 25421 16779
rect 25421 16745 25455 16779
rect 25455 16745 25464 16779
rect 25412 16736 25464 16745
rect 10968 16600 11020 16652
rect 11888 16600 11940 16652
rect 16120 16668 16172 16720
rect 16948 16668 17000 16720
rect 17776 16668 17828 16720
rect 18512 16668 18564 16720
rect 21732 16668 21784 16720
rect 14004 16643 14056 16652
rect 14004 16609 14013 16643
rect 14013 16609 14047 16643
rect 14047 16609 14056 16643
rect 15476 16643 15528 16652
rect 14004 16600 14056 16609
rect 15476 16609 15485 16643
rect 15485 16609 15519 16643
rect 15519 16609 15528 16643
rect 15476 16600 15528 16609
rect 15844 16600 15896 16652
rect 13268 16532 13320 16584
rect 13728 16532 13780 16584
rect 14188 16575 14240 16584
rect 14188 16541 14197 16575
rect 14197 16541 14231 16575
rect 14231 16541 14240 16575
rect 14188 16532 14240 16541
rect 16028 16532 16080 16584
rect 18052 16600 18104 16652
rect 19156 16643 19208 16652
rect 19156 16609 19165 16643
rect 19165 16609 19199 16643
rect 19199 16609 19208 16643
rect 19156 16600 19208 16609
rect 24952 16668 25004 16720
rect 17500 16532 17552 16584
rect 17868 16575 17920 16584
rect 17868 16541 17877 16575
rect 17877 16541 17911 16575
rect 17911 16541 17920 16575
rect 17868 16532 17920 16541
rect 18880 16464 18932 16516
rect 11152 16396 11204 16448
rect 12532 16439 12584 16448
rect 12532 16405 12541 16439
rect 12541 16405 12575 16439
rect 12575 16405 12584 16439
rect 12532 16396 12584 16405
rect 13636 16439 13688 16448
rect 13636 16405 13645 16439
rect 13645 16405 13679 16439
rect 13679 16405 13688 16439
rect 13636 16396 13688 16405
rect 14464 16396 14516 16448
rect 18788 16439 18840 16448
rect 18788 16405 18797 16439
rect 18797 16405 18831 16439
rect 18831 16405 18840 16439
rect 18788 16396 18840 16405
rect 20536 16396 20588 16448
rect 23020 16643 23072 16652
rect 23020 16609 23054 16643
rect 23054 16609 23072 16643
rect 23020 16600 23072 16609
rect 25504 16600 25556 16652
rect 25964 16600 26016 16652
rect 21364 16575 21416 16584
rect 21364 16541 21373 16575
rect 21373 16541 21407 16575
rect 21407 16541 21416 16575
rect 21364 16532 21416 16541
rect 21456 16575 21508 16584
rect 21456 16541 21465 16575
rect 21465 16541 21499 16575
rect 21499 16541 21508 16575
rect 21456 16532 21508 16541
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 10784 16235 10836 16244
rect 10784 16201 10793 16235
rect 10793 16201 10827 16235
rect 10827 16201 10836 16235
rect 10784 16192 10836 16201
rect 11888 16235 11940 16244
rect 11888 16201 11897 16235
rect 11897 16201 11931 16235
rect 11931 16201 11940 16235
rect 11888 16192 11940 16201
rect 13728 16235 13780 16244
rect 13728 16201 13737 16235
rect 13737 16201 13771 16235
rect 13771 16201 13780 16235
rect 13728 16192 13780 16201
rect 17500 16235 17552 16244
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 17776 16235 17828 16244
rect 17776 16201 17785 16235
rect 17785 16201 17819 16235
rect 17819 16201 17828 16235
rect 17776 16192 17828 16201
rect 19984 16192 20036 16244
rect 20352 16192 20404 16244
rect 21548 16192 21600 16244
rect 23480 16235 23532 16244
rect 23480 16201 23489 16235
rect 23489 16201 23523 16235
rect 23523 16201 23532 16235
rect 23480 16192 23532 16201
rect 23664 16235 23716 16244
rect 23664 16201 23673 16235
rect 23673 16201 23707 16235
rect 23707 16201 23716 16235
rect 23664 16192 23716 16201
rect 25964 16235 26016 16244
rect 25964 16201 25973 16235
rect 25973 16201 26007 16235
rect 26007 16201 26016 16235
rect 25964 16192 26016 16201
rect 10876 16124 10928 16176
rect 11152 16056 11204 16108
rect 12532 16056 12584 16108
rect 12900 16056 12952 16108
rect 13084 15988 13136 16040
rect 10876 15852 10928 15904
rect 17684 16124 17736 16176
rect 16856 16099 16908 16108
rect 16856 16065 16865 16099
rect 16865 16065 16899 16099
rect 16899 16065 16908 16099
rect 16856 16056 16908 16065
rect 18512 16099 18564 16108
rect 18512 16065 18521 16099
rect 18521 16065 18555 16099
rect 18555 16065 18564 16099
rect 18512 16056 18564 16065
rect 18604 16099 18656 16108
rect 18604 16065 18613 16099
rect 18613 16065 18647 16099
rect 18647 16065 18656 16099
rect 18604 16056 18656 16065
rect 21916 16056 21968 16108
rect 13820 15988 13872 16040
rect 14464 16031 14516 16040
rect 14464 15997 14498 16031
rect 14498 15997 14516 16031
rect 14464 15988 14516 15997
rect 16120 15988 16172 16040
rect 16672 16031 16724 16040
rect 16672 15997 16681 16031
rect 16681 15997 16715 16031
rect 16715 15997 16724 16031
rect 16672 15988 16724 15997
rect 17960 15988 18012 16040
rect 19340 15988 19392 16040
rect 22284 16031 22336 16040
rect 22284 15997 22293 16031
rect 22293 15997 22327 16031
rect 22327 15997 22336 16031
rect 22284 15988 22336 15997
rect 23020 15988 23072 16040
rect 24676 16056 24728 16108
rect 25412 16099 25464 16108
rect 25412 16065 25421 16099
rect 25421 16065 25455 16099
rect 25455 16065 25464 16099
rect 25412 16056 25464 16065
rect 14096 15920 14148 15972
rect 12716 15852 12768 15904
rect 14004 15895 14056 15904
rect 14004 15861 14013 15895
rect 14013 15861 14047 15895
rect 14047 15861 14056 15895
rect 14004 15852 14056 15861
rect 15568 15895 15620 15904
rect 15568 15861 15577 15895
rect 15577 15861 15611 15895
rect 15611 15861 15620 15895
rect 15568 15852 15620 15861
rect 16028 15852 16080 15904
rect 17960 15852 18012 15904
rect 23848 15920 23900 15972
rect 24952 15920 25004 15972
rect 22284 15852 22336 15904
rect 25044 15895 25096 15904
rect 25044 15861 25053 15895
rect 25053 15861 25087 15895
rect 25087 15861 25096 15895
rect 25044 15852 25096 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 10692 15580 10744 15632
rect 12532 15648 12584 15700
rect 12716 15648 12768 15700
rect 13084 15691 13136 15700
rect 13084 15657 13093 15691
rect 13093 15657 13127 15691
rect 13127 15657 13136 15691
rect 13084 15648 13136 15657
rect 13360 15648 13412 15700
rect 13636 15648 13688 15700
rect 14188 15691 14240 15700
rect 14188 15657 14197 15691
rect 14197 15657 14231 15691
rect 14231 15657 14240 15691
rect 14188 15648 14240 15657
rect 14464 15691 14516 15700
rect 14464 15657 14473 15691
rect 14473 15657 14507 15691
rect 14507 15657 14516 15691
rect 14464 15648 14516 15657
rect 15844 15648 15896 15700
rect 17684 15691 17736 15700
rect 17684 15657 17693 15691
rect 17693 15657 17727 15691
rect 17727 15657 17736 15691
rect 17684 15648 17736 15657
rect 18144 15691 18196 15700
rect 18144 15657 18153 15691
rect 18153 15657 18187 15691
rect 18187 15657 18196 15691
rect 18144 15648 18196 15657
rect 18880 15648 18932 15700
rect 21364 15648 21416 15700
rect 21732 15648 21784 15700
rect 22284 15648 22336 15700
rect 23848 15648 23900 15700
rect 25044 15648 25096 15700
rect 11060 15580 11112 15632
rect 16028 15580 16080 15632
rect 16672 15580 16724 15632
rect 17868 15580 17920 15632
rect 20720 15623 20772 15632
rect 12900 15555 12952 15564
rect 12900 15521 12909 15555
rect 12909 15521 12943 15555
rect 12943 15521 12952 15555
rect 12900 15512 12952 15521
rect 13176 15512 13228 15564
rect 16488 15555 16540 15564
rect 16488 15521 16497 15555
rect 16497 15521 16531 15555
rect 16531 15521 16540 15555
rect 16488 15512 16540 15521
rect 17408 15512 17460 15564
rect 20720 15589 20729 15623
rect 20729 15589 20763 15623
rect 20763 15589 20772 15623
rect 20720 15580 20772 15589
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 16304 15444 16356 15496
rect 16764 15487 16816 15496
rect 16764 15453 16773 15487
rect 16773 15453 16807 15487
rect 16807 15453 16816 15487
rect 16764 15444 16816 15453
rect 14372 15376 14424 15428
rect 17960 15376 18012 15428
rect 19984 15444 20036 15496
rect 20812 15512 20864 15564
rect 21732 15555 21784 15564
rect 21732 15521 21766 15555
rect 21766 15521 21784 15555
rect 21732 15512 21784 15521
rect 23848 15512 23900 15564
rect 20628 15444 20680 15496
rect 23480 15444 23532 15496
rect 24676 15512 24728 15564
rect 23756 15376 23808 15428
rect 10876 15308 10928 15360
rect 15752 15308 15804 15360
rect 24952 15351 25004 15360
rect 24952 15317 24961 15351
rect 24961 15317 24995 15351
rect 24995 15317 25004 15351
rect 24952 15308 25004 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 10692 15147 10744 15156
rect 10692 15113 10701 15147
rect 10701 15113 10735 15147
rect 10735 15113 10744 15147
rect 10692 15104 10744 15113
rect 13360 15104 13412 15156
rect 15384 15147 15436 15156
rect 15384 15113 15393 15147
rect 15393 15113 15427 15147
rect 15427 15113 15436 15147
rect 15384 15104 15436 15113
rect 16488 15104 16540 15156
rect 20536 15104 20588 15156
rect 23388 15104 23440 15156
rect 23756 15104 23808 15156
rect 11612 15036 11664 15088
rect 13544 15036 13596 15088
rect 12716 14968 12768 15020
rect 14372 15011 14424 15020
rect 14372 14977 14381 15011
rect 14381 14977 14415 15011
rect 14415 14977 14424 15011
rect 14372 14968 14424 14977
rect 14464 15011 14516 15020
rect 14464 14977 14473 15011
rect 14473 14977 14507 15011
rect 14507 14977 14516 15011
rect 14464 14968 14516 14977
rect 15292 14968 15344 15020
rect 12624 14900 12676 14952
rect 16764 14968 16816 15020
rect 19984 15036 20036 15088
rect 18604 15011 18656 15020
rect 18604 14977 18613 15011
rect 18613 14977 18647 15011
rect 18647 14977 18656 15011
rect 18604 14968 18656 14977
rect 20352 15011 20404 15020
rect 20352 14977 20361 15011
rect 20361 14977 20395 15011
rect 20395 14977 20404 15011
rect 20352 14968 20404 14977
rect 20812 15036 20864 15088
rect 22284 14968 22336 15020
rect 23940 14968 23992 15020
rect 10600 14832 10652 14884
rect 16948 14900 17000 14952
rect 22468 14900 22520 14952
rect 23020 14900 23072 14952
rect 23664 14900 23716 14952
rect 15568 14832 15620 14884
rect 18420 14875 18472 14884
rect 9864 14764 9916 14816
rect 18420 14841 18429 14875
rect 18429 14841 18463 14875
rect 18463 14841 18472 14875
rect 18420 14832 18472 14841
rect 20996 14875 21048 14884
rect 20996 14841 21005 14875
rect 21005 14841 21039 14875
rect 21039 14841 21048 14875
rect 20996 14832 21048 14841
rect 21180 14832 21232 14884
rect 23112 14832 23164 14884
rect 24492 14832 24544 14884
rect 24952 14832 25004 14884
rect 10968 14764 11020 14816
rect 13176 14807 13228 14816
rect 13176 14773 13185 14807
rect 13185 14773 13219 14807
rect 13219 14773 13228 14807
rect 13176 14764 13228 14773
rect 13912 14807 13964 14816
rect 13912 14773 13921 14807
rect 13921 14773 13955 14807
rect 13955 14773 13964 14807
rect 13912 14764 13964 14773
rect 17408 14807 17460 14816
rect 17408 14773 17417 14807
rect 17417 14773 17451 14807
rect 17451 14773 17460 14807
rect 17408 14764 17460 14773
rect 17776 14807 17828 14816
rect 17776 14773 17785 14807
rect 17785 14773 17819 14807
rect 17819 14773 17828 14807
rect 17776 14764 17828 14773
rect 18052 14807 18104 14816
rect 18052 14773 18061 14807
rect 18061 14773 18095 14807
rect 18095 14773 18104 14807
rect 18052 14764 18104 14773
rect 18512 14807 18564 14816
rect 18512 14773 18521 14807
rect 18521 14773 18555 14807
rect 18555 14773 18564 14807
rect 18512 14764 18564 14773
rect 20628 14764 20680 14816
rect 21272 14807 21324 14816
rect 21272 14773 21281 14807
rect 21281 14773 21315 14807
rect 21315 14773 21324 14807
rect 21272 14764 21324 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 9772 14560 9824 14612
rect 10968 14560 11020 14612
rect 11612 14603 11664 14612
rect 11612 14569 11621 14603
rect 11621 14569 11655 14603
rect 11655 14569 11664 14603
rect 11612 14560 11664 14569
rect 13912 14560 13964 14612
rect 14188 14560 14240 14612
rect 12348 14492 12400 14544
rect 15568 14560 15620 14612
rect 15844 14560 15896 14612
rect 16764 14603 16816 14612
rect 16764 14569 16773 14603
rect 16773 14569 16807 14603
rect 16807 14569 16816 14603
rect 16764 14560 16816 14569
rect 16948 14560 17000 14612
rect 10784 14467 10836 14476
rect 10784 14433 10793 14467
rect 10793 14433 10827 14467
rect 10827 14433 10836 14467
rect 10784 14424 10836 14433
rect 11612 14424 11664 14476
rect 12900 14424 12952 14476
rect 13360 14424 13412 14476
rect 13820 14424 13872 14476
rect 11060 14399 11112 14408
rect 11060 14365 11069 14399
rect 11069 14365 11103 14399
rect 11103 14365 11112 14399
rect 11060 14356 11112 14365
rect 12624 14399 12676 14408
rect 12624 14365 12633 14399
rect 12633 14365 12667 14399
rect 12667 14365 12676 14399
rect 12624 14356 12676 14365
rect 13912 14356 13964 14408
rect 12072 14331 12124 14340
rect 12072 14297 12081 14331
rect 12081 14297 12115 14331
rect 12115 14297 12124 14331
rect 12072 14288 12124 14297
rect 14372 14288 14424 14340
rect 13820 14220 13872 14272
rect 17868 14560 17920 14612
rect 18880 14560 18932 14612
rect 19984 14560 20036 14612
rect 20720 14560 20772 14612
rect 21732 14560 21784 14612
rect 23848 14603 23900 14612
rect 23848 14569 23857 14603
rect 23857 14569 23891 14603
rect 23891 14569 23900 14603
rect 23848 14560 23900 14569
rect 24860 14560 24912 14612
rect 18236 14492 18288 14544
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 15292 14288 15344 14340
rect 17868 14424 17920 14476
rect 20812 14492 20864 14544
rect 21364 14492 21416 14544
rect 22376 14492 22428 14544
rect 24952 14535 25004 14544
rect 24952 14501 24961 14535
rect 24961 14501 24995 14535
rect 24995 14501 25004 14535
rect 24952 14492 25004 14501
rect 21824 14424 21876 14476
rect 24032 14424 24084 14476
rect 17316 14356 17368 14408
rect 17684 14356 17736 14408
rect 20628 14356 20680 14408
rect 20812 14356 20864 14408
rect 21640 14356 21692 14408
rect 22284 14356 22336 14408
rect 23848 14356 23900 14408
rect 24492 14399 24544 14408
rect 24492 14365 24501 14399
rect 24501 14365 24535 14399
rect 24535 14365 24544 14399
rect 24492 14356 24544 14365
rect 23204 14288 23256 14340
rect 25504 14288 25556 14340
rect 16304 14263 16356 14272
rect 16304 14229 16313 14263
rect 16313 14229 16347 14263
rect 16347 14229 16356 14263
rect 16304 14220 16356 14229
rect 22284 14263 22336 14272
rect 22284 14229 22293 14263
rect 22293 14229 22327 14263
rect 22327 14229 22336 14263
rect 22284 14220 22336 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 11244 14016 11296 14068
rect 11612 14059 11664 14068
rect 11612 14025 11621 14059
rect 11621 14025 11655 14059
rect 11655 14025 11664 14059
rect 11612 14016 11664 14025
rect 12624 14016 12676 14068
rect 14464 14016 14516 14068
rect 15844 14016 15896 14068
rect 16396 14059 16448 14068
rect 16396 14025 16405 14059
rect 16405 14025 16439 14059
rect 16439 14025 16448 14059
rect 16396 14016 16448 14025
rect 13360 13991 13412 14000
rect 13360 13957 13369 13991
rect 13369 13957 13403 13991
rect 13403 13957 13412 13991
rect 13360 13948 13412 13957
rect 10968 13880 11020 13932
rect 13544 13923 13596 13932
rect 10140 13855 10192 13864
rect 10140 13821 10149 13855
rect 10149 13821 10183 13855
rect 10183 13821 10192 13855
rect 10140 13812 10192 13821
rect 10692 13744 10744 13796
rect 13544 13889 13553 13923
rect 13553 13889 13587 13923
rect 13587 13889 13596 13923
rect 13544 13880 13596 13889
rect 18052 14016 18104 14068
rect 18604 14016 18656 14068
rect 18880 14059 18932 14068
rect 18880 14025 18889 14059
rect 18889 14025 18923 14059
rect 18923 14025 18932 14059
rect 18880 14016 18932 14025
rect 21640 14059 21692 14068
rect 21640 14025 21649 14059
rect 21649 14025 21683 14059
rect 21683 14025 21692 14059
rect 21640 14016 21692 14025
rect 21824 14059 21876 14068
rect 21824 14025 21833 14059
rect 21833 14025 21867 14059
rect 21867 14025 21876 14059
rect 21824 14016 21876 14025
rect 23112 14059 23164 14068
rect 23112 14025 23121 14059
rect 23121 14025 23155 14059
rect 23155 14025 23164 14059
rect 23112 14016 23164 14025
rect 23848 14059 23900 14068
rect 23848 14025 23857 14059
rect 23857 14025 23891 14059
rect 23891 14025 23900 14059
rect 23848 14016 23900 14025
rect 20444 13948 20496 14000
rect 15844 13855 15896 13864
rect 15844 13821 15853 13855
rect 15853 13821 15887 13855
rect 15887 13821 15896 13855
rect 15844 13812 15896 13821
rect 13912 13744 13964 13796
rect 16580 13812 16632 13864
rect 18236 13812 18288 13864
rect 22100 13880 22152 13932
rect 23388 13880 23440 13932
rect 23664 13880 23716 13932
rect 23848 13880 23900 13932
rect 20812 13812 20864 13864
rect 21364 13855 21416 13864
rect 21364 13821 21373 13855
rect 21373 13821 21407 13855
rect 21407 13821 21416 13855
rect 21364 13812 21416 13821
rect 22284 13855 22336 13864
rect 22284 13821 22293 13855
rect 22293 13821 22327 13855
rect 22327 13821 22336 13855
rect 22284 13812 22336 13821
rect 24032 13812 24084 13864
rect 24952 13812 25004 13864
rect 19064 13744 19116 13796
rect 24400 13787 24452 13796
rect 24400 13753 24434 13787
rect 24434 13753 24452 13787
rect 24400 13744 24452 13753
rect 11704 13676 11756 13728
rect 13084 13719 13136 13728
rect 13084 13685 13093 13719
rect 13093 13685 13127 13719
rect 13127 13685 13136 13719
rect 13084 13676 13136 13685
rect 14188 13676 14240 13728
rect 22192 13719 22244 13728
rect 22192 13685 22201 13719
rect 22201 13685 22235 13719
rect 22235 13685 22244 13719
rect 22192 13676 22244 13685
rect 25504 13719 25556 13728
rect 25504 13685 25513 13719
rect 25513 13685 25547 13719
rect 25547 13685 25556 13719
rect 25504 13676 25556 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 11704 13515 11756 13524
rect 11704 13481 11713 13515
rect 11713 13481 11747 13515
rect 11747 13481 11756 13515
rect 11704 13472 11756 13481
rect 12348 13515 12400 13524
rect 12348 13481 12357 13515
rect 12357 13481 12391 13515
rect 12391 13481 12400 13515
rect 12348 13472 12400 13481
rect 13912 13472 13964 13524
rect 14832 13472 14884 13524
rect 15292 13515 15344 13524
rect 15292 13481 15301 13515
rect 15301 13481 15335 13515
rect 15335 13481 15344 13515
rect 15292 13472 15344 13481
rect 18236 13515 18288 13524
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 19064 13472 19116 13524
rect 20904 13515 20956 13524
rect 20904 13481 20913 13515
rect 20913 13481 20947 13515
rect 20947 13481 20956 13515
rect 20904 13472 20956 13481
rect 22192 13472 22244 13524
rect 23480 13515 23532 13524
rect 23480 13481 23489 13515
rect 23489 13481 23523 13515
rect 23523 13481 23532 13515
rect 23480 13472 23532 13481
rect 24676 13472 24728 13524
rect 16764 13404 16816 13456
rect 17960 13404 18012 13456
rect 19432 13404 19484 13456
rect 22100 13404 22152 13456
rect 10416 13336 10468 13388
rect 10876 13336 10928 13388
rect 12808 13379 12860 13388
rect 12808 13345 12817 13379
rect 12817 13345 12851 13379
rect 12851 13345 12860 13379
rect 12808 13336 12860 13345
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 16028 13336 16080 13388
rect 16948 13336 17000 13388
rect 19248 13336 19300 13388
rect 22376 13379 22428 13388
rect 22376 13345 22410 13379
rect 22410 13345 22428 13379
rect 24952 13379 25004 13388
rect 22376 13336 22428 13345
rect 24952 13345 24961 13379
rect 24961 13345 24995 13379
rect 24995 13345 25004 13379
rect 24952 13336 25004 13345
rect 25688 13336 25740 13388
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 9864 13268 9916 13320
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 14832 13268 14884 13320
rect 22008 13268 22060 13320
rect 25044 13311 25096 13320
rect 25044 13277 25053 13311
rect 25053 13277 25087 13311
rect 25087 13277 25096 13311
rect 25044 13268 25096 13277
rect 25504 13268 25556 13320
rect 25964 13268 26016 13320
rect 24400 13200 24452 13252
rect 25228 13200 25280 13252
rect 9864 13132 9916 13184
rect 16396 13175 16448 13184
rect 16396 13141 16405 13175
rect 16405 13141 16439 13175
rect 16439 13141 16448 13175
rect 16396 13132 16448 13141
rect 16580 13132 16632 13184
rect 16856 13132 16908 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 9680 12928 9732 12980
rect 10784 12971 10836 12980
rect 10416 12860 10468 12912
rect 10048 12792 10100 12844
rect 9496 12767 9548 12776
rect 9496 12733 9505 12767
rect 9505 12733 9539 12767
rect 9539 12733 9548 12767
rect 9496 12724 9548 12733
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 14464 12928 14516 12980
rect 14832 12928 14884 12980
rect 16028 12971 16080 12980
rect 16028 12937 16037 12971
rect 16037 12937 16071 12971
rect 16071 12937 16080 12971
rect 16028 12928 16080 12937
rect 16764 12928 16816 12980
rect 17408 12971 17460 12980
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 22192 12928 22244 12980
rect 23480 12971 23532 12980
rect 23480 12937 23489 12971
rect 23489 12937 23523 12971
rect 23523 12937 23532 12971
rect 23480 12928 23532 12937
rect 24768 12928 24820 12980
rect 25044 12928 25096 12980
rect 15200 12860 15252 12912
rect 16212 12860 16264 12912
rect 11244 12835 11296 12844
rect 11244 12801 11253 12835
rect 11253 12801 11287 12835
rect 11287 12801 11296 12835
rect 11244 12792 11296 12801
rect 11796 12835 11848 12844
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 12992 12792 13044 12844
rect 15476 12792 15528 12844
rect 12624 12724 12676 12776
rect 14556 12724 14608 12776
rect 16580 12792 16632 12844
rect 18328 12835 18380 12844
rect 18328 12801 18337 12835
rect 18337 12801 18371 12835
rect 18371 12801 18380 12835
rect 18328 12792 18380 12801
rect 19340 12792 19392 12844
rect 20720 12792 20772 12844
rect 22376 12792 22428 12844
rect 22652 12792 22704 12844
rect 25688 12903 25740 12912
rect 25688 12869 25697 12903
rect 25697 12869 25731 12903
rect 25731 12869 25740 12903
rect 25688 12860 25740 12869
rect 25964 12903 26016 12912
rect 25964 12869 25973 12903
rect 25973 12869 26007 12903
rect 26007 12869 26016 12903
rect 25964 12860 26016 12869
rect 10048 12656 10100 12708
rect 10324 12656 10376 12708
rect 15476 12656 15528 12708
rect 12256 12588 12308 12640
rect 12808 12588 12860 12640
rect 15660 12631 15712 12640
rect 15660 12597 15669 12631
rect 15669 12597 15703 12631
rect 15703 12597 15712 12631
rect 15660 12588 15712 12597
rect 16396 12724 16448 12776
rect 17868 12724 17920 12776
rect 18236 12724 18288 12776
rect 18788 12724 18840 12776
rect 20168 12724 20220 12776
rect 20904 12724 20956 12776
rect 22836 12724 22888 12776
rect 23664 12767 23716 12776
rect 23664 12733 23673 12767
rect 23673 12733 23707 12767
rect 23707 12733 23716 12767
rect 23664 12724 23716 12733
rect 17776 12699 17828 12708
rect 17776 12665 17785 12699
rect 17785 12665 17819 12699
rect 17819 12665 17828 12699
rect 17776 12656 17828 12665
rect 20720 12656 20772 12708
rect 24124 12656 24176 12708
rect 24676 12656 24728 12708
rect 16120 12588 16172 12640
rect 16764 12631 16816 12640
rect 16764 12597 16773 12631
rect 16773 12597 16807 12631
rect 16807 12597 16816 12631
rect 16764 12588 16816 12597
rect 19432 12631 19484 12640
rect 19432 12597 19441 12631
rect 19441 12597 19475 12631
rect 19475 12597 19484 12631
rect 19432 12588 19484 12597
rect 20904 12631 20956 12640
rect 20904 12597 20913 12631
rect 20913 12597 20947 12631
rect 20947 12597 20956 12631
rect 20904 12588 20956 12597
rect 22100 12588 22152 12640
rect 25228 12588 25280 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 10048 12384 10100 12436
rect 12624 12427 12676 12436
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 13452 12384 13504 12436
rect 13728 12384 13780 12436
rect 15292 12427 15344 12436
rect 15292 12393 15301 12427
rect 15301 12393 15335 12427
rect 15335 12393 15344 12427
rect 15292 12384 15344 12393
rect 15476 12384 15528 12436
rect 16488 12427 16540 12436
rect 1584 12316 1636 12368
rect 10140 12316 10192 12368
rect 15844 12316 15896 12368
rect 2044 12248 2096 12300
rect 9864 12248 9916 12300
rect 12440 12248 12492 12300
rect 13176 12291 13228 12300
rect 13176 12257 13185 12291
rect 13185 12257 13219 12291
rect 13219 12257 13228 12291
rect 13176 12248 13228 12257
rect 14372 12248 14424 12300
rect 15476 12248 15528 12300
rect 12348 12180 12400 12232
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 14188 12180 14240 12232
rect 14464 12180 14516 12232
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 16488 12393 16497 12427
rect 16497 12393 16531 12427
rect 16531 12393 16540 12427
rect 16488 12384 16540 12393
rect 17224 12427 17276 12436
rect 17224 12393 17233 12427
rect 17233 12393 17267 12427
rect 17267 12393 17276 12427
rect 17224 12384 17276 12393
rect 17500 12384 17552 12436
rect 17868 12384 17920 12436
rect 18236 12427 18288 12436
rect 18236 12393 18245 12427
rect 18245 12393 18279 12427
rect 18279 12393 18288 12427
rect 18236 12384 18288 12393
rect 19248 12427 19300 12436
rect 19248 12393 19257 12427
rect 19257 12393 19291 12427
rect 19291 12393 19300 12427
rect 19248 12384 19300 12393
rect 22100 12427 22152 12436
rect 22100 12393 22109 12427
rect 22109 12393 22143 12427
rect 22143 12393 22152 12427
rect 22100 12384 22152 12393
rect 22652 12384 22704 12436
rect 23848 12384 23900 12436
rect 20812 12316 20864 12368
rect 20996 12316 21048 12368
rect 19156 12291 19208 12300
rect 19156 12257 19165 12291
rect 19165 12257 19199 12291
rect 19199 12257 19208 12291
rect 19156 12248 19208 12257
rect 19432 12248 19484 12300
rect 19984 12248 20036 12300
rect 17316 12223 17368 12232
rect 15844 12180 15896 12189
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 17868 12180 17920 12232
rect 19524 12180 19576 12232
rect 19892 12223 19944 12232
rect 19892 12189 19901 12223
rect 19901 12189 19935 12223
rect 19935 12189 19944 12223
rect 19892 12180 19944 12189
rect 18604 12112 18656 12164
rect 20904 12248 20956 12300
rect 22008 12248 22060 12300
rect 23664 12316 23716 12368
rect 24768 12384 24820 12436
rect 25504 12316 25556 12368
rect 22468 12291 22520 12300
rect 22468 12257 22502 12291
rect 22502 12257 22520 12291
rect 22468 12248 22520 12257
rect 22928 12248 22980 12300
rect 23848 12248 23900 12300
rect 25044 12291 25096 12300
rect 25044 12257 25053 12291
rect 25053 12257 25087 12291
rect 25087 12257 25096 12291
rect 25044 12248 25096 12257
rect 25320 12248 25372 12300
rect 25228 12223 25280 12232
rect 25228 12189 25237 12223
rect 25237 12189 25271 12223
rect 25271 12189 25280 12223
rect 25228 12180 25280 12189
rect 2780 12087 2832 12096
rect 2780 12053 2789 12087
rect 2789 12053 2823 12087
rect 2823 12053 2832 12087
rect 2780 12044 2832 12053
rect 9588 12044 9640 12096
rect 11428 12044 11480 12096
rect 11796 12044 11848 12096
rect 15384 12044 15436 12096
rect 16580 12044 16632 12096
rect 18696 12087 18748 12096
rect 18696 12053 18705 12087
rect 18705 12053 18739 12087
rect 18739 12053 18748 12087
rect 18696 12044 18748 12053
rect 18788 12044 18840 12096
rect 24216 12087 24268 12096
rect 24216 12053 24225 12087
rect 24225 12053 24259 12087
rect 24259 12053 24268 12087
rect 24216 12044 24268 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 10140 11840 10192 11892
rect 13360 11840 13412 11892
rect 13544 11883 13596 11892
rect 13544 11849 13553 11883
rect 13553 11849 13587 11883
rect 13587 11849 13596 11883
rect 13544 11840 13596 11849
rect 14556 11772 14608 11824
rect 17316 11840 17368 11892
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 9588 11704 9640 11756
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 14004 11747 14056 11756
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 14832 11704 14884 11756
rect 16120 11772 16172 11824
rect 16488 11772 16540 11824
rect 16948 11772 17000 11824
rect 18788 11840 18840 11892
rect 22468 11883 22520 11892
rect 22468 11849 22477 11883
rect 22477 11849 22511 11883
rect 22511 11849 22520 11883
rect 22468 11840 22520 11849
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 20904 11704 20956 11756
rect 23664 11704 23716 11756
rect 25596 11747 25648 11756
rect 25596 11713 25605 11747
rect 25605 11713 25639 11747
rect 25639 11713 25648 11747
rect 25596 11704 25648 11713
rect 9128 11636 9180 11688
rect 13912 11679 13964 11688
rect 13912 11645 13921 11679
rect 13921 11645 13955 11679
rect 13955 11645 13964 11679
rect 13912 11636 13964 11645
rect 15384 11679 15436 11688
rect 15384 11645 15418 11679
rect 15418 11645 15436 11679
rect 15384 11636 15436 11645
rect 16120 11636 16172 11688
rect 16856 11636 16908 11688
rect 17960 11636 18012 11688
rect 19156 11636 19208 11688
rect 9956 11568 10008 11620
rect 14004 11568 14056 11620
rect 14188 11568 14240 11620
rect 18696 11568 18748 11620
rect 19248 11568 19300 11620
rect 19892 11568 19944 11620
rect 23112 11568 23164 11620
rect 24124 11636 24176 11688
rect 25044 11636 25096 11688
rect 24216 11568 24268 11620
rect 24768 11568 24820 11620
rect 2044 11543 2096 11552
rect 2044 11509 2053 11543
rect 2053 11509 2087 11543
rect 2087 11509 2096 11543
rect 2044 11500 2096 11509
rect 9220 11543 9272 11552
rect 9220 11509 9229 11543
rect 9229 11509 9263 11543
rect 9263 11509 9272 11543
rect 9220 11500 9272 11509
rect 9588 11543 9640 11552
rect 9588 11509 9597 11543
rect 9597 11509 9631 11543
rect 9631 11509 9640 11543
rect 9588 11500 9640 11509
rect 10784 11543 10836 11552
rect 10784 11509 10793 11543
rect 10793 11509 10827 11543
rect 10827 11509 10836 11543
rect 10784 11500 10836 11509
rect 10876 11500 10928 11552
rect 12532 11500 12584 11552
rect 12808 11500 12860 11552
rect 14372 11500 14424 11552
rect 15108 11500 15160 11552
rect 15844 11500 15896 11552
rect 23664 11500 23716 11552
rect 24032 11543 24084 11552
rect 24032 11509 24041 11543
rect 24041 11509 24075 11543
rect 24075 11509 24084 11543
rect 24032 11500 24084 11509
rect 25320 11500 25372 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 9128 11296 9180 11348
rect 9956 11339 10008 11348
rect 9956 11305 9965 11339
rect 9965 11305 9999 11339
rect 9999 11305 10008 11339
rect 9956 11296 10008 11305
rect 10784 11296 10836 11348
rect 13176 11296 13228 11348
rect 14464 11339 14516 11348
rect 14464 11305 14473 11339
rect 14473 11305 14507 11339
rect 14507 11305 14516 11339
rect 14464 11296 14516 11305
rect 15108 11339 15160 11348
rect 15108 11305 15117 11339
rect 15117 11305 15151 11339
rect 15151 11305 15160 11339
rect 15108 11296 15160 11305
rect 15476 11339 15528 11348
rect 15476 11305 15485 11339
rect 15485 11305 15519 11339
rect 15519 11305 15528 11339
rect 15476 11296 15528 11305
rect 15844 11296 15896 11348
rect 16212 11296 16264 11348
rect 16580 11339 16632 11348
rect 16580 11305 16589 11339
rect 16589 11305 16623 11339
rect 16623 11305 16632 11339
rect 16580 11296 16632 11305
rect 17500 11339 17552 11348
rect 17500 11305 17509 11339
rect 17509 11305 17543 11339
rect 17543 11305 17552 11339
rect 17500 11296 17552 11305
rect 19524 11296 19576 11348
rect 19984 11339 20036 11348
rect 19984 11305 19993 11339
rect 19993 11305 20027 11339
rect 20027 11305 20036 11339
rect 19984 11296 20036 11305
rect 20720 11296 20772 11348
rect 22284 11296 22336 11348
rect 23572 11296 23624 11348
rect 23848 11296 23900 11348
rect 25228 11296 25280 11348
rect 25780 11296 25832 11348
rect 12348 11271 12400 11280
rect 12348 11237 12357 11271
rect 12357 11237 12391 11271
rect 12391 11237 12400 11271
rect 12348 11228 12400 11237
rect 12624 11228 12676 11280
rect 14556 11228 14608 11280
rect 17960 11228 18012 11280
rect 19156 11228 19208 11280
rect 11060 11092 11112 11144
rect 11612 11135 11664 11144
rect 10968 11067 11020 11076
rect 10968 11033 10977 11067
rect 10977 11033 11011 11067
rect 11011 11033 11020 11067
rect 10968 11024 11020 11033
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 21732 11228 21784 11280
rect 22192 11228 22244 11280
rect 13084 11160 13136 11212
rect 16396 11160 16448 11212
rect 18788 11160 18840 11212
rect 18880 11160 18932 11212
rect 19524 11160 19576 11212
rect 20352 11160 20404 11212
rect 20904 11160 20956 11212
rect 24032 11203 24084 11212
rect 24032 11169 24041 11203
rect 24041 11169 24075 11203
rect 24075 11169 24084 11203
rect 24032 11160 24084 11169
rect 25136 11160 25188 11212
rect 16120 11135 16172 11144
rect 16120 11101 16129 11135
rect 16129 11101 16163 11135
rect 16163 11101 16172 11135
rect 16120 11092 16172 11101
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 18696 11092 18748 11144
rect 22560 11135 22612 11144
rect 15752 11024 15804 11076
rect 17868 11024 17920 11076
rect 22560 11101 22569 11135
rect 22569 11101 22603 11135
rect 22603 11101 22612 11135
rect 22560 11092 22612 11101
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 23572 11135 23624 11144
rect 22652 11092 22704 11101
rect 23572 11101 23581 11135
rect 23581 11101 23615 11135
rect 23615 11101 23624 11135
rect 23572 11092 23624 11101
rect 23756 11024 23808 11076
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 12440 10956 12492 11008
rect 14740 10956 14792 11008
rect 16948 10999 17000 11008
rect 16948 10965 16957 10999
rect 16957 10965 16991 10999
rect 16991 10965 17000 10999
rect 16948 10956 17000 10965
rect 21916 10956 21968 11008
rect 24216 10956 24268 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 8944 10795 8996 10804
rect 8944 10761 8953 10795
rect 8953 10761 8987 10795
rect 8987 10761 8996 10795
rect 8944 10752 8996 10761
rect 12532 10752 12584 10804
rect 13084 10752 13136 10804
rect 16120 10752 16172 10804
rect 16396 10795 16448 10804
rect 16396 10761 16405 10795
rect 16405 10761 16439 10795
rect 16439 10761 16448 10795
rect 16396 10752 16448 10761
rect 17868 10795 17920 10804
rect 17868 10761 17877 10795
rect 17877 10761 17911 10795
rect 17911 10761 17920 10795
rect 17868 10752 17920 10761
rect 18328 10795 18380 10804
rect 18328 10761 18337 10795
rect 18337 10761 18371 10795
rect 18371 10761 18380 10795
rect 18328 10752 18380 10761
rect 21364 10795 21416 10804
rect 21364 10761 21373 10795
rect 21373 10761 21407 10795
rect 21407 10761 21416 10795
rect 21364 10752 21416 10761
rect 22192 10752 22244 10804
rect 23664 10752 23716 10804
rect 24124 10752 24176 10804
rect 25136 10752 25188 10804
rect 11612 10684 11664 10736
rect 12256 10727 12308 10736
rect 12256 10693 12265 10727
rect 12265 10693 12299 10727
rect 12299 10693 12308 10727
rect 12256 10684 12308 10693
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 8944 10548 8996 10600
rect 10048 10548 10100 10600
rect 10784 10412 10836 10464
rect 10968 10412 11020 10464
rect 11336 10412 11388 10464
rect 23848 10684 23900 10736
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 14740 10591 14792 10600
rect 14740 10557 14774 10591
rect 14774 10557 14792 10591
rect 14740 10548 14792 10557
rect 16120 10548 16172 10600
rect 17592 10548 17644 10600
rect 18604 10548 18656 10600
rect 19432 10548 19484 10600
rect 20352 10548 20404 10600
rect 15752 10480 15804 10532
rect 16672 10480 16724 10532
rect 19064 10480 19116 10532
rect 20444 10480 20496 10532
rect 21732 10591 21784 10600
rect 21732 10557 21741 10591
rect 21741 10557 21775 10591
rect 21775 10557 21784 10591
rect 21732 10548 21784 10557
rect 24124 10591 24176 10600
rect 24124 10557 24158 10591
rect 24158 10557 24176 10591
rect 24124 10548 24176 10557
rect 23756 10480 23808 10532
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 13820 10455 13872 10464
rect 13820 10421 13829 10455
rect 13829 10421 13863 10455
rect 13863 10421 13872 10455
rect 13820 10412 13872 10421
rect 18696 10455 18748 10464
rect 18696 10421 18705 10455
rect 18705 10421 18739 10455
rect 18739 10421 18748 10455
rect 18696 10412 18748 10421
rect 19340 10412 19392 10464
rect 21916 10412 21968 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 11060 10208 11112 10260
rect 12256 10208 12308 10260
rect 12716 10208 12768 10260
rect 13820 10208 13872 10260
rect 17500 10208 17552 10260
rect 18604 10251 18656 10260
rect 18604 10217 18613 10251
rect 18613 10217 18647 10251
rect 18647 10217 18656 10251
rect 18604 10208 18656 10217
rect 19064 10208 19116 10260
rect 19340 10208 19392 10260
rect 19984 10208 20036 10260
rect 20352 10251 20404 10260
rect 20352 10217 20361 10251
rect 20361 10217 20395 10251
rect 20395 10217 20404 10251
rect 20352 10208 20404 10217
rect 22468 10251 22520 10260
rect 22468 10217 22477 10251
rect 22477 10217 22511 10251
rect 22511 10217 22520 10251
rect 22468 10208 22520 10217
rect 23572 10251 23624 10260
rect 23572 10217 23581 10251
rect 23581 10217 23615 10251
rect 23615 10217 23624 10251
rect 23572 10208 23624 10217
rect 24860 10208 24912 10260
rect 14372 10140 14424 10192
rect 17408 10140 17460 10192
rect 24032 10140 24084 10192
rect 11060 10115 11112 10124
rect 11060 10081 11094 10115
rect 11094 10081 11112 10115
rect 11060 10072 11112 10081
rect 11796 10072 11848 10124
rect 12624 10072 12676 10124
rect 13636 10115 13688 10124
rect 13636 10081 13645 10115
rect 13645 10081 13679 10115
rect 13679 10081 13688 10115
rect 13636 10072 13688 10081
rect 9956 10004 10008 10056
rect 13360 10004 13412 10056
rect 16212 10047 16264 10056
rect 13452 9936 13504 9988
rect 16212 10013 16221 10047
rect 16221 10013 16255 10047
rect 16255 10013 16264 10047
rect 16212 10004 16264 10013
rect 15844 9936 15896 9988
rect 17316 10072 17368 10124
rect 19616 10115 19668 10124
rect 19616 10081 19625 10115
rect 19625 10081 19659 10115
rect 19659 10081 19668 10115
rect 19616 10072 19668 10081
rect 21088 10072 21140 10124
rect 23664 10072 23716 10124
rect 17776 10047 17828 10056
rect 17776 10013 17785 10047
rect 17785 10013 17819 10047
rect 17819 10013 17828 10047
rect 17776 10004 17828 10013
rect 19984 10004 20036 10056
rect 21364 10047 21416 10056
rect 21364 10013 21373 10047
rect 21373 10013 21407 10047
rect 21407 10013 21416 10047
rect 21364 10004 21416 10013
rect 21456 10047 21508 10056
rect 21456 10013 21465 10047
rect 21465 10013 21499 10047
rect 21499 10013 21508 10047
rect 21456 10004 21508 10013
rect 23388 10004 23440 10056
rect 23572 10004 23624 10056
rect 24124 10047 24176 10056
rect 24124 10013 24133 10047
rect 24133 10013 24167 10047
rect 24167 10013 24176 10047
rect 24124 10004 24176 10013
rect 14464 9911 14516 9920
rect 14464 9877 14473 9911
rect 14473 9877 14507 9911
rect 14507 9877 14516 9911
rect 14464 9868 14516 9877
rect 15476 9911 15528 9920
rect 15476 9877 15485 9911
rect 15485 9877 15519 9911
rect 15519 9877 15528 9911
rect 15476 9868 15528 9877
rect 16672 9868 16724 9920
rect 19248 9911 19300 9920
rect 19248 9877 19257 9911
rect 19257 9877 19291 9911
rect 19291 9877 19300 9911
rect 19248 9868 19300 9877
rect 21272 9868 21324 9920
rect 22192 9868 22244 9920
rect 22560 9868 22612 9920
rect 23756 9868 23808 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 9956 9707 10008 9716
rect 9956 9673 9965 9707
rect 9965 9673 9999 9707
rect 9999 9673 10008 9707
rect 9956 9664 10008 9673
rect 10048 9664 10100 9716
rect 12900 9664 12952 9716
rect 14372 9707 14424 9716
rect 14372 9673 14381 9707
rect 14381 9673 14415 9707
rect 14415 9673 14424 9707
rect 14372 9664 14424 9673
rect 17316 9707 17368 9716
rect 17316 9673 17325 9707
rect 17325 9673 17359 9707
rect 17359 9673 17368 9707
rect 17316 9664 17368 9673
rect 17408 9664 17460 9716
rect 10876 9596 10928 9648
rect 11796 9639 11848 9648
rect 11796 9605 11805 9639
rect 11805 9605 11839 9639
rect 11839 9605 11848 9639
rect 11796 9596 11848 9605
rect 14004 9596 14056 9648
rect 15936 9596 15988 9648
rect 12716 9528 12768 9580
rect 13452 9571 13504 9580
rect 13452 9537 13461 9571
rect 13461 9537 13495 9571
rect 13495 9537 13504 9571
rect 13452 9528 13504 9537
rect 14464 9528 14516 9580
rect 15660 9528 15712 9580
rect 19616 9664 19668 9716
rect 20168 9664 20220 9716
rect 20352 9664 20404 9716
rect 22008 9639 22060 9648
rect 22008 9605 22017 9639
rect 22017 9605 22051 9639
rect 22051 9605 22060 9639
rect 22008 9596 22060 9605
rect 19340 9571 19392 9580
rect 10784 9460 10836 9512
rect 11244 9503 11296 9512
rect 11244 9469 11253 9503
rect 11253 9469 11287 9503
rect 11287 9469 11296 9503
rect 11244 9460 11296 9469
rect 14740 9503 14792 9512
rect 14740 9469 14749 9503
rect 14749 9469 14783 9503
rect 14783 9469 14792 9503
rect 14740 9460 14792 9469
rect 14832 9460 14884 9512
rect 16212 9460 16264 9512
rect 19340 9537 19349 9571
rect 19349 9537 19383 9571
rect 19383 9537 19392 9571
rect 19340 9528 19392 9537
rect 19432 9571 19484 9580
rect 19432 9537 19441 9571
rect 19441 9537 19475 9571
rect 19475 9537 19484 9571
rect 19432 9528 19484 9537
rect 23112 9596 23164 9648
rect 22468 9528 22520 9580
rect 23756 9571 23808 9580
rect 23756 9537 23765 9571
rect 23765 9537 23799 9571
rect 23799 9537 23808 9571
rect 23756 9528 23808 9537
rect 13176 9435 13228 9444
rect 13176 9401 13185 9435
rect 13185 9401 13219 9435
rect 13219 9401 13228 9435
rect 13176 9392 13228 9401
rect 14372 9392 14424 9444
rect 9680 9324 9732 9376
rect 12164 9324 12216 9376
rect 20076 9392 20128 9444
rect 21364 9435 21416 9444
rect 21364 9401 21373 9435
rect 21373 9401 21407 9435
rect 21407 9401 21416 9435
rect 21364 9392 21416 9401
rect 23664 9460 23716 9512
rect 23572 9392 23624 9444
rect 23940 9392 23992 9444
rect 15936 9367 15988 9376
rect 15936 9333 15945 9367
rect 15945 9333 15979 9367
rect 15979 9333 15988 9367
rect 15936 9324 15988 9333
rect 16028 9324 16080 9376
rect 17776 9324 17828 9376
rect 18328 9367 18380 9376
rect 18328 9333 18337 9367
rect 18337 9333 18371 9367
rect 18371 9333 18380 9367
rect 18328 9324 18380 9333
rect 19984 9324 20036 9376
rect 20812 9367 20864 9376
rect 20812 9333 20821 9367
rect 20821 9333 20855 9367
rect 20855 9333 20864 9367
rect 20812 9324 20864 9333
rect 23020 9367 23072 9376
rect 23020 9333 23029 9367
rect 23029 9333 23063 9367
rect 23063 9333 23072 9367
rect 23020 9324 23072 9333
rect 23664 9324 23716 9376
rect 24124 9324 24176 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 11060 9120 11112 9172
rect 13360 9163 13412 9172
rect 13360 9129 13369 9163
rect 13369 9129 13403 9163
rect 13403 9129 13412 9163
rect 13360 9120 13412 9129
rect 13452 9120 13504 9172
rect 14556 9120 14608 9172
rect 16028 9163 16080 9172
rect 16028 9129 16037 9163
rect 16037 9129 16071 9163
rect 16071 9129 16080 9163
rect 16028 9120 16080 9129
rect 16212 9120 16264 9172
rect 19248 9120 19300 9172
rect 21456 9163 21508 9172
rect 14372 9095 14424 9104
rect 14372 9061 14381 9095
rect 14381 9061 14415 9095
rect 14415 9061 14424 9095
rect 14372 9052 14424 9061
rect 9956 8984 10008 9036
rect 11336 9027 11388 9036
rect 11336 8993 11345 9027
rect 11345 8993 11379 9027
rect 11379 8993 11388 9027
rect 11336 8984 11388 8993
rect 11428 8984 11480 9036
rect 15660 9052 15712 9104
rect 17776 9052 17828 9104
rect 19984 9052 20036 9104
rect 17592 8984 17644 9036
rect 20168 8984 20220 9036
rect 10784 8959 10836 8968
rect 10784 8925 10793 8959
rect 10793 8925 10827 8959
rect 10827 8925 10836 8959
rect 10784 8916 10836 8925
rect 19340 8916 19392 8968
rect 20076 8916 20128 8968
rect 21456 9129 21465 9163
rect 21465 9129 21499 9163
rect 21499 9129 21508 9163
rect 21456 9120 21508 9129
rect 24124 9163 24176 9172
rect 24124 9129 24133 9163
rect 24133 9129 24167 9163
rect 24167 9129 24176 9163
rect 24124 9120 24176 9129
rect 21088 9095 21140 9104
rect 21088 9061 21097 9095
rect 21097 9061 21131 9095
rect 21131 9061 21140 9095
rect 21088 9052 21140 9061
rect 25044 9052 25096 9104
rect 22100 9027 22152 9036
rect 22100 8993 22134 9027
rect 22134 8993 22152 9027
rect 22100 8984 22152 8993
rect 24860 8984 24912 9036
rect 21548 8916 21600 8968
rect 23940 8916 23992 8968
rect 24768 8916 24820 8968
rect 25320 8848 25372 8900
rect 25688 8848 25740 8900
rect 12716 8823 12768 8832
rect 12716 8789 12725 8823
rect 12725 8789 12759 8823
rect 12759 8789 12768 8823
rect 12716 8780 12768 8789
rect 14832 8780 14884 8832
rect 19156 8780 19208 8832
rect 20536 8780 20588 8832
rect 23388 8780 23440 8832
rect 24124 8780 24176 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 11428 8619 11480 8628
rect 11428 8585 11437 8619
rect 11437 8585 11471 8619
rect 11471 8585 11480 8619
rect 11428 8576 11480 8585
rect 14648 8576 14700 8628
rect 17592 8619 17644 8628
rect 17592 8585 17601 8619
rect 17601 8585 17635 8619
rect 17635 8585 17644 8619
rect 17592 8576 17644 8585
rect 11336 8508 11388 8560
rect 14740 8508 14792 8560
rect 18880 8551 18932 8560
rect 15660 8483 15712 8492
rect 15660 8449 15669 8483
rect 15669 8449 15703 8483
rect 15703 8449 15712 8483
rect 15660 8440 15712 8449
rect 16672 8483 16724 8492
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 18880 8517 18889 8551
rect 18889 8517 18923 8551
rect 18923 8517 18932 8551
rect 18880 8508 18932 8517
rect 22100 8576 22152 8628
rect 24768 8508 24820 8560
rect 15936 8372 15988 8424
rect 19248 8415 19300 8424
rect 19248 8381 19257 8415
rect 19257 8381 19291 8415
rect 19291 8381 19300 8415
rect 19248 8372 19300 8381
rect 20168 8372 20220 8424
rect 20536 8372 20588 8424
rect 21548 8372 21600 8424
rect 23296 8372 23348 8424
rect 23756 8372 23808 8424
rect 24860 8372 24912 8424
rect 14832 8304 14884 8356
rect 20076 8304 20128 8356
rect 20812 8304 20864 8356
rect 21640 8304 21692 8356
rect 24216 8304 24268 8356
rect 25688 8347 25740 8356
rect 25688 8313 25697 8347
rect 25697 8313 25731 8347
rect 25731 8313 25740 8347
rect 25688 8304 25740 8313
rect 13544 8236 13596 8288
rect 19248 8236 19300 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 14188 8032 14240 8084
rect 15660 8075 15712 8084
rect 15660 8041 15669 8075
rect 15669 8041 15703 8075
rect 15703 8041 15712 8075
rect 15660 8032 15712 8041
rect 16396 8032 16448 8084
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 18328 8075 18380 8084
rect 18328 8041 18337 8075
rect 18337 8041 18371 8075
rect 18371 8041 18380 8075
rect 18328 8032 18380 8041
rect 19248 8032 19300 8084
rect 21272 8075 21324 8084
rect 21272 8041 21281 8075
rect 21281 8041 21315 8075
rect 21315 8041 21324 8075
rect 21272 8032 21324 8041
rect 25044 8032 25096 8084
rect 1492 7964 1544 8016
rect 9588 7964 9640 8016
rect 11888 7964 11940 8016
rect 13636 7964 13688 8016
rect 15936 7964 15988 8016
rect 24032 7964 24084 8016
rect 17224 7939 17276 7948
rect 17224 7905 17258 7939
rect 17258 7905 17276 7939
rect 17224 7896 17276 7905
rect 23296 7939 23348 7948
rect 13820 7871 13872 7880
rect 13820 7837 13829 7871
rect 13829 7837 13863 7871
rect 13863 7837 13872 7871
rect 13820 7828 13872 7837
rect 13176 7760 13228 7812
rect 16396 7828 16448 7880
rect 16580 7828 16632 7880
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 20076 7828 20128 7880
rect 21640 7828 21692 7880
rect 19340 7803 19392 7812
rect 19340 7769 19349 7803
rect 19349 7769 19383 7803
rect 19383 7769 19392 7803
rect 19340 7760 19392 7769
rect 13360 7735 13412 7744
rect 13360 7701 13369 7735
rect 13369 7701 13403 7735
rect 13403 7701 13412 7735
rect 13360 7692 13412 7701
rect 13544 7692 13596 7744
rect 16488 7692 16540 7744
rect 21456 7692 21508 7744
rect 21548 7692 21600 7744
rect 21916 7692 21968 7744
rect 23296 7905 23305 7939
rect 23305 7905 23339 7939
rect 23339 7905 23348 7939
rect 23296 7896 23348 7905
rect 23388 7896 23440 7948
rect 23572 7939 23624 7948
rect 23572 7905 23606 7939
rect 23606 7905 23624 7939
rect 23572 7896 23624 7905
rect 24860 7896 24912 7948
rect 24216 7692 24268 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 13176 7488 13228 7540
rect 15660 7488 15712 7540
rect 15936 7531 15988 7540
rect 15936 7497 15945 7531
rect 15945 7497 15979 7531
rect 15979 7497 15988 7531
rect 15936 7488 15988 7497
rect 17224 7488 17276 7540
rect 19340 7488 19392 7540
rect 20076 7531 20128 7540
rect 20076 7497 20085 7531
rect 20085 7497 20119 7531
rect 20119 7497 20128 7531
rect 20076 7488 20128 7497
rect 21272 7488 21324 7540
rect 25412 7531 25464 7540
rect 25412 7497 25421 7531
rect 25421 7497 25455 7531
rect 25455 7497 25464 7531
rect 25412 7488 25464 7497
rect 15108 7420 15160 7472
rect 19984 7420 20036 7472
rect 21640 7463 21692 7472
rect 21640 7429 21649 7463
rect 21649 7429 21683 7463
rect 21683 7429 21692 7463
rect 21640 7420 21692 7429
rect 16488 7395 16540 7404
rect 12624 7284 12676 7336
rect 13544 7327 13596 7336
rect 13544 7293 13553 7327
rect 13553 7293 13587 7327
rect 13587 7293 13596 7327
rect 13544 7284 13596 7293
rect 16488 7361 16497 7395
rect 16497 7361 16531 7395
rect 16531 7361 16540 7395
rect 16488 7352 16540 7361
rect 14740 7284 14792 7336
rect 16396 7284 16448 7336
rect 16672 7352 16724 7404
rect 17868 7352 17920 7404
rect 20904 7352 20956 7404
rect 21456 7352 21508 7404
rect 24216 7352 24268 7404
rect 18236 7284 18288 7336
rect 22192 7327 22244 7336
rect 22192 7293 22201 7327
rect 22201 7293 22235 7327
rect 22235 7293 22244 7327
rect 22192 7284 22244 7293
rect 24032 7327 24084 7336
rect 24032 7293 24041 7327
rect 24041 7293 24075 7327
rect 24075 7293 24084 7327
rect 24032 7284 24084 7293
rect 25228 7327 25280 7336
rect 25228 7293 25237 7327
rect 25237 7293 25271 7327
rect 25271 7293 25280 7327
rect 25228 7284 25280 7293
rect 15568 7216 15620 7268
rect 16212 7216 16264 7268
rect 17868 7259 17920 7268
rect 12532 7191 12584 7200
rect 12532 7157 12541 7191
rect 12541 7157 12575 7191
rect 12575 7157 12584 7191
rect 12532 7148 12584 7157
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 14924 7148 14976 7157
rect 17868 7225 17877 7259
rect 17877 7225 17911 7259
rect 17911 7225 17920 7259
rect 17868 7216 17920 7225
rect 19248 7216 19300 7268
rect 16580 7148 16632 7200
rect 19340 7148 19392 7200
rect 23388 7216 23440 7268
rect 20628 7191 20680 7200
rect 20628 7157 20637 7191
rect 20637 7157 20671 7191
rect 20671 7157 20680 7191
rect 20628 7148 20680 7157
rect 22376 7191 22428 7200
rect 22376 7157 22385 7191
rect 22385 7157 22419 7191
rect 22419 7157 22428 7191
rect 22376 7148 22428 7157
rect 23020 7148 23072 7200
rect 23572 7148 23624 7200
rect 24032 7148 24084 7200
rect 25412 7148 25464 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 13176 6987 13228 6996
rect 13176 6953 13185 6987
rect 13185 6953 13219 6987
rect 13219 6953 13228 6987
rect 13176 6944 13228 6953
rect 16212 6987 16264 6996
rect 16212 6953 16221 6987
rect 16221 6953 16255 6987
rect 16255 6953 16264 6987
rect 16212 6944 16264 6953
rect 17776 6944 17828 6996
rect 18420 6944 18472 6996
rect 20904 6944 20956 6996
rect 23296 6944 23348 6996
rect 25136 6987 25188 6996
rect 25136 6953 25145 6987
rect 25145 6953 25179 6987
rect 25179 6953 25188 6987
rect 25136 6944 25188 6953
rect 14924 6876 14976 6928
rect 16396 6876 16448 6928
rect 21272 6919 21324 6928
rect 12072 6851 12124 6860
rect 12072 6817 12106 6851
rect 12106 6817 12124 6851
rect 12072 6808 12124 6817
rect 14188 6851 14240 6860
rect 14188 6817 14197 6851
rect 14197 6817 14231 6851
rect 14231 6817 14240 6851
rect 14188 6808 14240 6817
rect 14832 6808 14884 6860
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 17132 6783 17184 6792
rect 17132 6749 17141 6783
rect 17141 6749 17175 6783
rect 17175 6749 17184 6783
rect 17132 6740 17184 6749
rect 17224 6783 17276 6792
rect 17224 6749 17233 6783
rect 17233 6749 17267 6783
rect 17267 6749 17276 6783
rect 17224 6740 17276 6749
rect 13820 6715 13872 6724
rect 13820 6681 13829 6715
rect 13829 6681 13863 6715
rect 13863 6681 13872 6715
rect 13820 6672 13872 6681
rect 15108 6672 15160 6724
rect 18696 6851 18748 6860
rect 18696 6817 18705 6851
rect 18705 6817 18739 6851
rect 18739 6817 18748 6851
rect 18696 6808 18748 6817
rect 19156 6808 19208 6860
rect 21272 6885 21281 6919
rect 21281 6885 21315 6919
rect 21315 6885 21324 6919
rect 21272 6876 21324 6885
rect 22652 6808 22704 6860
rect 25320 6808 25372 6860
rect 20168 6740 20220 6792
rect 20444 6740 20496 6792
rect 21548 6783 21600 6792
rect 21548 6749 21557 6783
rect 21557 6749 21591 6783
rect 21591 6749 21600 6783
rect 21548 6740 21600 6749
rect 23020 6740 23072 6792
rect 22008 6672 22060 6724
rect 23388 6672 23440 6724
rect 24952 6740 25004 6792
rect 25412 6783 25464 6792
rect 25412 6749 25421 6783
rect 25421 6749 25455 6783
rect 25455 6749 25464 6783
rect 25412 6740 25464 6749
rect 24216 6715 24268 6724
rect 24216 6681 24225 6715
rect 24225 6681 24259 6715
rect 24259 6681 24268 6715
rect 24216 6672 24268 6681
rect 14740 6604 14792 6656
rect 16488 6604 16540 6656
rect 16856 6604 16908 6656
rect 18696 6604 18748 6656
rect 19524 6604 19576 6656
rect 19616 6647 19668 6656
rect 19616 6613 19625 6647
rect 19625 6613 19659 6647
rect 19659 6613 19668 6647
rect 20904 6647 20956 6656
rect 19616 6604 19668 6613
rect 20904 6613 20913 6647
rect 20913 6613 20947 6647
rect 20947 6613 20956 6647
rect 20904 6604 20956 6613
rect 22928 6604 22980 6656
rect 23296 6604 23348 6656
rect 24124 6604 24176 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 12072 6400 12124 6452
rect 17776 6400 17828 6452
rect 21548 6400 21600 6452
rect 22652 6443 22704 6452
rect 22652 6409 22661 6443
rect 22661 6409 22695 6443
rect 22695 6409 22704 6443
rect 22652 6400 22704 6409
rect 23112 6443 23164 6452
rect 23112 6409 23121 6443
rect 23121 6409 23155 6443
rect 23155 6409 23164 6443
rect 23112 6400 23164 6409
rect 23664 6443 23716 6452
rect 23664 6409 23673 6443
rect 23673 6409 23707 6443
rect 23707 6409 23716 6443
rect 23664 6400 23716 6409
rect 24952 6400 25004 6452
rect 19156 6375 19208 6384
rect 19156 6341 19165 6375
rect 19165 6341 19199 6375
rect 19199 6341 19208 6375
rect 19156 6332 19208 6341
rect 23572 6332 23624 6384
rect 17868 6264 17920 6316
rect 18696 6307 18748 6316
rect 18696 6273 18705 6307
rect 18705 6273 18739 6307
rect 18739 6273 18748 6307
rect 18696 6264 18748 6273
rect 24216 6307 24268 6316
rect 24216 6273 24225 6307
rect 24225 6273 24259 6307
rect 24259 6273 24268 6307
rect 24216 6264 24268 6273
rect 11796 6196 11848 6248
rect 12624 6196 12676 6248
rect 16764 6239 16816 6248
rect 13176 6128 13228 6180
rect 16764 6205 16773 6239
rect 16773 6205 16807 6239
rect 16807 6205 16816 6239
rect 16764 6196 16816 6205
rect 18512 6239 18564 6248
rect 18512 6205 18521 6239
rect 18521 6205 18555 6239
rect 18555 6205 18564 6239
rect 18512 6196 18564 6205
rect 19616 6196 19668 6248
rect 20536 6239 20588 6248
rect 20536 6205 20545 6239
rect 20545 6205 20579 6239
rect 20579 6205 20588 6239
rect 20536 6196 20588 6205
rect 23112 6196 23164 6248
rect 24860 6196 24912 6248
rect 16304 6128 16356 6180
rect 14188 6060 14240 6112
rect 15476 6103 15528 6112
rect 15476 6069 15485 6103
rect 15485 6069 15519 6103
rect 15519 6069 15528 6103
rect 15476 6060 15528 6069
rect 15936 6103 15988 6112
rect 15936 6069 15945 6103
rect 15945 6069 15979 6103
rect 15979 6069 15988 6103
rect 15936 6060 15988 6069
rect 16396 6103 16448 6112
rect 16396 6069 16405 6103
rect 16405 6069 16439 6103
rect 16439 6069 16448 6103
rect 16396 6060 16448 6069
rect 16856 6103 16908 6112
rect 16856 6069 16865 6103
rect 16865 6069 16899 6103
rect 16899 6069 16908 6103
rect 16856 6060 16908 6069
rect 17500 6060 17552 6112
rect 19340 6128 19392 6180
rect 21456 6128 21508 6180
rect 23572 6128 23624 6180
rect 25504 6171 25556 6180
rect 25504 6137 25513 6171
rect 25513 6137 25547 6171
rect 25547 6137 25556 6171
rect 25504 6128 25556 6137
rect 17868 6060 17920 6112
rect 19524 6060 19576 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 13360 5856 13412 5908
rect 14832 5856 14884 5908
rect 16856 5856 16908 5908
rect 17132 5856 17184 5908
rect 17868 5856 17920 5908
rect 19248 5856 19300 5908
rect 20444 5856 20496 5908
rect 20812 5856 20864 5908
rect 20904 5856 20956 5908
rect 22008 5856 22060 5908
rect 23020 5899 23072 5908
rect 23020 5865 23029 5899
rect 23029 5865 23063 5899
rect 23063 5865 23072 5899
rect 23020 5856 23072 5865
rect 24216 5856 24268 5908
rect 25136 5899 25188 5908
rect 25136 5865 25145 5899
rect 25145 5865 25179 5899
rect 25179 5865 25188 5899
rect 25136 5856 25188 5865
rect 25412 5899 25464 5908
rect 25412 5865 25421 5899
rect 25421 5865 25455 5899
rect 25455 5865 25464 5899
rect 25412 5856 25464 5865
rect 12532 5788 12584 5840
rect 13820 5788 13872 5840
rect 17224 5788 17276 5840
rect 19064 5788 19116 5840
rect 19524 5788 19576 5840
rect 20536 5788 20588 5840
rect 21916 5831 21968 5840
rect 21916 5797 21925 5831
rect 21925 5797 21959 5831
rect 21959 5797 21968 5831
rect 21916 5788 21968 5797
rect 22836 5788 22888 5840
rect 13176 5720 13228 5772
rect 16028 5763 16080 5772
rect 11336 5695 11388 5704
rect 11336 5661 11345 5695
rect 11345 5661 11379 5695
rect 11379 5661 11388 5695
rect 11336 5652 11388 5661
rect 12440 5652 12492 5704
rect 13636 5652 13688 5704
rect 16028 5729 16062 5763
rect 16062 5729 16080 5763
rect 16028 5720 16080 5729
rect 18236 5763 18288 5772
rect 18236 5729 18245 5763
rect 18245 5729 18279 5763
rect 18279 5729 18288 5763
rect 18236 5720 18288 5729
rect 20720 5720 20772 5772
rect 23572 5788 23624 5840
rect 12624 5584 12676 5636
rect 13084 5516 13136 5568
rect 21364 5652 21416 5704
rect 20536 5584 20588 5636
rect 21548 5584 21600 5636
rect 14740 5516 14792 5568
rect 15936 5516 15988 5568
rect 17224 5516 17276 5568
rect 18512 5516 18564 5568
rect 20904 5559 20956 5568
rect 20904 5525 20913 5559
rect 20913 5525 20947 5559
rect 20947 5525 20956 5559
rect 20904 5516 20956 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 13820 5355 13872 5364
rect 13820 5321 13829 5355
rect 13829 5321 13863 5355
rect 13863 5321 13872 5355
rect 13820 5312 13872 5321
rect 14188 5355 14240 5364
rect 14188 5321 14197 5355
rect 14197 5321 14231 5355
rect 14231 5321 14240 5355
rect 14188 5312 14240 5321
rect 16028 5312 16080 5364
rect 16856 5312 16908 5364
rect 17960 5312 18012 5364
rect 19064 5355 19116 5364
rect 19064 5321 19073 5355
rect 19073 5321 19107 5355
rect 19107 5321 19116 5355
rect 19064 5312 19116 5321
rect 21364 5312 21416 5364
rect 22100 5312 22152 5364
rect 22744 5312 22796 5364
rect 23572 5312 23624 5364
rect 24768 5312 24820 5364
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 13360 5108 13412 5160
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 18420 5151 18472 5160
rect 18420 5117 18429 5151
rect 18429 5117 18463 5151
rect 18463 5117 18472 5151
rect 18420 5108 18472 5117
rect 18696 5219 18748 5228
rect 18696 5185 18705 5219
rect 18705 5185 18739 5219
rect 18739 5185 18748 5219
rect 18696 5176 18748 5185
rect 19524 5108 19576 5160
rect 24032 5176 24084 5228
rect 26884 5244 26936 5296
rect 24676 5219 24728 5228
rect 24676 5185 24685 5219
rect 24685 5185 24719 5219
rect 24719 5185 24728 5219
rect 24676 5176 24728 5185
rect 20536 5108 20588 5160
rect 22744 5108 22796 5160
rect 25228 5151 25280 5160
rect 25228 5117 25237 5151
rect 25237 5117 25271 5151
rect 25271 5117 25280 5151
rect 25228 5108 25280 5117
rect 14740 5040 14792 5092
rect 24124 5040 24176 5092
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 12808 4972 12860 5024
rect 17040 5015 17092 5024
rect 17040 4981 17049 5015
rect 17049 4981 17083 5015
rect 17083 4981 17092 5015
rect 17040 4972 17092 4981
rect 18052 4972 18104 5024
rect 22652 5015 22704 5024
rect 22652 4981 22661 5015
rect 22661 4981 22695 5015
rect 22695 4981 22704 5015
rect 22652 4972 22704 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 12440 4768 12492 4820
rect 12900 4768 12952 4820
rect 13176 4768 13228 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 14004 4768 14056 4820
rect 14372 4768 14424 4820
rect 16396 4811 16448 4820
rect 16396 4777 16405 4811
rect 16405 4777 16439 4811
rect 16439 4777 16448 4811
rect 16396 4768 16448 4777
rect 17776 4768 17828 4820
rect 18052 4811 18104 4820
rect 18052 4777 18061 4811
rect 18061 4777 18095 4811
rect 18095 4777 18104 4811
rect 18052 4768 18104 4777
rect 19248 4811 19300 4820
rect 19248 4777 19257 4811
rect 19257 4777 19291 4811
rect 19291 4777 19300 4811
rect 19248 4768 19300 4777
rect 20536 4768 20588 4820
rect 20720 4811 20772 4820
rect 20720 4777 20729 4811
rect 20729 4777 20763 4811
rect 20763 4777 20772 4811
rect 20720 4768 20772 4777
rect 20812 4768 20864 4820
rect 21088 4768 21140 4820
rect 22560 4768 22612 4820
rect 22836 4811 22888 4820
rect 22836 4777 22845 4811
rect 22845 4777 22879 4811
rect 22879 4777 22888 4811
rect 22836 4768 22888 4777
rect 23572 4768 23624 4820
rect 24216 4768 24268 4820
rect 13268 4700 13320 4752
rect 15844 4700 15896 4752
rect 12164 4632 12216 4684
rect 13820 4632 13872 4684
rect 15384 4632 15436 4684
rect 16028 4632 16080 4684
rect 19984 4632 20036 4684
rect 20812 4632 20864 4684
rect 24124 4700 24176 4752
rect 23296 4675 23348 4684
rect 23296 4641 23305 4675
rect 23305 4641 23339 4675
rect 23339 4641 23348 4675
rect 23296 4632 23348 4641
rect 23388 4632 23440 4684
rect 12716 4607 12768 4616
rect 12716 4573 12725 4607
rect 12725 4573 12759 4607
rect 12759 4573 12768 4607
rect 12716 4564 12768 4573
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 17224 4564 17276 4616
rect 18604 4607 18656 4616
rect 18604 4573 18613 4607
rect 18613 4573 18647 4607
rect 18647 4573 18656 4607
rect 18604 4564 18656 4573
rect 21456 4607 21508 4616
rect 21456 4573 21465 4607
rect 21465 4573 21499 4607
rect 21499 4573 21508 4607
rect 21456 4564 21508 4573
rect 13084 4496 13136 4548
rect 15936 4539 15988 4548
rect 15936 4505 15945 4539
rect 15945 4505 15979 4539
rect 15979 4505 15988 4539
rect 15936 4496 15988 4505
rect 16764 4496 16816 4548
rect 11428 4428 11480 4480
rect 12072 4471 12124 4480
rect 12072 4437 12081 4471
rect 12081 4437 12115 4471
rect 12115 4437 12124 4471
rect 12072 4428 12124 4437
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 15384 4428 15436 4480
rect 19524 4471 19576 4480
rect 19524 4437 19533 4471
rect 19533 4437 19567 4471
rect 19567 4437 19576 4471
rect 19524 4428 19576 4437
rect 20076 4428 20128 4480
rect 22468 4471 22520 4480
rect 22468 4437 22477 4471
rect 22477 4437 22511 4471
rect 22511 4437 22520 4471
rect 22468 4428 22520 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 14280 4224 14332 4276
rect 16028 4267 16080 4276
rect 16028 4233 16037 4267
rect 16037 4233 16071 4267
rect 16071 4233 16080 4267
rect 16028 4224 16080 4233
rect 19984 4224 20036 4276
rect 20812 4224 20864 4276
rect 21088 4224 21140 4276
rect 23480 4224 23532 4276
rect 21640 4156 21692 4208
rect 22284 4156 22336 4208
rect 22468 4156 22520 4208
rect 9128 4088 9180 4140
rect 9680 4088 9732 4140
rect 12072 4088 12124 4140
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 13636 4131 13688 4140
rect 13636 4097 13645 4131
rect 13645 4097 13679 4131
rect 13679 4097 13688 4131
rect 13636 4088 13688 4097
rect 14464 4088 14516 4140
rect 15292 4131 15344 4140
rect 15292 4097 15301 4131
rect 15301 4097 15335 4131
rect 15335 4097 15344 4131
rect 15292 4088 15344 4097
rect 11428 4020 11480 4072
rect 12348 4020 12400 4072
rect 11244 3884 11296 3936
rect 11428 3927 11480 3936
rect 11428 3893 11437 3927
rect 11437 3893 11471 3927
rect 11471 3893 11480 3927
rect 11428 3884 11480 3893
rect 11796 3884 11848 3936
rect 12164 3884 12216 3936
rect 14372 4020 14424 4072
rect 16304 4088 16356 4140
rect 17684 4088 17736 4140
rect 18788 4131 18840 4140
rect 16396 4020 16448 4072
rect 18788 4097 18797 4131
rect 18797 4097 18831 4131
rect 18831 4097 18840 4131
rect 18788 4088 18840 4097
rect 20444 4131 20496 4140
rect 20444 4097 20453 4131
rect 20453 4097 20487 4131
rect 20487 4097 20496 4131
rect 20444 4088 20496 4097
rect 23388 4156 23440 4208
rect 23296 4088 23348 4140
rect 24308 4131 24360 4140
rect 20260 4063 20312 4072
rect 20260 4029 20269 4063
rect 20269 4029 20303 4063
rect 20303 4029 20312 4063
rect 20260 4020 20312 4029
rect 20628 4020 20680 4072
rect 22560 4020 22612 4072
rect 23388 4020 23440 4072
rect 24032 4020 24084 4072
rect 24308 4097 24317 4131
rect 24317 4097 24351 4131
rect 24351 4097 24360 4131
rect 24308 4088 24360 4097
rect 24952 4088 25004 4140
rect 25044 4063 25096 4072
rect 25044 4029 25053 4063
rect 25053 4029 25087 4063
rect 25087 4029 25096 4063
rect 25044 4020 25096 4029
rect 25320 4020 25372 4072
rect 12900 3952 12952 4004
rect 15844 3952 15896 4004
rect 12532 3884 12584 3936
rect 13452 3884 13504 3936
rect 15568 3927 15620 3936
rect 15568 3893 15577 3927
rect 15577 3893 15611 3927
rect 15611 3893 15620 3927
rect 15568 3884 15620 3893
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 18696 3927 18748 3936
rect 18696 3893 18705 3927
rect 18705 3893 18739 3927
rect 18739 3893 18748 3927
rect 18696 3884 18748 3893
rect 20536 3952 20588 4004
rect 19984 3884 20036 3936
rect 22284 3884 22336 3936
rect 24032 3927 24084 3936
rect 24032 3893 24041 3927
rect 24041 3893 24075 3927
rect 24075 3893 24084 3927
rect 24032 3884 24084 3893
rect 24768 3884 24820 3936
rect 25412 3927 25464 3936
rect 25412 3893 25421 3927
rect 25421 3893 25455 3927
rect 25455 3893 25464 3927
rect 25412 3884 25464 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 11152 3723 11204 3732
rect 11152 3689 11161 3723
rect 11161 3689 11195 3723
rect 11195 3689 11204 3723
rect 11152 3680 11204 3689
rect 12072 3680 12124 3732
rect 13084 3680 13136 3732
rect 13452 3723 13504 3732
rect 13452 3689 13461 3723
rect 13461 3689 13495 3723
rect 13495 3689 13504 3723
rect 13452 3680 13504 3689
rect 14004 3723 14056 3732
rect 14004 3689 14013 3723
rect 14013 3689 14047 3723
rect 14047 3689 14056 3723
rect 14004 3680 14056 3689
rect 14372 3723 14424 3732
rect 14372 3689 14381 3723
rect 14381 3689 14415 3723
rect 14415 3689 14424 3723
rect 14372 3680 14424 3689
rect 17224 3723 17276 3732
rect 17224 3689 17233 3723
rect 17233 3689 17267 3723
rect 17267 3689 17276 3723
rect 17224 3680 17276 3689
rect 19340 3680 19392 3732
rect 19984 3680 20036 3732
rect 20260 3723 20312 3732
rect 20260 3689 20269 3723
rect 20269 3689 20303 3723
rect 20303 3689 20312 3723
rect 20260 3680 20312 3689
rect 21456 3680 21508 3732
rect 23296 3723 23348 3732
rect 23296 3689 23305 3723
rect 23305 3689 23339 3723
rect 23339 3689 23348 3723
rect 23296 3680 23348 3689
rect 24216 3680 24268 3732
rect 24952 3680 25004 3732
rect 11244 3612 11296 3664
rect 12256 3612 12308 3664
rect 12716 3612 12768 3664
rect 13544 3612 13596 3664
rect 15292 3612 15344 3664
rect 9956 3544 10008 3596
rect 11520 3544 11572 3596
rect 12624 3544 12676 3596
rect 15384 3544 15436 3596
rect 17500 3544 17552 3596
rect 21916 3544 21968 3596
rect 22744 3544 22796 3596
rect 24124 3587 24176 3596
rect 24124 3553 24147 3587
rect 24147 3553 24176 3587
rect 24124 3544 24176 3553
rect 17776 3519 17828 3528
rect 17776 3485 17785 3519
rect 17785 3485 17819 3519
rect 17819 3485 17828 3519
rect 17776 3476 17828 3485
rect 23296 3476 23348 3528
rect 10048 3451 10100 3460
rect 10048 3417 10057 3451
rect 10057 3417 10091 3451
rect 10091 3417 10100 3451
rect 10048 3408 10100 3417
rect 16764 3408 16816 3460
rect 17500 3408 17552 3460
rect 19892 3408 19944 3460
rect 20720 3408 20772 3460
rect 11980 3383 12032 3392
rect 11980 3349 11989 3383
rect 11989 3349 12023 3383
rect 12023 3349 12032 3383
rect 11980 3340 12032 3349
rect 15292 3340 15344 3392
rect 18052 3340 18104 3392
rect 18788 3340 18840 3392
rect 22744 3383 22796 3392
rect 22744 3349 22753 3383
rect 22753 3349 22787 3383
rect 22787 3349 22796 3383
rect 22744 3340 22796 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 9864 3136 9916 3188
rect 11428 3179 11480 3188
rect 11428 3145 11437 3179
rect 11437 3145 11471 3179
rect 11471 3145 11480 3179
rect 11428 3136 11480 3145
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 12256 3179 12308 3188
rect 12256 3145 12265 3179
rect 12265 3145 12299 3179
rect 12299 3145 12308 3179
rect 12256 3136 12308 3145
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 15660 3136 15712 3188
rect 16304 3136 16356 3188
rect 17500 3179 17552 3188
rect 17500 3145 17509 3179
rect 17509 3145 17543 3179
rect 17543 3145 17552 3179
rect 17500 3136 17552 3145
rect 18972 3136 19024 3188
rect 23572 3136 23624 3188
rect 24124 3136 24176 3188
rect 25044 3136 25096 3188
rect 10324 3111 10376 3120
rect 10324 3077 10333 3111
rect 10333 3077 10367 3111
rect 10367 3077 10376 3111
rect 10324 3068 10376 3077
rect 11520 3068 11572 3120
rect 15292 3068 15344 3120
rect 16120 3068 16172 3120
rect 21364 3068 21416 3120
rect 11888 2932 11940 2984
rect 12624 2932 12676 2984
rect 16764 3043 16816 3052
rect 16764 3009 16773 3043
rect 16773 3009 16807 3043
rect 16807 3009 16816 3043
rect 16764 3000 16816 3009
rect 18236 3000 18288 3052
rect 16488 2932 16540 2984
rect 19524 3000 19576 3052
rect 23848 3043 23900 3052
rect 19248 2932 19300 2984
rect 19892 2975 19944 2984
rect 19892 2941 19901 2975
rect 19901 2941 19935 2975
rect 19935 2941 19944 2975
rect 19892 2932 19944 2941
rect 23848 3009 23857 3043
rect 23857 3009 23891 3043
rect 23891 3009 23900 3043
rect 23848 3000 23900 3009
rect 20720 2932 20772 2984
rect 22928 2975 22980 2984
rect 22928 2941 22937 2975
rect 22937 2941 22971 2975
rect 22971 2941 22980 2975
rect 22928 2932 22980 2941
rect 23572 2932 23624 2984
rect 25136 2932 25188 2984
rect 13176 2907 13228 2916
rect 13176 2873 13185 2907
rect 13185 2873 13219 2907
rect 13219 2873 13228 2907
rect 13176 2864 13228 2873
rect 9956 2839 10008 2848
rect 9956 2805 9965 2839
rect 9965 2805 9999 2839
rect 9999 2805 10008 2839
rect 9956 2796 10008 2805
rect 12716 2839 12768 2848
rect 12716 2805 12725 2839
rect 12725 2805 12759 2839
rect 12759 2805 12768 2839
rect 12716 2796 12768 2805
rect 16672 2864 16724 2916
rect 19432 2864 19484 2916
rect 25228 2907 25280 2916
rect 25228 2873 25237 2907
rect 25237 2873 25271 2907
rect 25271 2873 25280 2907
rect 25228 2864 25280 2873
rect 16304 2796 16356 2848
rect 21916 2839 21968 2848
rect 21916 2805 21925 2839
rect 21925 2805 21959 2839
rect 21959 2805 21968 2839
rect 21916 2796 21968 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 11244 2592 11296 2644
rect 12072 2635 12124 2644
rect 12072 2601 12081 2635
rect 12081 2601 12115 2635
rect 12115 2601 12124 2635
rect 12072 2592 12124 2601
rect 12624 2592 12676 2644
rect 12808 2499 12860 2508
rect 12808 2465 12817 2499
rect 12817 2465 12851 2499
rect 12851 2465 12860 2499
rect 14648 2592 14700 2644
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 19524 2592 19576 2644
rect 20720 2635 20772 2644
rect 20720 2601 20729 2635
rect 20729 2601 20763 2635
rect 20763 2601 20772 2635
rect 20720 2592 20772 2601
rect 22008 2635 22060 2644
rect 22008 2601 22017 2635
rect 22017 2601 22051 2635
rect 22051 2601 22060 2635
rect 22008 2592 22060 2601
rect 24584 2592 24636 2644
rect 24860 2592 24912 2644
rect 19248 2524 19300 2576
rect 12808 2456 12860 2465
rect 15384 2456 15436 2508
rect 12440 2388 12492 2440
rect 14280 2431 14332 2440
rect 14280 2397 14289 2431
rect 14289 2397 14323 2431
rect 14323 2397 14332 2431
rect 14280 2388 14332 2397
rect 16396 2456 16448 2508
rect 17776 2499 17828 2508
rect 17776 2465 17785 2499
rect 17785 2465 17819 2499
rect 17819 2465 17828 2499
rect 17776 2456 17828 2465
rect 18420 2499 18472 2508
rect 18420 2465 18429 2499
rect 18429 2465 18463 2499
rect 18463 2465 18472 2499
rect 18420 2456 18472 2465
rect 20168 2456 20220 2508
rect 16120 2431 16172 2440
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 23756 2456 23808 2508
rect 16120 2388 16172 2397
rect 9220 2363 9272 2372
rect 9220 2329 9229 2363
rect 9229 2329 9263 2363
rect 9263 2329 9272 2363
rect 9220 2320 9272 2329
rect 22744 2388 22796 2440
rect 24492 2388 24544 2440
rect 8760 2295 8812 2304
rect 8760 2261 8769 2295
rect 8769 2261 8803 2295
rect 8803 2261 8812 2295
rect 8760 2252 8812 2261
rect 10968 2252 11020 2304
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 15384 2252 15436 2304
rect 16488 2252 16540 2304
rect 17592 2252 17644 2304
rect 23756 2295 23808 2304
rect 23756 2261 23765 2295
rect 23765 2261 23799 2295
rect 23799 2261 23808 2295
rect 23756 2252 23808 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 21272 552 21324 604
rect 23480 552 23532 604
<< metal2 >>
rect 294 27520 350 28000
rect 938 27520 994 28000
rect 1582 27520 1638 28000
rect 2318 27520 2374 28000
rect 2962 27520 3018 28000
rect 3698 27520 3754 28000
rect 4342 27520 4398 28000
rect 4986 27520 5042 28000
rect 5722 27520 5778 28000
rect 6366 27520 6422 28000
rect 7102 27520 7158 28000
rect 7746 27520 7802 28000
rect 8390 27520 8446 28000
rect 9126 27520 9182 28000
rect 9770 27520 9826 28000
rect 10506 27520 10562 28000
rect 11150 27520 11206 28000
rect 11886 27520 11942 28000
rect 12530 27520 12586 28000
rect 13174 27520 13230 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15290 27520 15346 28000
rect 15934 27520 15990 28000
rect 16578 27520 16634 28000
rect 17314 27520 17370 28000
rect 17958 27520 18014 28000
rect 18694 27520 18750 28000
rect 19338 27520 19394 28000
rect 20074 27520 20130 28000
rect 20718 27520 20774 28000
rect 21362 27520 21418 28000
rect 22098 27520 22154 28000
rect 22742 27520 22798 28000
rect 23110 27704 23166 27713
rect 23110 27639 23166 27648
rect 308 27418 336 27520
rect 308 27390 428 27418
rect 400 12889 428 27390
rect 952 24177 980 27520
rect 938 24168 994 24177
rect 938 24103 994 24112
rect 1596 22681 1624 27520
rect 1582 22672 1638 22681
rect 1582 22607 1638 22616
rect 1582 13968 1638 13977
rect 1582 13903 1638 13912
rect 386 12880 442 12889
rect 386 12815 442 12824
rect 1490 12472 1546 12481
rect 1490 12407 1546 12416
rect 1504 8022 1532 12407
rect 1596 12374 1624 13903
rect 2332 12481 2360 27520
rect 2976 21457 3004 27520
rect 2962 21448 3018 21457
rect 2962 21383 3018 21392
rect 3712 20505 3740 27520
rect 4356 24313 4384 27520
rect 4342 24304 4398 24313
rect 4342 24239 4398 24248
rect 5000 23361 5028 27520
rect 5736 25242 5764 27520
rect 5736 25214 6040 25242
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 4986 23352 5042 23361
rect 4986 23287 5042 23296
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 3698 20496 3754 20505
rect 3698 20431 3754 20440
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6012 17921 6040 25214
rect 6380 24721 6408 27520
rect 6366 24712 6422 24721
rect 6366 24647 6422 24656
rect 7116 20942 7144 27520
rect 7760 22817 7788 27520
rect 7746 22808 7802 22817
rect 7746 22743 7802 22752
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8220 21486 8248 21830
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 8208 21480 8260 21486
rect 8208 21422 8260 21428
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7668 19310 7696 21422
rect 8404 21162 8432 27520
rect 9140 24857 9168 27520
rect 9126 24848 9182 24857
rect 9126 24783 9182 24792
rect 9678 24712 9734 24721
rect 9678 24647 9734 24656
rect 9586 23352 9642 23361
rect 9586 23287 9642 23296
rect 9600 22001 9628 23287
rect 9586 21992 9642 22001
rect 9586 21927 9642 21936
rect 8484 21412 8536 21418
rect 8484 21354 8536 21360
rect 8220 21146 8432 21162
rect 8208 21140 8432 21146
rect 8260 21134 8432 21140
rect 8208 21082 8260 21088
rect 8220 20602 8248 21082
rect 8496 20942 8524 21354
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8484 20936 8536 20942
rect 9692 20913 9720 24647
rect 9784 23633 9812 27520
rect 10520 25786 10548 27520
rect 10520 25758 11008 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 9770 23624 9826 23633
rect 9770 23559 9826 23568
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10692 23180 10744 23186
rect 10692 23122 10744 23128
rect 10048 22976 10100 22982
rect 10048 22918 10100 22924
rect 9864 22500 9916 22506
rect 9864 22442 9916 22448
rect 9876 22234 9904 22442
rect 9864 22228 9916 22234
rect 9864 22170 9916 22176
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9784 21146 9812 22034
rect 9876 21162 9904 22170
rect 10060 21894 10088 22918
rect 10598 22808 10654 22817
rect 10598 22743 10600 22752
rect 10652 22743 10654 22752
rect 10600 22714 10652 22720
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10152 21729 10180 22374
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10704 22234 10732 23122
rect 10782 22944 10838 22953
rect 10782 22879 10838 22888
rect 10796 22778 10824 22879
rect 10874 22808 10930 22817
rect 10784 22772 10836 22778
rect 10874 22743 10930 22752
rect 10784 22714 10836 22720
rect 10692 22228 10744 22234
rect 10692 22170 10744 22176
rect 10232 22092 10284 22098
rect 10232 22034 10284 22040
rect 10138 21720 10194 21729
rect 10138 21655 10194 21664
rect 10140 21480 10192 21486
rect 10244 21468 10272 22034
rect 10192 21440 10272 21468
rect 10140 21422 10192 21428
rect 10152 21350 10180 21422
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 9772 21140 9824 21146
rect 9876 21134 10088 21162
rect 9772 21082 9824 21088
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 8484 20878 8536 20884
rect 9678 20904 9734 20913
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8312 20262 8340 20878
rect 8496 20262 8524 20878
rect 9678 20839 9734 20848
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9692 20466 9720 20742
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9588 20392 9640 20398
rect 9784 20346 9812 20946
rect 9640 20340 9812 20346
rect 9588 20334 9812 20340
rect 9600 20318 9812 20334
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 9036 20256 9088 20262
rect 9036 20198 9088 20204
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7668 18698 7696 19246
rect 7656 18692 7708 18698
rect 7656 18634 7708 18640
rect 5998 17912 6054 17921
rect 5998 17847 6054 17856
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 8312 16017 8340 20198
rect 9048 19514 9076 20198
rect 9036 19508 9088 19514
rect 9036 19450 9088 19456
rect 9600 19417 9628 20318
rect 9876 20058 9904 21014
rect 10060 20890 10088 21134
rect 10152 21078 10180 21286
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10140 21072 10192 21078
rect 10140 21014 10192 21020
rect 10060 20862 10272 20890
rect 9954 20768 10010 20777
rect 9954 20703 10010 20712
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9586 19408 9642 19417
rect 9586 19343 9642 19352
rect 9494 18864 9550 18873
rect 9494 18799 9496 18808
rect 9548 18799 9550 18808
rect 9496 18770 9548 18776
rect 9508 17882 9536 18770
rect 9692 18766 9720 19790
rect 9770 19272 9826 19281
rect 9770 19207 9826 19216
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9692 17542 9720 18702
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 8298 16008 8354 16017
rect 8298 15943 8354 15952
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 9784 14618 9812 19207
rect 9968 18986 9996 20703
rect 10244 20466 10272 20862
rect 10704 20602 10732 21286
rect 10784 20868 10836 20874
rect 10784 20810 10836 20816
rect 10692 20596 10744 20602
rect 10692 20538 10744 20544
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10152 20058 10180 20402
rect 10244 20330 10272 20402
rect 10704 20398 10732 20538
rect 10796 20466 10824 20810
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10232 20324 10284 20330
rect 10232 20266 10284 20272
rect 10888 20210 10916 22743
rect 10980 20641 11008 25758
rect 11164 22574 11192 27520
rect 11334 24576 11390 24585
rect 11334 24511 11390 24520
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 11150 21584 11206 21593
rect 11150 21519 11152 21528
rect 11204 21519 11206 21528
rect 11152 21490 11204 21496
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 11072 21146 11100 21286
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 10966 20632 11022 20641
rect 10966 20567 11022 20576
rect 11256 20534 11284 20946
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 10704 20182 10916 20210
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 10704 19394 10732 20182
rect 10874 20088 10930 20097
rect 10874 20023 10930 20032
rect 10888 19990 10916 20023
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10888 19514 10916 19926
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 9876 18958 9996 18986
rect 10060 19366 10732 19394
rect 9876 17746 9904 18958
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9968 18290 9996 18770
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 9876 13326 9904 14758
rect 9954 13968 10010 13977
rect 9954 13903 10010 13912
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 9692 12986 9720 13262
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9126 12880 9182 12889
rect 9126 12815 9182 12824
rect 2318 12472 2374 12481
rect 2318 12407 2374 12416
rect 1584 12368 1636 12374
rect 1584 12310 1636 12316
rect 1596 11898 1624 12310
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 2056 11558 2084 12242
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 2056 11121 2084 11494
rect 2042 11112 2098 11121
rect 2042 11047 2098 11056
rect 2792 10713 2820 12038
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 9140 11694 9168 12815
rect 9496 12776 9548 12782
rect 9494 12744 9496 12753
rect 9548 12744 9550 12753
rect 9494 12679 9550 12688
rect 9876 12306 9904 13126
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9600 11762 9628 12038
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9128 11688 9180 11694
rect 9600 11665 9628 11698
rect 9128 11630 9180 11636
rect 9586 11656 9642 11665
rect 9140 11354 9168 11630
rect 9586 11591 9642 11600
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9232 11257 9260 11494
rect 9218 11248 9274 11257
rect 9218 11183 9274 11192
rect 8942 11112 8998 11121
rect 8942 11047 8998 11056
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 8956 10810 8984 11047
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 2778 10704 2834 10713
rect 2778 10639 2834 10648
rect 8956 10606 8984 10746
rect 9600 10713 9628 11494
rect 9876 11121 9904 12242
rect 9968 11778 9996 13903
rect 10060 12850 10088 19366
rect 10692 19236 10744 19242
rect 10692 19178 10744 19184
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10152 18329 10180 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10704 18426 10732 19178
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10796 18970 10824 19110
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10138 18320 10194 18329
rect 10138 18255 10194 18264
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10138 17912 10194 17921
rect 10289 17904 10585 17924
rect 10138 17847 10194 17856
rect 10152 17814 10180 17847
rect 10140 17808 10192 17814
rect 10140 17750 10192 17756
rect 10888 17762 10916 19450
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 10980 18698 11008 19314
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 11152 18624 11204 18630
rect 10980 18572 11152 18578
rect 10980 18566 11204 18572
rect 10980 18550 11192 18566
rect 10980 17882 11008 18550
rect 11348 18086 11376 24511
rect 11900 24449 11928 27520
rect 11886 24440 11942 24449
rect 11886 24375 11942 24384
rect 12162 24304 12218 24313
rect 12162 24239 12218 24248
rect 11796 22976 11848 22982
rect 11796 22918 11848 22924
rect 11808 22778 11836 22918
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11888 22568 11940 22574
rect 11888 22510 11940 22516
rect 11520 20936 11572 20942
rect 11518 20904 11520 20913
rect 11572 20904 11574 20913
rect 11518 20839 11574 20848
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 10152 17202 10180 17750
rect 10784 17740 10836 17746
rect 10888 17734 11008 17762
rect 10784 17682 10836 17688
rect 10796 17270 10824 17682
rect 10980 17678 11008 17734
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 11334 17640 11390 17649
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10784 17264 10836 17270
rect 10782 17232 10784 17241
rect 10836 17232 10838 17241
rect 10140 17196 10192 17202
rect 10888 17218 10916 17478
rect 10980 17338 11008 17614
rect 11334 17575 11390 17584
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10888 17190 11008 17218
rect 11348 17202 11376 17575
rect 10782 17167 10838 17176
rect 10140 17138 10192 17144
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10796 16250 10824 16730
rect 10980 16658 11008 17190
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11060 17128 11112 17134
rect 11440 17082 11468 20198
rect 11900 19802 11928 22510
rect 12176 21026 12204 24239
rect 12544 23361 12572 27520
rect 12806 24712 12862 24721
rect 12806 24647 12862 24656
rect 12820 23866 12848 24647
rect 12808 23860 12860 23866
rect 12808 23802 12860 23808
rect 13188 23610 13216 27520
rect 13726 24440 13782 24449
rect 13726 24375 13728 24384
rect 13780 24375 13782 24384
rect 13728 24346 13780 24352
rect 13924 24342 13952 27520
rect 14186 24848 14242 24857
rect 14186 24783 14242 24792
rect 14370 24848 14426 24857
rect 14370 24783 14426 24792
rect 13912 24336 13964 24342
rect 13912 24278 13964 24284
rect 14200 24274 14228 24783
rect 14384 24614 14412 24783
rect 14568 24721 14596 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14554 24712 14610 24721
rect 14554 24647 14610 24656
rect 14372 24608 14424 24614
rect 14372 24550 14424 24556
rect 14556 24608 14608 24614
rect 14556 24550 14608 24556
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14188 24268 14240 24274
rect 14188 24210 14240 24216
rect 13096 23582 13216 23610
rect 13726 23624 13782 23633
rect 13452 23588 13504 23594
rect 12530 23352 12586 23361
rect 12530 23287 12586 23296
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12254 22536 12310 22545
rect 12636 22506 12664 23258
rect 12716 22976 12768 22982
rect 12714 22944 12716 22953
rect 12900 22976 12952 22982
rect 12768 22944 12770 22953
rect 12900 22918 12952 22924
rect 12714 22879 12770 22888
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12728 22574 12756 22714
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12254 22471 12310 22480
rect 12624 22500 12676 22506
rect 12268 22234 12296 22471
rect 12624 22442 12676 22448
rect 12256 22228 12308 22234
rect 12256 22170 12308 22176
rect 12912 22166 12940 22918
rect 12992 22228 13044 22234
rect 12992 22170 13044 22176
rect 12900 22160 12952 22166
rect 12900 22102 12952 22108
rect 12714 21720 12770 21729
rect 12714 21655 12716 21664
rect 12768 21655 12770 21664
rect 12716 21626 12768 21632
rect 12728 21486 12756 21626
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 12624 21344 12676 21350
rect 12624 21286 12676 21292
rect 12176 21010 12296 21026
rect 12176 21004 12308 21010
rect 12176 20998 12256 21004
rect 12256 20946 12308 20952
rect 12268 20262 12296 20946
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12544 20398 12572 20742
rect 12532 20392 12584 20398
rect 12346 20360 12402 20369
rect 12532 20334 12584 20340
rect 12346 20295 12402 20304
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 11900 19774 12020 19802
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11900 18426 11928 19654
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11060 17070 11112 17076
rect 11072 16794 11100 17070
rect 11348 17054 11468 17082
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10876 16176 10928 16182
rect 10876 16118 10928 16124
rect 10888 15910 10916 16118
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10612 14890 10640 15438
rect 10704 15162 10732 15574
rect 10888 15366 10916 15846
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10600 14884 10652 14890
rect 10600 14826 10652 14832
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10060 12442 10088 12650
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10152 12374 10180 13806
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10336 12714 10364 13262
rect 10428 12918 10456 13330
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 10152 11898 10180 12310
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 9968 11750 10180 11778
rect 9956 11620 10008 11626
rect 9956 11562 10008 11568
rect 9968 11354 9996 11562
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9862 11112 9918 11121
rect 9862 11047 9918 11056
rect 9310 10704 9366 10713
rect 9310 10639 9312 10648
rect 9364 10639 9366 10648
rect 9586 10704 9642 10713
rect 9586 10639 9642 10648
rect 9312 10610 9364 10616
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 4986 10160 5042 10169
rect 4986 10095 5042 10104
rect 2318 8936 2374 8945
rect 2318 8871 2374 8880
rect 1492 8016 1544 8022
rect 1492 7958 1544 7964
rect 294 4448 350 4457
rect 294 4383 350 4392
rect 308 480 336 4383
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 952 480 980 4111
rect 1582 2544 1638 2553
rect 1582 2479 1638 2488
rect 1596 480 1624 2479
rect 2332 480 2360 8871
rect 3790 7984 3846 7993
rect 3790 7919 3846 7928
rect 3698 6896 3754 6905
rect 3698 6831 3754 6840
rect 2962 5264 3018 5273
rect 2962 5199 3018 5208
rect 2976 480 3004 5199
rect 3712 4729 3740 6831
rect 3698 4720 3754 4729
rect 3698 4655 3754 4664
rect 3804 4604 3832 7919
rect 4342 7440 4398 7449
rect 4342 7375 4398 7384
rect 3712 4576 3832 4604
rect 3712 480 3740 4576
rect 4356 480 4384 7375
rect 5000 480 5028 10095
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 9968 9722 9996 9998
rect 10060 9722 10088 10542
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 7102 8528 7158 8537
rect 7102 8463 7158 8472
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6366 6760 6422 6769
rect 6366 6695 6422 6704
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5722 1864 5778 1873
rect 5722 1799 5778 1808
rect 5736 480 5764 1799
rect 6380 480 6408 6695
rect 7116 480 7144 8463
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 7746 7848 7802 7857
rect 7746 7783 7802 7792
rect 7760 480 7788 7783
rect 9600 6361 9628 7958
rect 9586 6352 9642 6361
rect 9586 6287 9642 6296
rect 9692 4146 9720 9318
rect 9770 9072 9826 9081
rect 9968 9042 9996 9658
rect 9770 9007 9826 9016
rect 9956 9036 10008 9042
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 8390 3360 8446 3369
rect 8390 3295 8446 3304
rect 8404 480 8432 3295
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8772 1601 8800 2246
rect 8758 1592 8814 1601
rect 8758 1527 8814 1536
rect 9140 480 9168 4082
rect 9218 2408 9274 2417
rect 9218 2343 9220 2352
rect 9272 2343 9274 2352
rect 9220 2314 9272 2320
rect 9784 480 9812 9007
rect 9956 8978 10008 8984
rect 9862 6352 9918 6361
rect 9862 6287 9918 6296
rect 9876 3194 9904 6287
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9968 2854 9996 3538
rect 10046 3496 10102 3505
rect 10046 3431 10048 3440
rect 10100 3431 10102 3440
rect 10048 3402 10100 3408
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9968 2553 9996 2790
rect 9954 2544 10010 2553
rect 10152 2530 10180 11750
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10704 5522 10732 13738
rect 10796 12986 10824 14418
rect 10888 13394 10916 15302
rect 10980 14822 11008 16594
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 11164 16114 11192 16390
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10968 14612 11020 14618
rect 11072 14600 11100 15574
rect 11020 14572 11100 14600
rect 10968 14554 11020 14560
rect 10980 13938 11008 14554
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 11072 13433 11100 14350
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11058 13424 11114 13433
rect 10876 13388 10928 13394
rect 11058 13359 11114 13368
rect 10876 13330 10928 13336
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 11256 12850 11284 14010
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11348 12322 11376 17054
rect 11164 12294 11376 12322
rect 10966 12064 11022 12073
rect 10966 11999 11022 12008
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10796 11354 10824 11494
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10470 10824 10950
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10888 9654 10916 11494
rect 10980 11082 11008 11999
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 10146 11008 10406
rect 11072 10266 11100 11086
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10980 10130 11100 10146
rect 10980 10124 11112 10130
rect 10980 10118 11060 10124
rect 11060 10066 11112 10072
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10796 8974 10824 9454
rect 11072 9178 11100 10066
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10784 8968 10836 8974
rect 10782 8936 10784 8945
rect 10836 8936 10838 8945
rect 10782 8871 10838 8880
rect 11164 7449 11192 12294
rect 11532 12186 11560 18022
rect 11794 17232 11850 17241
rect 11794 17167 11850 17176
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11624 14618 11652 15030
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11624 14074 11652 14418
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11716 13530 11744 13670
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11808 13410 11836 17167
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11900 16289 11928 16594
rect 11886 16280 11942 16289
rect 11886 16215 11888 16224
rect 11940 16215 11942 16224
rect 11888 16186 11940 16192
rect 11256 12158 11560 12186
rect 11256 10282 11284 12158
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11348 10470 11376 11698
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11256 10254 11376 10282
rect 11242 9616 11298 9625
rect 11242 9551 11298 9560
rect 11256 9518 11284 9551
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11348 9330 11376 10254
rect 11256 9302 11376 9330
rect 11150 7440 11206 7449
rect 11150 7375 11206 7384
rect 11164 6610 11192 7375
rect 11256 6769 11284 9302
rect 11440 9042 11468 12038
rect 11532 11937 11560 12158
rect 11716 13382 11836 13410
rect 11518 11928 11574 11937
rect 11518 11863 11574 11872
rect 11716 11234 11744 13382
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11808 12102 11836 12786
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11716 11206 11928 11234
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11624 10742 11652 11086
rect 11702 10976 11758 10985
rect 11702 10911 11758 10920
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11518 9072 11574 9081
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11428 9036 11480 9042
rect 11518 9007 11574 9016
rect 11428 8978 11480 8984
rect 11348 8566 11376 8978
rect 11440 8634 11468 8978
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11242 6760 11298 6769
rect 11242 6695 11298 6704
rect 11164 6582 11284 6610
rect 10704 5494 11100 5522
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 11072 3482 11100 5494
rect 11256 4162 11284 6582
rect 11336 5704 11388 5710
rect 11334 5672 11336 5681
rect 11388 5672 11390 5681
rect 11334 5607 11390 5616
rect 11336 5024 11388 5030
rect 11334 4992 11336 5001
rect 11388 4992 11390 5001
rect 11334 4927 11390 4936
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 11256 4134 11376 4162
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11164 3641 11192 3674
rect 11256 3670 11284 3878
rect 11244 3664 11296 3670
rect 11150 3632 11206 3641
rect 11244 3606 11296 3612
rect 11150 3567 11206 3576
rect 11348 3482 11376 4134
rect 11440 4078 11468 4422
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11428 3936 11480 3942
rect 11426 3904 11428 3913
rect 11480 3904 11482 3913
rect 11426 3839 11482 3848
rect 11426 3768 11482 3777
rect 11426 3703 11482 3712
rect 11072 3454 11192 3482
rect 10324 3120 10376 3126
rect 10322 3088 10324 3097
rect 10376 3088 10378 3097
rect 10322 3023 10378 3032
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10152 2502 10548 2530
rect 9954 2479 10010 2488
rect 10520 480 10548 2502
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 1465 11008 2246
rect 10966 1456 11022 1465
rect 10966 1391 11022 1400
rect 11164 480 11192 3454
rect 11256 3454 11376 3482
rect 11256 2650 11284 3454
rect 11440 3194 11468 3703
rect 11532 3602 11560 9007
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11532 3126 11560 3538
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 11716 2836 11744 10911
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11808 9654 11836 10066
rect 11796 9648 11848 9654
rect 11796 9590 11848 9596
rect 11900 8022 11928 11206
rect 11992 9353 12020 19774
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12070 17912 12126 17921
rect 12070 17847 12072 17856
rect 12124 17847 12126 17856
rect 12072 17818 12124 17824
rect 12176 17542 12204 19110
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12268 18426 12296 18770
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12268 17678 12296 18362
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12176 17202 12204 17478
rect 12268 17338 12296 17614
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12268 16726 12296 17274
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 12070 15736 12126 15745
rect 12070 15671 12126 15680
rect 12084 14346 12112 15671
rect 12360 15552 12388 20295
rect 12544 20233 12572 20334
rect 12530 20224 12586 20233
rect 12530 20159 12586 20168
rect 12636 19961 12664 21286
rect 12820 20482 12848 21354
rect 12912 21146 12940 22102
rect 13004 21418 13032 22170
rect 13096 21554 13124 23582
rect 13726 23559 13782 23568
rect 13452 23530 13504 23536
rect 13268 23180 13320 23186
rect 13268 23122 13320 23128
rect 13280 22234 13308 23122
rect 13358 22672 13414 22681
rect 13358 22607 13414 22616
rect 13268 22228 13320 22234
rect 13268 22170 13320 22176
rect 13268 22092 13320 22098
rect 13268 22034 13320 22040
rect 13280 21690 13308 22034
rect 13268 21684 13320 21690
rect 13268 21626 13320 21632
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 12820 20454 12940 20482
rect 12808 20324 12860 20330
rect 12808 20266 12860 20272
rect 12622 19952 12678 19961
rect 12622 19887 12678 19896
rect 12438 18320 12494 18329
rect 12438 18255 12494 18264
rect 12452 18222 12480 18255
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12452 17882 12480 18158
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 16114 12572 16390
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12544 15706 12572 16050
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12636 15586 12664 19887
rect 12820 19718 12848 20266
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12820 19310 12848 19654
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12728 18290 12756 18702
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12714 18184 12770 18193
rect 12714 18119 12716 18128
rect 12768 18119 12770 18128
rect 12716 18090 12768 18096
rect 12912 17746 12940 20454
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12728 15706 12756 15846
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12268 15524 12388 15552
rect 12544 15558 12664 15586
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 12268 12730 12296 15524
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12360 13530 12388 14486
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12268 12702 12388 12730
rect 12256 12640 12308 12646
rect 12084 12588 12256 12594
rect 12084 12582 12308 12588
rect 12084 12566 12296 12582
rect 11978 9344 12034 9353
rect 11978 9279 12034 9288
rect 11888 8016 11940 8022
rect 11888 7958 11940 7964
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11808 6254 11836 6734
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11900 5556 11928 7958
rect 12084 7018 12112 12566
rect 12360 12458 12388 12702
rect 12176 12430 12388 12458
rect 12176 9382 12204 12430
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12360 11286 12388 12174
rect 12348 11280 12400 11286
rect 12346 11248 12348 11257
rect 12452 11268 12480 12242
rect 12544 11558 12572 15558
rect 12728 15026 12756 15642
rect 12912 15570 12940 16050
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12636 14414 12664 14894
rect 12912 14482 12940 15506
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12636 14074 12664 14350
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12714 12880 12770 12889
rect 12714 12815 12770 12824
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12636 12442 12664 12718
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12636 12073 12664 12378
rect 12622 12064 12678 12073
rect 12622 11999 12678 12008
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12624 11280 12676 11286
rect 12400 11248 12402 11257
rect 12452 11240 12624 11268
rect 12624 11222 12676 11228
rect 12346 11183 12402 11192
rect 12440 11008 12492 11014
rect 12492 10956 12572 10962
rect 12440 10950 12572 10956
rect 12452 10934 12572 10950
rect 12544 10810 12572 10934
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 12268 10266 12296 10678
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12636 10130 12664 11222
rect 12728 10266 12756 12815
rect 12820 12646 12848 13330
rect 13004 12850 13032 21082
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 13096 19990 13124 20742
rect 13188 20058 13216 20878
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 13084 19984 13136 19990
rect 13084 19926 13136 19932
rect 13096 19514 13124 19926
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 13096 16266 13124 17682
rect 13174 17096 13230 17105
rect 13174 17031 13176 17040
rect 13228 17031 13230 17040
rect 13176 17002 13228 17008
rect 13188 16794 13216 17002
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 13280 16590 13308 21490
rect 13372 20942 13400 22607
rect 13464 21146 13492 23530
rect 13544 23520 13596 23526
rect 13544 23462 13596 23468
rect 13556 23322 13584 23462
rect 13544 23316 13596 23322
rect 13544 23258 13596 23264
rect 13544 23112 13596 23118
rect 13740 23089 13768 23559
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 13544 23054 13596 23060
rect 13726 23080 13782 23089
rect 13556 22438 13584 23054
rect 13726 23015 13782 23024
rect 13544 22432 13596 22438
rect 13544 22374 13596 22380
rect 13556 21554 13584 22374
rect 14016 22098 14044 23462
rect 14108 22982 14136 24210
rect 14278 24168 14334 24177
rect 14278 24103 14334 24112
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14108 22817 14136 22918
rect 14094 22808 14150 22817
rect 14094 22743 14150 22752
rect 14004 22092 14056 22098
rect 14004 22034 14056 22040
rect 14016 21690 14044 22034
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13556 21146 13584 21490
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 13740 20346 13768 20878
rect 14002 20496 14058 20505
rect 14002 20431 14058 20440
rect 13820 20392 13872 20398
rect 13648 20340 13820 20346
rect 13648 20334 13872 20340
rect 13648 20318 13860 20334
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13372 19417 13400 19654
rect 13358 19408 13414 19417
rect 13358 19343 13414 19352
rect 13464 18970 13492 19790
rect 13648 19242 13676 20318
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13832 20097 13860 20198
rect 13818 20088 13874 20097
rect 13818 20023 13874 20032
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13464 18426 13492 18906
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13648 17678 13676 19178
rect 13740 18816 13768 19858
rect 13912 19780 13964 19786
rect 13912 19722 13964 19728
rect 13924 19310 13952 19722
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13740 18788 13860 18816
rect 13832 18630 13860 18788
rect 13924 18630 13952 19246
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13832 17921 13860 18566
rect 13818 17912 13874 17921
rect 13818 17847 13874 17856
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13450 16960 13506 16969
rect 13450 16895 13506 16904
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13096 16238 13308 16266
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 13096 15706 13124 15982
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13188 14822 13216 15506
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13096 12730 13124 13670
rect 13188 13297 13216 14758
rect 13280 14385 13308 16238
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13372 15162 13400 15642
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13266 14376 13322 14385
rect 13266 14311 13322 14320
rect 13280 13818 13308 14311
rect 13372 14006 13400 14418
rect 13360 14000 13412 14006
rect 13358 13968 13360 13977
rect 13412 13968 13414 13977
rect 13358 13903 13414 13912
rect 13280 13790 13400 13818
rect 13174 13288 13230 13297
rect 13372 13274 13400 13790
rect 13174 13223 13230 13232
rect 13280 13246 13400 13274
rect 13004 12702 13124 12730
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12898 12608 12954 12617
rect 12898 12543 12954 12552
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12728 9586 12756 10202
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 11992 6990 12112 7018
rect 11992 6905 12020 6990
rect 11978 6896 12034 6905
rect 11978 6831 12034 6840
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12084 6769 12112 6802
rect 12070 6760 12126 6769
rect 12070 6695 12126 6704
rect 12084 6458 12112 6695
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12544 5846 12572 7142
rect 12636 6254 12664 7278
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 11900 5528 12020 5556
rect 11886 5400 11942 5409
rect 11886 5335 11942 5344
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 3369 11836 3878
rect 11794 3360 11850 3369
rect 11794 3295 11850 3304
rect 11900 3194 11928 5335
rect 11992 3618 12020 5528
rect 12452 4826 12480 5646
rect 12636 5642 12664 6190
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12084 4146 12112 4422
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12084 3738 12112 4082
rect 12176 3942 12204 4626
rect 12728 4622 12756 8774
rect 12820 7857 12848 11494
rect 12912 10554 12940 12543
rect 13004 10690 13032 12702
rect 13188 12617 13216 13223
rect 13174 12608 13230 12617
rect 13174 12543 13230 12552
rect 13174 12336 13230 12345
rect 13174 12271 13176 12280
rect 13228 12271 13230 12280
rect 13176 12242 13228 12248
rect 13188 11354 13216 12242
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 13096 10810 13124 11154
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 13004 10662 13124 10690
rect 12912 10526 13032 10554
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12912 9722 12940 10406
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12806 7848 12862 7857
rect 12806 7783 12862 7792
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12728 4434 12756 4558
rect 12452 4406 12756 4434
rect 12452 4298 12480 4406
rect 12268 4270 12480 4298
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 12268 3670 12296 4270
rect 12348 4072 12400 4078
rect 12400 4020 12480 4026
rect 12348 4014 12480 4020
rect 12360 3998 12480 4014
rect 12256 3664 12308 3670
rect 11992 3590 12112 3618
rect 12256 3606 12308 3612
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11900 2990 11928 3130
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11716 2808 11928 2836
rect 11992 2825 12020 3334
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 1873 11652 2246
rect 11610 1864 11666 1873
rect 11610 1799 11666 1808
rect 11900 480 11928 2808
rect 11978 2816 12034 2825
rect 11978 2751 12034 2760
rect 12084 2650 12112 3590
rect 12268 3194 12296 3606
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12452 2446 12480 3998
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12544 480 12572 3878
rect 12714 3768 12770 3777
rect 12714 3703 12770 3712
rect 12728 3670 12756 3703
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12636 2990 12664 3538
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12636 2650 12664 2926
rect 12716 2848 12768 2854
rect 12714 2816 12716 2825
rect 12768 2816 12770 2825
rect 12714 2751 12770 2760
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12820 2514 12848 4966
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12912 4010 12940 4762
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 12898 3768 12954 3777
rect 12898 3703 12954 3712
rect 12912 2689 12940 3703
rect 13004 2836 13032 10526
rect 13096 7721 13124 10662
rect 13174 9480 13230 9489
rect 13174 9415 13176 9424
rect 13228 9415 13230 9424
rect 13176 9386 13228 9392
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13082 7712 13138 7721
rect 13082 7647 13138 7656
rect 13188 7546 13216 7754
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13188 7002 13216 7482
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13188 6186 13216 6938
rect 13176 6180 13228 6186
rect 13176 6122 13228 6128
rect 13188 5778 13216 6122
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 13096 5166 13124 5510
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13188 4826 13216 5714
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13280 4758 13308 13246
rect 13358 12608 13414 12617
rect 13358 12543 13414 12552
rect 13372 12238 13400 12543
rect 13464 12442 13492 16895
rect 13648 16794 13676 17614
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13648 15706 13676 16390
rect 13740 16250 13768 16526
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13740 15609 13768 16186
rect 13820 16040 13872 16046
rect 13924 16028 13952 18566
rect 14016 18358 14044 20431
rect 14292 19825 14320 24103
rect 14370 23352 14426 23361
rect 14370 23287 14426 23296
rect 14278 19816 14334 19825
rect 14278 19751 14334 19760
rect 14384 18850 14412 23287
rect 14464 21888 14516 21894
rect 14464 21830 14516 21836
rect 14476 20806 14504 21830
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14108 18822 14412 18850
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 14016 16658 14044 16730
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 13872 16000 13952 16028
rect 13820 15982 13872 15988
rect 13726 15600 13782 15609
rect 13726 15535 13782 15544
rect 13832 15484 13860 15982
rect 14016 15910 14044 16594
rect 14108 16561 14136 18822
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14200 17882 14228 18022
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14292 17746 14320 18702
rect 14476 18578 14504 18906
rect 14384 18550 14504 18578
rect 14384 17814 14412 18550
rect 14462 18320 14518 18329
rect 14462 18255 14518 18264
rect 14476 18222 14504 18255
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14372 17808 14424 17814
rect 14372 17750 14424 17756
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14280 16992 14332 16998
rect 14384 16980 14412 17750
rect 14332 16952 14412 16980
rect 14280 16934 14332 16940
rect 14200 16590 14228 16934
rect 14188 16584 14240 16590
rect 14094 16552 14150 16561
rect 14188 16526 14240 16532
rect 14094 16487 14150 16496
rect 14200 16289 14228 16526
rect 14186 16280 14242 16289
rect 14186 16215 14242 16224
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 13556 15456 13860 15484
rect 13556 15094 13584 15456
rect 13544 15088 13596 15094
rect 13544 15030 13596 15036
rect 13818 15056 13874 15065
rect 13556 13938 13584 15030
rect 13818 14991 13874 15000
rect 13832 14482 13860 14991
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13924 14618 13952 14758
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 14016 14521 14044 15846
rect 14002 14512 14058 14521
rect 13820 14476 13872 14482
rect 14002 14447 14058 14456
rect 13820 14418 13872 14424
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13820 14272 13872 14278
rect 13740 14232 13820 14260
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13740 12442 13768 14232
rect 13820 14214 13872 14220
rect 13818 13968 13874 13977
rect 13818 13903 13874 13912
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13542 12200 13598 12209
rect 13372 11898 13400 12174
rect 13542 12135 13598 12144
rect 13556 11898 13584 12135
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13832 10554 13860 13903
rect 13924 13802 13952 14350
rect 13912 13796 13964 13802
rect 13912 13738 13964 13744
rect 13924 13530 13952 13738
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13910 11928 13966 11937
rect 13910 11863 13966 11872
rect 13924 11694 13952 11863
rect 14002 11792 14058 11801
rect 14002 11727 14004 11736
rect 14056 11727 14058 11736
rect 14004 11698 14056 11704
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 14004 11620 14056 11626
rect 14004 11562 14056 11568
rect 13832 10526 13952 10554
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 10266 13860 10406
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13358 10160 13414 10169
rect 13358 10095 13414 10104
rect 13636 10124 13688 10130
rect 13372 10062 13400 10095
rect 13636 10066 13688 10072
rect 13360 10056 13412 10062
rect 13648 10033 13676 10066
rect 13360 9998 13412 10004
rect 13634 10024 13690 10033
rect 13372 9178 13400 9998
rect 13452 9988 13504 9994
rect 13634 9959 13690 9968
rect 13452 9930 13504 9936
rect 13464 9586 13492 9930
rect 13924 9625 13952 10526
rect 14016 10441 14044 11562
rect 14002 10432 14058 10441
rect 14002 10367 14058 10376
rect 14002 10024 14058 10033
rect 14002 9959 14058 9968
rect 14016 9654 14044 9959
rect 14004 9648 14056 9654
rect 13910 9616 13966 9625
rect 13452 9580 13504 9586
rect 14004 9590 14056 9596
rect 13910 9551 13966 9560
rect 13452 9522 13504 9528
rect 13464 9178 13492 9522
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13450 7984 13506 7993
rect 13450 7919 13506 7928
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13372 5914 13400 7686
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13372 5166 13400 5850
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13268 4752 13320 4758
rect 13268 4694 13320 4700
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 13096 4146 13124 4490
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13096 3738 13124 4082
rect 13280 3777 13308 4694
rect 13464 3942 13492 7919
rect 13556 7750 13584 8230
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13648 7857 13676 7958
rect 13820 7880 13872 7886
rect 13634 7848 13690 7857
rect 13820 7822 13872 7828
rect 13634 7783 13690 7792
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13556 7342 13584 7686
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13832 6730 13860 7822
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13648 4826 13676 5646
rect 13832 5370 13860 5782
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13818 5128 13874 5137
rect 13818 5063 13874 5072
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13832 4690 13860 5063
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 13820 4684 13872 4690
rect 13648 4644 13820 4672
rect 13648 4593 13676 4644
rect 13820 4626 13872 4632
rect 13634 4584 13690 4593
rect 13634 4519 13690 4528
rect 13648 4146 13676 4519
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13266 3768 13322 3777
rect 13084 3732 13136 3738
rect 13542 3768 13598 3777
rect 13266 3703 13322 3712
rect 13452 3732 13504 3738
rect 13084 3674 13136 3680
rect 14016 3738 14044 4762
rect 13542 3703 13598 3712
rect 14004 3732 14056 3738
rect 13452 3674 13504 3680
rect 13464 3194 13492 3674
rect 13556 3670 13584 3703
rect 14004 3674 14056 3680
rect 13544 3664 13596 3670
rect 14108 3618 14136 15914
rect 14200 15706 14228 16215
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14188 14612 14240 14618
rect 14292 14600 14320 16934
rect 14476 16538 14504 18022
rect 14568 16697 14596 24550
rect 15304 24426 15332 27520
rect 15948 24857 15976 27520
rect 16304 25356 16356 25362
rect 16304 25298 16356 25304
rect 15934 24848 15990 24857
rect 15934 24783 15990 24792
rect 16316 24614 16344 25298
rect 16592 24698 16620 27520
rect 17328 25498 17356 27520
rect 17316 25492 17368 25498
rect 17316 25434 17368 25440
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 16500 24682 16620 24698
rect 16856 24744 16908 24750
rect 16856 24686 16908 24692
rect 16488 24676 16620 24682
rect 16540 24670 16620 24676
rect 16488 24618 16540 24624
rect 16304 24608 16356 24614
rect 16304 24550 16356 24556
rect 15120 24410 15332 24426
rect 15108 24404 15332 24410
rect 15160 24398 15332 24404
rect 15108 24346 15160 24352
rect 15752 24268 15804 24274
rect 15752 24210 15804 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15764 23866 15792 24210
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15290 23352 15346 23361
rect 14648 23316 14700 23322
rect 15290 23287 15346 23296
rect 14648 23258 14700 23264
rect 14660 23118 14688 23258
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 14660 22642 14688 23054
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14660 21894 14688 22578
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14844 22098 14872 22374
rect 14832 22092 14884 22098
rect 14832 22034 14884 22040
rect 14738 21992 14794 22001
rect 14738 21927 14794 21936
rect 14752 21894 14780 21927
rect 14648 21888 14700 21894
rect 14648 21830 14700 21836
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14752 21486 14780 21830
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14740 21480 14792 21486
rect 14646 21448 14702 21457
rect 14740 21422 14792 21428
rect 14646 21383 14648 21392
rect 14700 21383 14702 21392
rect 14648 21354 14700 21360
rect 14752 21298 14780 21422
rect 14660 21270 14780 21298
rect 14832 21344 14884 21350
rect 14832 21286 14884 21292
rect 14554 16688 14610 16697
rect 14554 16623 14610 16632
rect 14476 16510 14596 16538
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14476 16046 14504 16390
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14476 15706 14504 15982
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 14384 15026 14412 15370
rect 14476 15026 14504 15642
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 14240 14572 14320 14600
rect 14188 14554 14240 14560
rect 14200 13734 14228 14554
rect 14384 14346 14412 14962
rect 14372 14340 14424 14346
rect 14372 14282 14424 14288
rect 14476 14074 14504 14962
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14568 13954 14596 16510
rect 14292 13926 14596 13954
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14200 11626 14228 12174
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14186 11384 14242 11393
rect 14186 11319 14242 11328
rect 14200 8242 14228 11319
rect 14292 9432 14320 13926
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14384 11558 14412 12242
rect 14476 12238 14504 12922
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14384 11393 14412 11494
rect 14370 11384 14426 11393
rect 14476 11354 14504 12174
rect 14568 11830 14596 12718
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14370 11319 14426 11328
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14568 11286 14596 11766
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14464 10600 14516 10606
rect 14568 10588 14596 11222
rect 14516 10560 14596 10588
rect 14464 10542 14516 10548
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 14384 9722 14412 10134
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14476 9586 14504 9862
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14372 9444 14424 9450
rect 14292 9404 14372 9432
rect 14372 9386 14424 9392
rect 14384 9110 14412 9386
rect 14568 9178 14596 10560
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14372 9104 14424 9110
rect 14370 9072 14372 9081
rect 14424 9072 14426 9081
rect 14370 9007 14426 9016
rect 14660 8786 14688 21270
rect 14844 21146 14872 21286
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 14752 19700 14780 20946
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14844 20584 14872 20742
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14844 20556 14964 20584
rect 14936 20398 14964 20556
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 14936 19786 14964 20334
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 14832 19712 14884 19718
rect 14752 19672 14832 19700
rect 14832 19654 14884 19660
rect 14738 19408 14794 19417
rect 14738 19343 14794 19352
rect 14752 17882 14780 19343
rect 14844 19281 14872 19654
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14830 19272 14886 19281
rect 14830 19207 14886 19216
rect 14844 18873 14872 19207
rect 15304 18970 15332 23287
rect 15396 23186 15424 23462
rect 15384 23180 15436 23186
rect 15384 23122 15436 23128
rect 15568 22024 15620 22030
rect 15566 21992 15568 22001
rect 15620 21992 15622 22001
rect 15476 21956 15528 21962
rect 15566 21927 15622 21936
rect 15476 21898 15528 21904
rect 15488 21078 15516 21898
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15658 20496 15714 20505
rect 15658 20431 15714 20440
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15396 19514 15424 19858
rect 15474 19816 15530 19825
rect 15474 19751 15530 19760
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 14830 18864 14886 18873
rect 14830 18799 14886 18808
rect 15290 18728 15346 18737
rect 15290 18663 15292 18672
rect 15344 18663 15346 18672
rect 15292 18634 15344 18640
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14844 18426 14872 18566
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15488 18426 15516 19751
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15384 18080 15436 18086
rect 14830 18048 14886 18057
rect 15384 18022 15436 18028
rect 14830 17983 14886 17992
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14752 17338 14780 17682
rect 14844 17678 14872 17983
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 15304 16794 15332 17682
rect 15396 17202 15424 18022
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 15026 15332 16730
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15488 15745 15516 16594
rect 15672 16130 15700 20431
rect 15764 19514 15792 23802
rect 16040 23186 16068 24142
rect 16028 23180 16080 23186
rect 16028 23122 16080 23128
rect 15934 22808 15990 22817
rect 15934 22743 15990 22752
rect 15844 20324 15896 20330
rect 15844 20266 15896 20272
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 15750 19408 15806 19417
rect 15750 19343 15806 19352
rect 15764 18970 15792 19343
rect 15752 18964 15804 18970
rect 15752 18906 15804 18912
rect 15856 18766 15884 20266
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15856 18426 15884 18702
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15844 18148 15896 18154
rect 15844 18090 15896 18096
rect 15856 17746 15884 18090
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 15752 17536 15804 17542
rect 15856 17524 15884 17682
rect 15804 17496 15884 17524
rect 15752 17478 15804 17484
rect 15856 16998 15884 17496
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15856 16658 15884 16934
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15672 16102 15792 16130
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15474 15736 15530 15745
rect 15474 15671 15530 15680
rect 15474 15600 15530 15609
rect 15474 15535 15530 15544
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15304 13530 15332 14282
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 14844 13326 14872 13466
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14844 12986 14872 13262
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15212 12322 15240 12854
rect 15290 12744 15346 12753
rect 15290 12679 15346 12688
rect 15304 12442 15332 12679
rect 15396 12481 15424 15098
rect 15488 12850 15516 15535
rect 15580 14890 15608 15846
rect 15764 15450 15792 16102
rect 15856 15706 15884 16594
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15764 15422 15884 15450
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15568 14884 15620 14890
rect 15568 14826 15620 14832
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15382 12472 15438 12481
rect 15292 12436 15344 12442
rect 15488 12442 15516 12650
rect 15382 12407 15438 12416
rect 15476 12436 15528 12442
rect 15292 12378 15344 12384
rect 15476 12378 15528 12384
rect 15212 12294 15332 12322
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14738 11112 14794 11121
rect 14738 11047 14794 11056
rect 14752 11014 14780 11047
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14752 10606 14780 10950
rect 14740 10600 14792 10606
rect 14844 10577 14872 11698
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 11354 15148 11494
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14740 10542 14792 10548
rect 14830 10568 14886 10577
rect 14830 10503 14886 10512
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14738 9616 14794 9625
rect 14738 9551 14794 9560
rect 14752 9518 14780 9551
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14844 8838 14872 9454
rect 14568 8758 14688 8786
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14200 8214 14412 8242
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14200 6866 14228 8026
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14278 6760 14334 6769
rect 14278 6695 14334 6704
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14200 5370 14228 6054
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14292 4622 14320 6695
rect 14384 4826 14412 8214
rect 14462 6896 14518 6905
rect 14462 6831 14518 6840
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14292 4282 14320 4558
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14476 4146 14504 6831
rect 14568 5409 14596 8758
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14554 5400 14610 5409
rect 14554 5335 14610 5344
rect 14568 4865 14596 5335
rect 14554 4856 14610 4865
rect 14554 4791 14610 4800
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14384 3738 14412 4014
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 13544 3606 13596 3612
rect 14016 3590 14136 3618
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13174 2952 13230 2961
rect 13174 2887 13176 2896
rect 13228 2887 13230 2896
rect 13176 2858 13228 2864
rect 13004 2808 13124 2836
rect 12898 2680 12954 2689
rect 13096 2666 13124 2808
rect 14016 2666 14044 3590
rect 13096 2638 13216 2666
rect 12898 2615 12954 2624
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 13188 480 13216 2638
rect 13924 2638 14044 2666
rect 14660 2650 14688 8570
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 14752 7342 14780 8502
rect 14844 8362 14872 8774
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 14936 6934 14964 7142
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14752 5574 14780 6598
rect 14844 6225 14872 6802
rect 14936 6769 14964 6870
rect 14922 6760 14978 6769
rect 15120 6730 15148 7414
rect 14922 6695 14978 6704
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14830 6216 14886 6225
rect 14830 6151 14886 6160
rect 14844 5914 14872 6151
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14752 5098 14780 5510
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14752 4486 14780 5034
rect 15304 4593 15332 12294
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15396 11694 15424 12038
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15488 11354 15516 12242
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15382 10432 15438 10441
rect 15382 10367 15438 10376
rect 15396 9761 15424 10367
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15382 9752 15438 9761
rect 15382 9687 15438 9696
rect 15382 9344 15438 9353
rect 15382 9279 15438 9288
rect 15396 4690 15424 9279
rect 15488 9217 15516 9862
rect 15474 9208 15530 9217
rect 15474 9143 15530 9152
rect 15580 7274 15608 14554
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15672 12646 15700 13330
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15672 9897 15700 12582
rect 15764 12345 15792 15302
rect 15856 14618 15884 15422
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 14074 15884 14350
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15856 12374 15884 13806
rect 15948 12617 15976 22743
rect 16040 22234 16068 23122
rect 16118 22944 16174 22953
rect 16118 22879 16174 22888
rect 16028 22228 16080 22234
rect 16028 22170 16080 22176
rect 16132 22114 16160 22879
rect 16040 22086 16160 22114
rect 16040 17649 16068 22086
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16120 19236 16172 19242
rect 16120 19178 16172 19184
rect 16132 18630 16160 19178
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16026 17640 16082 17649
rect 16026 17575 16082 17584
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 16040 16590 16068 17478
rect 16132 16726 16160 18566
rect 16120 16720 16172 16726
rect 16120 16662 16172 16668
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 16040 15910 16068 16526
rect 16132 16046 16160 16662
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 16040 15638 16068 15846
rect 16028 15632 16080 15638
rect 16028 15574 16080 15580
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16040 12986 16068 13330
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16040 12889 16068 12922
rect 16026 12880 16082 12889
rect 16026 12815 16082 12824
rect 16132 12764 16160 15982
rect 16224 12918 16252 19450
rect 16316 15881 16344 24550
rect 16396 24336 16448 24342
rect 16396 24278 16448 24284
rect 16408 23866 16436 24278
rect 16488 24064 16540 24070
rect 16488 24006 16540 24012
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 16500 22794 16528 24006
rect 16684 23662 16712 24006
rect 16868 23730 16896 24686
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16672 23656 16724 23662
rect 16672 23598 16724 23604
rect 16500 22778 16620 22794
rect 16500 22772 16632 22778
rect 16500 22766 16580 22772
rect 16580 22714 16632 22720
rect 16592 22234 16620 22714
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16948 21888 17000 21894
rect 16948 21830 17000 21836
rect 16960 21554 16988 21830
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 16408 21010 16436 21422
rect 16488 21344 16540 21350
rect 16488 21286 16540 21292
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 16408 20262 16436 20946
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16500 20074 16528 21286
rect 16672 20324 16724 20330
rect 16672 20266 16724 20272
rect 16500 20046 16620 20074
rect 16684 20058 16712 20266
rect 16776 20058 16804 21286
rect 16868 21146 16896 21286
rect 16960 21146 16988 21490
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 17052 20482 17080 24754
rect 17972 24614 18000 27520
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17408 24064 17460 24070
rect 17408 24006 17460 24012
rect 17592 24064 17644 24070
rect 17592 24006 17644 24012
rect 17132 23860 17184 23866
rect 17132 23802 17184 23808
rect 16960 20454 17080 20482
rect 16592 19990 16620 20046
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16776 19514 16804 19994
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16762 19272 16818 19281
rect 16762 19207 16818 19216
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16408 17542 16436 19110
rect 16776 18834 16804 19207
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16580 18216 16632 18222
rect 16500 18176 16580 18204
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16500 17338 16528 18176
rect 16580 18158 16632 18164
rect 16684 17814 16712 18634
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 16776 17610 16804 18770
rect 16960 18290 16988 20454
rect 17144 20369 17172 23802
rect 17420 22982 17448 24006
rect 17500 23656 17552 23662
rect 17500 23598 17552 23604
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17316 22092 17368 22098
rect 17316 22034 17368 22040
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17130 20360 17186 20369
rect 17040 20324 17092 20330
rect 17130 20295 17186 20304
rect 17040 20266 17092 20272
rect 17052 19378 17080 20266
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 17236 19258 17264 21354
rect 17328 21350 17356 22034
rect 17420 22030 17448 22918
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17420 21690 17448 21966
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17328 19310 17356 21286
rect 17408 21140 17460 21146
rect 17408 21082 17460 21088
rect 17420 20602 17448 21082
rect 17408 20596 17460 20602
rect 17408 20538 17460 20544
rect 17420 19514 17448 20538
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17052 19230 17264 19258
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16764 17604 16816 17610
rect 16764 17546 16816 17552
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16408 16794 16436 16934
rect 16396 16788 16448 16794
rect 16396 16730 16448 16736
rect 16394 16688 16450 16697
rect 16394 16623 16450 16632
rect 16302 15872 16358 15881
rect 16302 15807 16358 15816
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16316 14278 16344 15438
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16040 12736 16160 12764
rect 15934 12608 15990 12617
rect 15934 12543 15990 12552
rect 15934 12472 15990 12481
rect 15934 12407 15990 12416
rect 15844 12368 15896 12374
rect 15750 12336 15806 12345
rect 15844 12310 15896 12316
rect 15750 12271 15806 12280
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15764 11082 15792 12174
rect 15856 11558 15884 12174
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 15658 9888 15714 9897
rect 15658 9823 15714 9832
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15672 9110 15700 9522
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15672 8498 15700 9046
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15672 7546 15700 8026
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15290 4584 15346 4593
rect 15290 4519 15346 4528
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15304 4146 15332 4519
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15292 3664 15344 3670
rect 15292 3606 15344 3612
rect 15304 3398 15332 3606
rect 15396 3602 15424 4422
rect 15488 4049 15516 6054
rect 15566 4312 15622 4321
rect 15566 4247 15622 4256
rect 15474 4040 15530 4049
rect 15474 3975 15530 3984
rect 15580 3942 15608 4247
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15474 3496 15530 3505
rect 15474 3431 15530 3440
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15304 3126 15332 3334
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 14648 2644 14700 2650
rect 13924 480 13952 2638
rect 14648 2586 14700 2592
rect 14278 2544 14334 2553
rect 14278 2479 14334 2488
rect 15384 2508 15436 2514
rect 14292 2446 14320 2479
rect 15384 2450 15436 2456
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 15396 2310 15424 2450
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15396 1737 15424 2246
rect 15382 1728 15438 1737
rect 15382 1663 15438 1672
rect 14554 1592 14610 1601
rect 14554 1527 14610 1536
rect 14568 480 14596 1527
rect 15488 626 15516 3431
rect 15672 3194 15700 6734
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15764 1057 15792 10474
rect 15856 9994 15884 11290
rect 15844 9988 15896 9994
rect 15844 9930 15896 9936
rect 15842 9888 15898 9897
rect 15842 9823 15898 9832
rect 15856 8242 15884 9823
rect 15948 9654 15976 12407
rect 15936 9648 15988 9654
rect 15936 9590 15988 9596
rect 16040 9466 16068 12736
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16132 11830 16160 12582
rect 16210 12336 16266 12345
rect 16210 12271 16266 12280
rect 16120 11824 16172 11830
rect 16120 11766 16172 11772
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16132 11150 16160 11630
rect 16224 11354 16252 12271
rect 16316 11665 16344 14214
rect 16408 14074 16436 16623
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16776 15994 16804 17546
rect 16960 16726 16988 18022
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 16854 16552 16910 16561
rect 16854 16487 16910 16496
rect 16868 16114 16896 16487
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16684 15745 16712 15982
rect 16776 15966 16896 15994
rect 16670 15736 16726 15745
rect 16670 15671 16726 15680
rect 16672 15632 16724 15638
rect 16672 15574 16724 15580
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16500 15473 16528 15506
rect 16486 15464 16542 15473
rect 16486 15399 16542 15408
rect 16500 15162 16528 15399
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16486 14784 16542 14793
rect 16486 14719 16542 14728
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16408 12889 16436 13126
rect 16394 12880 16450 12889
rect 16394 12815 16450 12824
rect 16396 12776 16448 12782
rect 16394 12744 16396 12753
rect 16448 12744 16450 12753
rect 16394 12679 16450 12688
rect 16500 12594 16528 14719
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16592 13190 16620 13806
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16408 12566 16528 12594
rect 16302 11656 16358 11665
rect 16302 11591 16358 11600
rect 16212 11348 16264 11354
rect 16408 11336 16436 12566
rect 16488 12436 16540 12442
rect 16592 12424 16620 12786
rect 16540 12396 16620 12424
rect 16488 12378 16540 12384
rect 16592 12345 16620 12396
rect 16578 12336 16634 12345
rect 16578 12271 16634 12280
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 16212 11290 16264 11296
rect 16316 11308 16436 11336
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16132 10810 16160 11086
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16132 10606 16160 10746
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16316 10305 16344 11308
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16408 10810 16436 11154
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16302 10296 16358 10305
rect 16302 10231 16358 10240
rect 16500 10146 16528 11766
rect 16592 11354 16620 12038
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16684 10538 16712 15574
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16776 15026 16804 15438
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16776 14618 16804 14962
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16776 13462 16804 14554
rect 16764 13456 16816 13462
rect 16764 13398 16816 13404
rect 16776 12986 16804 13398
rect 16868 13190 16896 15966
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16960 14618 16988 14894
rect 17052 14793 17080 19230
rect 17512 19156 17540 23598
rect 17604 23254 17632 24006
rect 17696 23866 17724 24210
rect 17684 23860 17736 23866
rect 17684 23802 17736 23808
rect 17592 23248 17644 23254
rect 17592 23190 17644 23196
rect 17604 22778 17632 23190
rect 17592 22772 17644 22778
rect 17592 22714 17644 22720
rect 17682 20224 17738 20233
rect 17682 20159 17738 20168
rect 17696 19854 17724 20159
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17696 19310 17724 19790
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17328 19128 17540 19156
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17144 17542 17172 17682
rect 17236 17649 17264 18566
rect 17222 17640 17278 17649
rect 17222 17575 17278 17584
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17144 17202 17172 17478
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17038 14784 17094 14793
rect 17038 14719 17094 14728
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 17328 14414 17356 19128
rect 17788 18952 17816 24550
rect 17958 24440 18014 24449
rect 18708 24410 18736 27520
rect 18972 25356 19024 25362
rect 18972 25298 19024 25304
rect 18984 24614 19012 25298
rect 19352 25242 19380 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19352 25214 19564 25242
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19248 24744 19300 24750
rect 19444 24698 19472 25094
rect 19300 24692 19472 24698
rect 19248 24686 19472 24692
rect 19260 24670 19472 24686
rect 18972 24608 19024 24614
rect 18972 24550 19024 24556
rect 17958 24375 17960 24384
rect 18012 24375 18014 24384
rect 18696 24404 18748 24410
rect 17960 24346 18012 24352
rect 18696 24346 18748 24352
rect 17972 23474 18000 24346
rect 18984 24177 19012 24550
rect 19156 24268 19208 24274
rect 19156 24210 19208 24216
rect 18970 24168 19026 24177
rect 18328 24132 18380 24138
rect 18970 24103 19026 24112
rect 18328 24074 18380 24080
rect 18340 23662 18368 24074
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 17880 23446 18000 23474
rect 17880 23322 17908 23446
rect 18064 23322 18092 23598
rect 19168 23594 19196 24210
rect 19156 23588 19208 23594
rect 19156 23530 19208 23536
rect 19168 23361 19196 23530
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19154 23352 19210 23361
rect 17868 23316 17920 23322
rect 17868 23258 17920 23264
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 19064 23316 19116 23322
rect 19154 23287 19210 23296
rect 19064 23258 19116 23264
rect 18420 23112 18472 23118
rect 18420 23054 18472 23060
rect 18432 22778 18460 23054
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 18420 22772 18472 22778
rect 18420 22714 18472 22720
rect 17880 21962 17908 22714
rect 19076 22574 19104 23258
rect 19352 23118 19380 23462
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19352 22574 19380 23054
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 17868 21956 17920 21962
rect 17868 21898 17920 21904
rect 18064 21486 18092 22374
rect 18512 21956 18564 21962
rect 18512 21898 18564 21904
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 18156 21554 18184 21830
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 18064 21146 18092 21422
rect 18524 21418 18552 21898
rect 19076 21894 19104 22510
rect 19064 21888 19116 21894
rect 19064 21830 19116 21836
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19076 21486 19104 21830
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 18512 21412 18564 21418
rect 18512 21354 18564 21360
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18052 21140 18104 21146
rect 18052 21082 18104 21088
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17972 20584 18000 20946
rect 17880 20556 18000 20584
rect 17880 20262 17908 20556
rect 18156 20482 18184 21082
rect 18064 20454 18276 20482
rect 18064 20398 18092 20454
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17880 19700 17908 20198
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 17880 19672 18000 19700
rect 17512 18924 17816 18952
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17420 15570 17448 18226
rect 17512 16590 17540 18924
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 17604 18068 17632 18770
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17696 18222 17724 18702
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 17684 18080 17736 18086
rect 17604 18040 17684 18068
rect 17684 18022 17736 18028
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17512 16250 17540 16526
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17420 14822 17448 15506
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17420 13977 17448 14758
rect 17406 13968 17462 13977
rect 17406 13903 17462 13912
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16776 12209 16804 12582
rect 16762 12200 16818 12209
rect 16762 12135 16818 12144
rect 16868 11694 16896 13126
rect 16960 11830 16988 13330
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16946 11112 17002 11121
rect 16946 11047 17002 11056
rect 16960 11014 16988 11047
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16672 10532 16724 10538
rect 16672 10474 16724 10480
rect 16316 10118 16528 10146
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16224 9518 16252 9998
rect 16212 9512 16264 9518
rect 16040 9438 16160 9466
rect 16212 9454 16264 9460
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 15948 8430 15976 9318
rect 16040 9178 16068 9318
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15856 8214 15976 8242
rect 15948 8022 15976 8214
rect 15936 8016 15988 8022
rect 15936 7958 15988 7964
rect 15948 7721 15976 7958
rect 15934 7712 15990 7721
rect 15934 7647 15990 7656
rect 15948 7546 15976 7647
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15842 5672 15898 5681
rect 15842 5607 15898 5616
rect 15856 4758 15884 5607
rect 15948 5574 15976 6054
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 16040 5370 16068 5714
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 15844 4752 15896 4758
rect 15844 4694 15896 4700
rect 15856 4010 15884 4694
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 15934 4584 15990 4593
rect 15934 4519 15936 4528
rect 15988 4519 15990 4528
rect 15936 4490 15988 4496
rect 16040 4282 16068 4626
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 15844 4004 15896 4010
rect 15844 3946 15896 3952
rect 16132 3924 16160 9438
rect 16224 9178 16252 9454
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16316 7585 16344 10118
rect 16672 9920 16724 9926
rect 16486 9888 16542 9897
rect 16672 9862 16724 9868
rect 16486 9823 16542 9832
rect 16394 9752 16450 9761
rect 16394 9687 16450 9696
rect 16408 8090 16436 9687
rect 16500 8537 16528 9823
rect 16486 8528 16542 8537
rect 16684 8498 16712 9862
rect 16486 8463 16542 8472
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16684 8090 16712 8434
rect 17236 8129 17264 12378
rect 17316 12232 17368 12238
rect 17314 12200 17316 12209
rect 17368 12200 17370 12209
rect 17314 12135 17370 12144
rect 17328 11898 17356 12135
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17314 11656 17370 11665
rect 17314 11591 17370 11600
rect 17328 11257 17356 11591
rect 17420 11529 17448 12922
rect 17512 12442 17540 16186
rect 17696 16182 17724 18022
rect 17868 17604 17920 17610
rect 17868 17546 17920 17552
rect 17880 17270 17908 17546
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17972 17134 18000 19672
rect 18064 19174 18092 19858
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18064 18970 18092 19110
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17868 16788 17920 16794
rect 17920 16748 18000 16776
rect 17868 16730 17920 16736
rect 17776 16720 17828 16726
rect 17776 16662 17828 16668
rect 17788 16250 17816 16662
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17776 16244 17828 16250
rect 17776 16186 17828 16192
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17696 15609 17724 15642
rect 17880 15638 17908 16526
rect 17972 16046 18000 16748
rect 18064 16658 18092 17138
rect 18052 16652 18104 16658
rect 18052 16594 18104 16600
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 18050 16008 18106 16017
rect 18050 15943 18106 15952
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17868 15632 17920 15638
rect 17682 15600 17738 15609
rect 17868 15574 17920 15580
rect 17682 15535 17738 15544
rect 17972 15434 18000 15846
rect 18064 15586 18092 15943
rect 18156 15706 18184 18770
rect 18248 18698 18276 20454
rect 18328 20256 18380 20262
rect 18328 20198 18380 20204
rect 18340 19854 18368 20198
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18432 19242 18460 21286
rect 19076 21146 19104 21422
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18524 19310 18552 20742
rect 19076 20398 19104 20946
rect 19168 20942 19196 21490
rect 19260 21457 19288 21830
rect 19246 21448 19302 21457
rect 19246 21383 19302 21392
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 18696 20392 18748 20398
rect 18696 20334 18748 20340
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 18708 19718 18736 20334
rect 19168 20330 19196 20878
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 19168 19990 19196 20266
rect 19156 19984 19208 19990
rect 19156 19926 19208 19932
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18420 19236 18472 19242
rect 18420 19178 18472 19184
rect 18236 18692 18288 18698
rect 18236 18634 18288 18640
rect 18248 18290 18276 18634
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18248 17882 18276 18226
rect 18432 18154 18460 18566
rect 18420 18148 18472 18154
rect 18420 18090 18472 18096
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 18248 17678 18276 17818
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18248 16794 18276 17070
rect 18340 16794 18368 17682
rect 18602 17504 18658 17513
rect 18602 17439 18658 17448
rect 18616 17134 18644 17439
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18708 16998 18736 19654
rect 18970 19544 19026 19553
rect 18970 19479 19026 19488
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18800 18057 18828 18702
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 18892 18329 18920 18566
rect 18878 18320 18934 18329
rect 18878 18255 18934 18264
rect 18786 18048 18842 18057
rect 18786 17983 18842 17992
rect 18878 17232 18934 17241
rect 18878 17167 18880 17176
rect 18932 17167 18934 17176
rect 18880 17138 18932 17144
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 18524 16726 18552 16934
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18512 16720 18564 16726
rect 18512 16662 18564 16668
rect 18524 16114 18552 16662
rect 18616 16114 18644 16730
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18326 15872 18382 15881
rect 18326 15807 18382 15816
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18064 15558 18184 15586
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17972 15314 18000 15370
rect 17880 15286 18000 15314
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17512 11898 17540 12378
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17406 11520 17462 11529
rect 17406 11455 17462 11464
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17314 11248 17370 11257
rect 17314 11183 17370 11192
rect 17328 10130 17356 11183
rect 17406 10704 17462 10713
rect 17406 10639 17462 10648
rect 17420 10198 17448 10639
rect 17512 10266 17540 11290
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17604 10606 17632 11086
rect 17696 10690 17724 14350
rect 17788 13841 17816 14758
rect 17880 14618 17908 15286
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17774 13832 17830 13841
rect 17880 13818 17908 14418
rect 18064 14074 18092 14758
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17880 13790 18000 13818
rect 17774 13767 17830 13776
rect 17972 13462 18000 13790
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17788 10849 17816 12650
rect 17880 12442 17908 12718
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17880 11082 17908 12174
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17972 11286 18000 11630
rect 17960 11280 18012 11286
rect 17960 11222 18012 11228
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17774 10840 17830 10849
rect 17880 10810 17908 11018
rect 17774 10775 17830 10784
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17696 10662 17908 10690
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17408 10192 17460 10198
rect 17408 10134 17460 10140
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 9722 17356 10066
rect 17420 9722 17448 10134
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17788 9382 17816 9998
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17788 9110 17816 9318
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17604 8634 17632 8978
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17222 8120 17278 8129
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16672 8084 16724 8090
rect 17222 8055 17278 8064
rect 16672 8026 16724 8032
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16302 7576 16358 7585
rect 16302 7511 16358 7520
rect 16408 7342 16436 7822
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 7449 16528 7686
rect 16486 7440 16542 7449
rect 16486 7375 16488 7384
rect 16540 7375 16542 7384
rect 16488 7346 16540 7352
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 16224 7002 16252 7210
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16224 5681 16252 6938
rect 16408 6934 16436 7278
rect 16592 7206 16620 7822
rect 17236 7546 17264 7890
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16396 6928 16448 6934
rect 16592 6882 16620 7142
rect 16396 6870 16448 6876
rect 16500 6854 16620 6882
rect 16500 6662 16528 6854
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16304 6180 16356 6186
rect 16304 6122 16356 6128
rect 16210 5672 16266 5681
rect 16210 5607 16266 5616
rect 16316 4146 16344 6122
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16408 4826 16436 6054
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16408 4078 16436 4762
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 15934 3904 15990 3913
rect 16132 3896 16436 3924
rect 15934 3839 15990 3848
rect 15750 1048 15806 1057
rect 15750 983 15806 992
rect 15304 598 15516 626
rect 15304 480 15332 598
rect 15948 480 15976 3839
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 16132 2446 16160 3062
rect 16316 2854 16344 3130
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 16408 2514 16436 3896
rect 16578 3088 16634 3097
rect 16578 3023 16634 3032
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16408 2145 16436 2450
rect 16500 2310 16528 2926
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16394 2136 16450 2145
rect 16394 2071 16450 2080
rect 16592 480 16620 3023
rect 16684 2922 16712 7346
rect 17236 7313 17264 7482
rect 17880 7410 17908 10662
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17222 7304 17278 7313
rect 17222 7239 17278 7248
rect 17868 7268 17920 7274
rect 17868 7210 17920 7216
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16776 4554 16804 6190
rect 16868 6118 16896 6598
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16868 5914 16896 6054
rect 17144 5914 17172 6734
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17236 5846 17264 6734
rect 17788 6458 17816 6938
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17880 6322 17908 7210
rect 18156 6905 18184 15558
rect 18236 14544 18288 14550
rect 18236 14486 18288 14492
rect 18248 13870 18276 14486
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18248 13530 18276 13806
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18340 12850 18368 15807
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18418 14920 18474 14929
rect 18418 14855 18420 14864
rect 18472 14855 18474 14864
rect 18420 14826 18472 14832
rect 18512 14816 18564 14822
rect 18510 14784 18512 14793
rect 18564 14784 18566 14793
rect 18510 14719 18566 14728
rect 18616 14074 18644 14962
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18708 13977 18736 16934
rect 18880 16516 18932 16522
rect 18880 16458 18932 16464
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18694 13968 18750 13977
rect 18694 13903 18750 13912
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18800 12782 18828 16390
rect 18892 15706 18920 16458
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18892 14618 18920 15642
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18892 14074 18920 14554
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18248 12442 18276 12718
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18694 12336 18750 12345
rect 18694 12271 18750 12280
rect 18510 12200 18566 12209
rect 18510 12135 18566 12144
rect 18604 12164 18656 12170
rect 18326 10976 18382 10985
rect 18326 10911 18382 10920
rect 18340 10810 18368 10911
rect 18328 10804 18380 10810
rect 18380 10764 18460 10792
rect 18328 10746 18380 10752
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 18340 8090 18368 9318
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18142 6896 18198 6905
rect 18142 6831 18198 6840
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17500 6112 17552 6118
rect 17868 6112 17920 6118
rect 17500 6054 17552 6060
rect 17788 6060 17868 6066
rect 17788 6054 17920 6060
rect 17224 5840 17276 5846
rect 16854 5808 16910 5817
rect 17224 5782 17276 5788
rect 16854 5743 16910 5752
rect 16868 5370 16896 5743
rect 17236 5574 17264 5782
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16868 5166 16896 5306
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 17052 4729 17080 4966
rect 17038 4720 17094 4729
rect 17038 4655 17094 4664
rect 17236 4622 17264 5510
rect 17512 5137 17540 6054
rect 17788 6038 17908 6054
rect 17682 5264 17738 5273
rect 17682 5199 17738 5208
rect 17498 5128 17554 5137
rect 17498 5063 17554 5072
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 16764 4548 16816 4554
rect 16764 4490 16816 4496
rect 17236 3738 17264 4558
rect 17696 4146 17724 5199
rect 17788 4826 17816 6038
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17880 5352 17908 5850
rect 18248 5778 18276 7278
rect 18432 7002 18460 10764
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18524 6254 18552 12135
rect 18604 12106 18656 12112
rect 18616 11762 18644 12106
rect 18708 12102 18736 12271
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18708 11626 18736 12038
rect 18800 11898 18828 12038
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18800 11218 18828 11834
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18880 11212 18932 11218
rect 18880 11154 18932 11160
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18616 10266 18644 10542
rect 18708 10470 18736 11086
rect 18892 10985 18920 11154
rect 18878 10976 18934 10985
rect 18878 10911 18934 10920
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18708 6866 18736 10406
rect 18880 8560 18932 8566
rect 18880 8502 18932 8508
rect 18892 8401 18920 8502
rect 18878 8392 18934 8401
rect 18878 8327 18934 8336
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18708 6322 18736 6598
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18524 5574 18552 6190
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 17960 5364 18012 5370
rect 17880 5324 17960 5352
rect 17960 5306 18012 5312
rect 18418 5264 18474 5273
rect 18708 5234 18736 6258
rect 18418 5199 18474 5208
rect 18696 5228 18748 5234
rect 18432 5166 18460 5199
rect 18696 5170 18748 5176
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18064 4865 18092 4966
rect 18050 4856 18106 4865
rect 17776 4820 17828 4826
rect 18050 4791 18052 4800
rect 17776 4762 17828 4768
rect 18104 4791 18106 4800
rect 18052 4762 18104 4768
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17314 4040 17370 4049
rect 17314 3975 17370 3984
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 16764 3460 16816 3466
rect 16764 3402 16816 3408
rect 16776 3058 16804 3402
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 17222 2000 17278 2009
rect 17222 1935 17278 1944
rect 17236 1737 17264 1935
rect 17222 1728 17278 1737
rect 17222 1663 17278 1672
rect 17328 480 17356 3975
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 17958 3632 18014 3641
rect 17500 3596 17552 3602
rect 17958 3567 18014 3576
rect 17500 3538 17552 3544
rect 17512 3466 17540 3538
rect 17776 3528 17828 3534
rect 17774 3496 17776 3505
rect 17828 3496 17830 3505
rect 17500 3460 17552 3466
rect 17774 3431 17830 3440
rect 17500 3402 17552 3408
rect 17512 3194 17540 3402
rect 17500 3188 17552 3194
rect 17500 3130 17552 3136
rect 17774 2544 17830 2553
rect 17774 2479 17776 2488
rect 17828 2479 17830 2488
rect 17776 2450 17828 2456
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17604 1601 17632 2246
rect 17590 1592 17646 1601
rect 17590 1527 17646 1536
rect 17972 480 18000 3567
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 2650 18092 3334
rect 18248 3058 18276 3878
rect 18418 3496 18474 3505
rect 18418 3431 18474 3440
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 18432 2514 18460 3431
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 18616 2417 18644 4558
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18708 3641 18736 3878
rect 18694 3632 18750 3641
rect 18694 3567 18750 3576
rect 18800 3398 18828 4082
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18984 3194 19012 19479
rect 19352 18970 19380 19858
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 19260 18465 19288 18770
rect 19246 18456 19302 18465
rect 19246 18391 19302 18400
rect 19248 18080 19300 18086
rect 19300 18040 19380 18068
rect 19248 18022 19300 18028
rect 19352 17882 19380 18040
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19156 17060 19208 17066
rect 19156 17002 19208 17008
rect 19168 16697 19196 17002
rect 19260 16998 19288 17029
rect 19248 16992 19300 16998
rect 19246 16960 19248 16969
rect 19300 16960 19302 16969
rect 19246 16895 19302 16904
rect 19260 16794 19288 16895
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19154 16688 19210 16697
rect 19154 16623 19156 16632
rect 19208 16623 19210 16632
rect 19156 16594 19208 16600
rect 19352 16046 19380 17070
rect 19340 16040 19392 16046
rect 19076 15988 19340 15994
rect 19076 15982 19392 15988
rect 19076 15966 19380 15982
rect 19076 13802 19104 15966
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 19076 13530 19104 13738
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 19444 13462 19472 24670
rect 19536 23866 19564 25214
rect 20088 24682 20116 27520
rect 20168 25356 20220 25362
rect 20168 25298 20220 25304
rect 20076 24676 20128 24682
rect 20076 24618 20128 24624
rect 20180 24614 20208 25298
rect 20260 24744 20312 24750
rect 20258 24712 20260 24721
rect 20312 24712 20314 24721
rect 20258 24647 20314 24656
rect 20168 24608 20220 24614
rect 20074 24576 20130 24585
rect 19622 24508 19918 24528
rect 20168 24550 20220 24556
rect 20628 24608 20680 24614
rect 20732 24596 20760 27520
rect 20680 24568 20760 24596
rect 20628 24550 20680 24556
rect 20074 24511 20130 24520
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20088 24342 20116 24511
rect 20076 24336 20128 24342
rect 20076 24278 20128 24284
rect 19982 24168 20038 24177
rect 19982 24103 20038 24112
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19800 23112 19852 23118
rect 19800 23054 19852 23060
rect 19890 23080 19946 23089
rect 19812 22681 19840 23054
rect 19890 23015 19946 23024
rect 19798 22672 19854 22681
rect 19798 22607 19854 22616
rect 19904 22574 19932 23015
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19524 22228 19576 22234
rect 19524 22170 19576 22176
rect 19536 21146 19564 22170
rect 19708 22092 19760 22098
rect 19708 22034 19760 22040
rect 19720 21690 19748 22034
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19708 21684 19760 21690
rect 19708 21626 19760 21632
rect 19904 21554 19932 21966
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19524 21140 19576 21146
rect 19524 21082 19576 21088
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19798 19952 19854 19961
rect 19798 19887 19854 19896
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19628 19417 19656 19790
rect 19614 19408 19670 19417
rect 19614 19343 19670 19352
rect 19812 19310 19840 19887
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19536 18426 19564 18702
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19996 17377 20024 24103
rect 20076 23656 20128 23662
rect 20076 23598 20128 23604
rect 20088 22030 20116 23598
rect 20180 22817 20208 24550
rect 21376 24410 21404 27520
rect 22112 24834 22140 27520
rect 22756 25498 22784 27520
rect 22744 25492 22796 25498
rect 22744 25434 22796 25440
rect 22376 25356 22428 25362
rect 22376 25298 22428 25304
rect 22560 25356 22612 25362
rect 22560 25298 22612 25304
rect 22020 24806 22140 24834
rect 21916 24744 21968 24750
rect 21916 24686 21968 24692
rect 21928 24614 21956 24686
rect 22020 24682 22048 24806
rect 22008 24676 22060 24682
rect 22008 24618 22060 24624
rect 22388 24614 22416 25298
rect 22572 24886 22600 25298
rect 22560 24880 22612 24886
rect 22560 24822 22612 24828
rect 22468 24744 22520 24750
rect 22468 24686 22520 24692
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 22376 24608 22428 24614
rect 22480 24585 22508 24686
rect 22376 24550 22428 24556
rect 22466 24576 22522 24585
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 21732 24268 21784 24274
rect 21732 24210 21784 24216
rect 21744 23526 21772 24210
rect 21928 23746 21956 24550
rect 21928 23718 22048 23746
rect 21732 23520 21784 23526
rect 21638 23488 21694 23497
rect 21732 23462 21784 23468
rect 21638 23423 21694 23432
rect 20260 23180 20312 23186
rect 20260 23122 20312 23128
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20166 22808 20222 22817
rect 20166 22743 20222 22752
rect 20168 22568 20220 22574
rect 20168 22510 20220 22516
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 20088 21690 20116 21830
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 20088 17542 20116 18566
rect 20180 17660 20208 22510
rect 20272 22166 20300 23122
rect 20824 22545 20852 23122
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 20810 22536 20866 22545
rect 20810 22471 20812 22480
rect 20864 22471 20866 22480
rect 20812 22442 20864 22448
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20260 22160 20312 22166
rect 20260 22102 20312 22108
rect 20442 22128 20498 22137
rect 20732 22098 20760 22374
rect 20916 22234 20944 22918
rect 21008 22817 21036 23054
rect 20994 22808 21050 22817
rect 20994 22743 20996 22752
rect 21048 22743 21050 22752
rect 20996 22714 21048 22720
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 20904 22228 20956 22234
rect 20904 22170 20956 22176
rect 20442 22063 20498 22072
rect 20720 22092 20772 22098
rect 20180 17632 20300 17660
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 19982 17368 20038 17377
rect 19982 17303 20038 17312
rect 20088 17134 20116 17478
rect 20166 17368 20222 17377
rect 20166 17303 20222 17312
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20074 16416 20130 16425
rect 20074 16351 20130 16360
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19996 15502 20024 16186
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19996 15094 20024 15438
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19996 14618 20024 15030
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19260 12442 19288 13330
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 19168 11694 19196 12242
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19168 11286 19196 11630
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19260 11506 19288 11562
rect 19352 11506 19380 12786
rect 19522 12744 19578 12753
rect 19522 12679 19578 12688
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19444 12306 19472 12582
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19536 12238 19564 12679
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19260 11478 19380 11506
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19062 10568 19118 10577
rect 19062 10503 19064 10512
rect 19116 10503 19118 10512
rect 19064 10474 19116 10480
rect 19076 10266 19104 10474
rect 19352 10470 19380 11478
rect 19536 11354 19564 12174
rect 19904 11626 19932 12174
rect 19892 11620 19944 11626
rect 19892 11562 19944 11568
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19996 11354 20024 12242
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 19352 10033 19380 10202
rect 19338 10024 19394 10033
rect 19338 9959 19394 9968
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9178 19288 9862
rect 19352 9586 19380 9959
rect 19444 9586 19472 10542
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19156 8832 19208 8838
rect 19156 8774 19208 8780
rect 19168 7698 19196 8774
rect 19260 8430 19288 9114
rect 19340 8968 19392 8974
rect 19340 8910 19392 8916
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19248 8288 19300 8294
rect 19248 8230 19300 8236
rect 19260 8090 19288 8230
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19352 7857 19380 8910
rect 19432 7880 19484 7886
rect 19338 7848 19394 7857
rect 19432 7822 19484 7828
rect 19338 7783 19340 7792
rect 19392 7783 19394 7792
rect 19340 7754 19392 7760
rect 19168 7670 19380 7698
rect 19352 7546 19380 7670
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 19168 6390 19196 6802
rect 19156 6384 19208 6390
rect 19154 6352 19156 6361
rect 19208 6352 19210 6361
rect 19154 6287 19210 6296
rect 19260 5914 19288 7210
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19352 6186 19380 7142
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 19076 5370 19104 5782
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 19246 5128 19302 5137
rect 19246 5063 19302 5072
rect 19260 4826 19288 5063
rect 19338 4992 19394 5001
rect 19338 4927 19394 4936
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19154 3768 19210 3777
rect 19352 3738 19380 4927
rect 19154 3703 19210 3712
rect 19340 3732 19392 3738
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 18970 2680 19026 2689
rect 18970 2615 19026 2624
rect 18602 2408 18658 2417
rect 18602 2343 18658 2352
rect 18984 2145 19012 2615
rect 19168 2394 19196 3703
rect 19340 3674 19392 3680
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19260 2582 19288 2926
rect 19444 2922 19472 7822
rect 19536 6882 19564 11154
rect 19982 10704 20038 10713
rect 19982 10639 20038 10648
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19996 10266 20024 10639
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19628 9722 19656 10066
rect 19984 10056 20036 10062
rect 19706 10024 19762 10033
rect 19984 9998 20036 10004
rect 19706 9959 19762 9968
rect 19720 9761 19748 9959
rect 19706 9752 19762 9761
rect 19616 9716 19668 9722
rect 19706 9687 19762 9696
rect 19616 9658 19668 9664
rect 19996 9382 20024 9998
rect 20088 9602 20116 16351
rect 20180 12782 20208 17303
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 20180 9722 20208 12718
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20272 9625 20300 17632
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20364 16794 20392 17002
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20364 16250 20392 16730
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20350 15600 20406 15609
rect 20350 15535 20406 15544
rect 20364 15026 20392 15535
rect 20456 15042 20484 22063
rect 20720 22034 20772 22040
rect 20732 21894 20760 22034
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20916 21690 20944 21966
rect 20904 21684 20956 21690
rect 20904 21626 20956 21632
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20548 21146 20576 21422
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20732 20058 20760 20538
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20548 18630 20576 19858
rect 20824 19514 20852 20810
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20916 20505 20944 20742
rect 21008 20534 21036 20810
rect 20996 20528 21048 20534
rect 20902 20496 20958 20505
rect 20996 20470 21048 20476
rect 20902 20431 20958 20440
rect 20902 20360 20958 20369
rect 20902 20295 20904 20304
rect 20956 20295 20958 20304
rect 20904 20266 20956 20272
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 20916 19922 20944 19994
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 21100 19292 21128 22510
rect 21468 22098 21496 23054
rect 21548 22432 21600 22438
rect 21548 22374 21600 22380
rect 21560 22166 21588 22374
rect 21548 22160 21600 22166
rect 21548 22102 21600 22108
rect 21456 22092 21508 22098
rect 21456 22034 21508 22040
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21178 20360 21234 20369
rect 21178 20295 21234 20304
rect 21192 19825 21220 20295
rect 21284 20058 21312 21626
rect 21454 21584 21510 21593
rect 21454 21519 21510 21528
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 21376 20602 21404 20878
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21178 19816 21234 19825
rect 21178 19751 21234 19760
rect 21100 19264 21220 19292
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20536 18624 20588 18630
rect 20536 18566 20588 18572
rect 20718 18456 20774 18465
rect 20718 18391 20720 18400
rect 20772 18391 20774 18400
rect 20720 18362 20772 18368
rect 20536 16448 20588 16454
rect 20536 16390 20588 16396
rect 20548 15162 20576 16390
rect 20720 15632 20772 15638
rect 20718 15600 20720 15609
rect 20772 15600 20774 15609
rect 20718 15535 20774 15544
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20628 15496 20680 15502
rect 20680 15456 20760 15484
rect 20628 15438 20680 15444
rect 20536 15156 20588 15162
rect 20536 15098 20588 15104
rect 20352 15020 20404 15026
rect 20456 15014 20576 15042
rect 20352 14962 20404 14968
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 20352 11212 20404 11218
rect 20352 11154 20404 11160
rect 20364 10606 20392 11154
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 20364 10266 20392 10542
rect 20456 10538 20484 13942
rect 20548 12481 20576 15014
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20640 14414 20668 14758
rect 20732 14618 20760 15456
rect 20824 15094 20852 15506
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20824 14550 20852 15030
rect 20812 14544 20864 14550
rect 20812 14486 20864 14492
rect 20628 14408 20680 14414
rect 20812 14408 20864 14414
rect 20680 14368 20760 14396
rect 20628 14350 20680 14356
rect 20732 12850 20760 14368
rect 20812 14350 20864 14356
rect 20824 13870 20852 14350
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20534 12472 20590 12481
rect 20534 12407 20590 12416
rect 20732 11354 20760 12650
rect 20824 12374 20852 13806
rect 20916 13530 20944 19110
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 20996 18148 21048 18154
rect 20996 18090 21048 18096
rect 21008 14890 21036 18090
rect 21100 18086 21128 18770
rect 21192 18766 21220 19264
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 21192 18086 21220 18702
rect 21364 18352 21416 18358
rect 21362 18320 21364 18329
rect 21416 18320 21418 18329
rect 21362 18255 21418 18264
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21100 16153 21128 18022
rect 21180 17740 21232 17746
rect 21180 17682 21232 17688
rect 21192 17338 21220 17682
rect 21468 17490 21496 21519
rect 21548 20460 21600 20466
rect 21548 20402 21600 20408
rect 21560 19990 21588 20402
rect 21548 19984 21600 19990
rect 21548 19926 21600 19932
rect 21560 19514 21588 19926
rect 21548 19508 21600 19514
rect 21548 19450 21600 19456
rect 21560 18902 21588 19450
rect 21652 18970 21680 23423
rect 21744 21865 21772 23462
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21928 22574 21956 22918
rect 21916 22568 21968 22574
rect 21822 22536 21878 22545
rect 21916 22510 21968 22516
rect 21822 22471 21878 22480
rect 21730 21856 21786 21865
rect 21730 21791 21786 21800
rect 21836 19553 21864 22471
rect 21916 21344 21968 21350
rect 21916 21286 21968 21292
rect 21928 20602 21956 21286
rect 22020 21026 22048 23718
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 22112 22642 22140 23054
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22296 21486 22324 21830
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 22020 20998 22232 21026
rect 22008 20936 22060 20942
rect 22060 20884 22140 20890
rect 22008 20878 22140 20884
rect 22020 20862 22140 20878
rect 21916 20596 21968 20602
rect 21916 20538 21968 20544
rect 22112 20058 22140 20862
rect 22204 20369 22232 20998
rect 22190 20360 22246 20369
rect 22190 20295 22246 20304
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 21822 19544 21878 19553
rect 21822 19479 21878 19488
rect 22020 19446 22048 19994
rect 22008 19440 22060 19446
rect 22008 19382 22060 19388
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 21836 19258 21864 19314
rect 21836 19230 21956 19258
rect 21824 19168 21876 19174
rect 21824 19110 21876 19116
rect 21640 18964 21692 18970
rect 21640 18906 21692 18912
rect 21548 18896 21600 18902
rect 21548 18838 21600 18844
rect 21468 17462 21680 17490
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21468 16590 21496 17274
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21456 16584 21508 16590
rect 21508 16532 21588 16538
rect 21456 16526 21588 16532
rect 21086 16144 21142 16153
rect 21086 16079 21142 16088
rect 21376 15706 21404 16526
rect 21468 16510 21588 16526
rect 21560 16250 21588 16510
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 20996 14884 21048 14890
rect 20996 14826 21048 14832
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 20902 13288 20958 13297
rect 20902 13223 20958 13232
rect 20916 12782 20944 13223
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20812 12368 20864 12374
rect 20812 12310 20864 12316
rect 20916 12306 20944 12582
rect 20996 12368 21048 12374
rect 20996 12310 21048 12316
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20810 12200 20866 12209
rect 20810 12135 20866 12144
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20444 10532 20496 10538
rect 20444 10474 20496 10480
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20352 9716 20404 9722
rect 20352 9658 20404 9664
rect 20258 9616 20314 9625
rect 20088 9574 20208 9602
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19996 9110 20024 9318
rect 19984 9104 20036 9110
rect 19984 9046 20036 9052
rect 20088 8974 20116 9386
rect 20180 9042 20208 9574
rect 20258 9551 20314 9560
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 20088 8362 20116 8910
rect 20180 8430 20208 8978
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20088 7970 20116 8298
rect 20180 8265 20208 8366
rect 20166 8256 20222 8265
rect 20166 8191 20222 8200
rect 20364 7993 20392 9658
rect 20824 9466 20852 12135
rect 20916 11762 20944 12242
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20916 11218 20944 11698
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20824 9438 20944 9466
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20548 8430 20576 8774
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20824 8362 20852 9318
rect 20812 8356 20864 8362
rect 20812 8298 20864 8304
rect 19996 7942 20116 7970
rect 20350 7984 20406 7993
rect 19996 7478 20024 7942
rect 20350 7919 20406 7928
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 20088 7546 20116 7822
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 19984 7472 20036 7478
rect 19984 7414 20036 7420
rect 20916 7410 20944 9438
rect 21008 8922 21036 12310
rect 21086 10160 21142 10169
rect 21086 10095 21088 10104
rect 21140 10095 21142 10104
rect 21088 10066 21140 10072
rect 21100 9761 21128 10066
rect 21086 9752 21142 9761
rect 21086 9687 21142 9696
rect 21100 9110 21128 9687
rect 21088 9104 21140 9110
rect 21088 9046 21140 9052
rect 21008 8894 21128 8922
rect 20994 8392 21050 8401
rect 20994 8327 21050 8336
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19536 6854 19656 6882
rect 19628 6662 19656 6854
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19616 6656 19668 6662
rect 19616 6598 19668 6604
rect 19536 6118 19564 6598
rect 19628 6254 19656 6598
rect 19616 6248 19668 6254
rect 19614 6216 19616 6225
rect 19668 6216 19670 6225
rect 19614 6151 19670 6160
rect 19628 6125 19656 6151
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19536 5846 19564 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5840 19576 5846
rect 19524 5782 19576 5788
rect 19536 5166 19564 5782
rect 19982 5672 20038 5681
rect 19982 5607 20038 5616
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19536 4486 19564 5102
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4690 20024 5607
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19536 3505 19564 4422
rect 19996 4282 20024 4626
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19996 3738 20024 3878
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19522 3496 19578 3505
rect 19522 3431 19578 3440
rect 19890 3496 19946 3505
rect 19890 3431 19892 3440
rect 19944 3431 19946 3440
rect 19892 3402 19944 3408
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19430 2816 19486 2825
rect 19430 2751 19486 2760
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 19168 2366 19380 2394
rect 18970 2136 19026 2145
rect 18970 2071 19026 2080
rect 18694 1456 18750 1465
rect 18694 1391 18750 1400
rect 18708 480 18736 1391
rect 19352 480 19380 2366
rect 19444 1442 19472 2751
rect 19536 2650 19564 2994
rect 19904 2990 19932 3402
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 20088 2825 20116 4422
rect 20074 2816 20130 2825
rect 19622 2748 19918 2768
rect 20074 2751 20130 2760
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 20180 2514 20208 6734
rect 20456 5914 20484 6734
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20548 5846 20576 6190
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 20536 5636 20588 5642
rect 20536 5578 20588 5584
rect 20548 5166 20576 5578
rect 20536 5160 20588 5166
rect 20456 5108 20536 5114
rect 20456 5102 20588 5108
rect 20456 5086 20576 5102
rect 20456 4146 20484 5086
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20272 3738 20300 4014
rect 20548 4010 20576 4762
rect 20640 4078 20668 7142
rect 20916 7002 20944 7346
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20916 5914 20944 6598
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20732 4826 20760 5714
rect 20824 4826 20852 5850
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20916 5137 20944 5510
rect 20902 5128 20958 5137
rect 20902 5063 20958 5072
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20812 4820 20864 4826
rect 20812 4762 20864 4768
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20824 4457 20852 4626
rect 21008 4457 21036 8327
rect 21100 6497 21128 8894
rect 21086 6488 21142 6497
rect 21086 6423 21142 6432
rect 21100 4826 21128 6423
rect 21088 4820 21140 4826
rect 21088 4762 21140 4768
rect 20810 4448 20866 4457
rect 20810 4383 20866 4392
rect 20994 4448 21050 4457
rect 20994 4383 21050 4392
rect 20824 4282 20852 4383
rect 21100 4282 21128 4762
rect 20812 4276 20864 4282
rect 20812 4218 20864 4224
rect 21088 4276 21140 4282
rect 21088 4218 21140 4224
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20536 4004 20588 4010
rect 20536 3946 20588 3952
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 21192 3641 21220 14826
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21284 14385 21312 14758
rect 21364 14544 21416 14550
rect 21362 14512 21364 14521
rect 21416 14512 21418 14521
rect 21652 14498 21680 17462
rect 21732 16720 21784 16726
rect 21732 16662 21784 16668
rect 21744 15706 21772 16662
rect 21732 15700 21784 15706
rect 21732 15642 21784 15648
rect 21732 15564 21784 15570
rect 21732 15506 21784 15512
rect 21744 15337 21772 15506
rect 21730 15328 21786 15337
rect 21730 15263 21786 15272
rect 21744 14618 21772 15263
rect 21836 15065 21864 19110
rect 21928 18170 21956 19230
rect 22020 19174 22048 19382
rect 22192 19304 22244 19310
rect 22192 19246 22244 19252
rect 22008 19168 22060 19174
rect 22008 19110 22060 19116
rect 22098 18728 22154 18737
rect 22098 18663 22154 18672
rect 22112 18426 22140 18663
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 22112 18222 22140 18362
rect 22100 18216 22152 18222
rect 21928 18142 22048 18170
rect 22100 18158 22152 18164
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21928 16114 21956 18022
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 22020 15416 22048 18142
rect 21928 15388 22048 15416
rect 21822 15056 21878 15065
rect 21822 14991 21878 15000
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21652 14470 21772 14498
rect 21362 14447 21418 14456
rect 21270 14376 21326 14385
rect 21270 14311 21326 14320
rect 21376 13870 21404 14447
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21652 14074 21680 14350
rect 21640 14068 21692 14074
rect 21640 14010 21692 14016
rect 21364 13864 21416 13870
rect 21362 13832 21364 13841
rect 21416 13832 21418 13841
rect 21362 13767 21418 13776
rect 21744 11286 21772 14470
rect 21824 14476 21876 14482
rect 21824 14418 21876 14424
rect 21836 14074 21864 14418
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21928 13954 21956 15388
rect 22204 15314 22232 19246
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22296 17241 22324 17478
rect 22282 17232 22338 17241
rect 22282 17167 22338 17176
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22296 16046 22324 16730
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22284 15904 22336 15910
rect 22284 15846 22336 15852
rect 22296 15706 22324 15846
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22020 15286 22232 15314
rect 22020 14929 22048 15286
rect 22296 15026 22324 15642
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22006 14920 22062 14929
rect 22006 14855 22062 14864
rect 22296 14414 22324 14962
rect 22388 14550 22416 24550
rect 22466 24511 22522 24520
rect 22468 21004 22520 21010
rect 22468 20946 22520 20952
rect 22480 20534 22508 20946
rect 22468 20528 22520 20534
rect 22468 20470 22520 20476
rect 22572 19242 22600 24822
rect 23124 24410 23152 27639
rect 23478 27520 23534 28000
rect 24122 27520 24178 28000
rect 24766 27520 24822 28000
rect 25502 27520 25558 28000
rect 26146 27520 26202 28000
rect 26882 27520 26938 28000
rect 27526 27520 27582 28000
rect 23202 27160 23258 27169
rect 23202 27095 23258 27104
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 23020 24268 23072 24274
rect 23020 24210 23072 24216
rect 23032 23526 23060 24210
rect 23216 23866 23244 27095
rect 23296 24608 23348 24614
rect 23492 24596 23520 27520
rect 23662 26616 23718 26625
rect 23662 26551 23718 26560
rect 23348 24568 23520 24596
rect 23296 24550 23348 24556
rect 23676 24410 23704 26551
rect 24136 25430 24164 27520
rect 24780 26058 24808 27520
rect 24596 26030 24808 26058
rect 24596 25498 24624 26030
rect 24766 25936 24822 25945
rect 24766 25871 24822 25880
rect 24780 25498 24808 25871
rect 24584 25492 24636 25498
rect 24584 25434 24636 25440
rect 24768 25492 24820 25498
rect 24768 25434 24820 25440
rect 24124 25424 24176 25430
rect 24124 25366 24176 25372
rect 24766 25392 24822 25401
rect 23940 25356 23992 25362
rect 24766 25327 24822 25336
rect 23940 25298 23992 25304
rect 23848 24744 23900 24750
rect 23848 24686 23900 24692
rect 23664 24404 23716 24410
rect 23664 24346 23716 24352
rect 23386 24304 23442 24313
rect 23386 24239 23442 24248
rect 23480 24268 23532 24274
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 23020 23520 23072 23526
rect 23020 23462 23072 23468
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 22940 22438 22968 23122
rect 22928 22432 22980 22438
rect 22928 22374 22980 22380
rect 22650 21584 22706 21593
rect 22650 21519 22706 21528
rect 22664 21146 22692 21519
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22650 21040 22706 21049
rect 22650 20975 22706 20984
rect 22664 20602 22692 20975
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 22836 20392 22888 20398
rect 22836 20334 22888 20340
rect 22650 19816 22706 19825
rect 22650 19751 22706 19760
rect 22560 19236 22612 19242
rect 22560 19178 22612 19184
rect 22664 19174 22692 19751
rect 22652 19168 22704 19174
rect 22652 19110 22704 19116
rect 22742 19000 22798 19009
rect 22742 18935 22744 18944
rect 22796 18935 22798 18944
rect 22744 18906 22796 18912
rect 22560 18828 22612 18834
rect 22560 18770 22612 18776
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22480 14958 22508 18226
rect 22572 18193 22600 18770
rect 22558 18184 22614 18193
rect 22558 18119 22614 18128
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22664 17338 22692 17682
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22756 16794 22784 16934
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22376 14544 22428 14550
rect 22376 14486 22428 14492
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 21836 13926 21956 13954
rect 22100 13932 22152 13938
rect 21732 11280 21784 11286
rect 21652 11240 21732 11268
rect 21454 10976 21510 10985
rect 21454 10911 21510 10920
rect 21362 10840 21418 10849
rect 21362 10775 21364 10784
rect 21416 10775 21418 10784
rect 21364 10746 21416 10752
rect 21468 10305 21496 10911
rect 21454 10296 21510 10305
rect 21454 10231 21510 10240
rect 21364 10056 21416 10062
rect 21364 9998 21416 10004
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21284 8090 21312 9862
rect 21376 9489 21404 9998
rect 21362 9480 21418 9489
rect 21362 9415 21364 9424
rect 21416 9415 21418 9424
rect 21364 9386 21416 9392
rect 21376 8945 21404 9386
rect 21468 9178 21496 9998
rect 21652 9897 21680 11240
rect 21732 11222 21784 11228
rect 21730 10976 21786 10985
rect 21730 10911 21786 10920
rect 21744 10606 21772 10911
rect 21732 10600 21784 10606
rect 21732 10542 21784 10548
rect 21638 9888 21694 9897
rect 21638 9823 21694 9832
rect 21456 9172 21508 9178
rect 21456 9114 21508 9120
rect 21548 8968 21600 8974
rect 21362 8936 21418 8945
rect 21548 8910 21600 8916
rect 21362 8871 21418 8880
rect 21560 8430 21588 8910
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21284 7546 21312 8026
rect 21560 7750 21588 8366
rect 21640 8356 21692 8362
rect 21640 8298 21692 8304
rect 21652 7886 21680 8298
rect 21640 7880 21692 7886
rect 21640 7822 21692 7828
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21468 7410 21496 7686
rect 21652 7478 21680 7822
rect 21730 7712 21786 7721
rect 21730 7647 21786 7656
rect 21640 7472 21692 7478
rect 21744 7449 21772 7647
rect 21640 7414 21692 7420
rect 21730 7440 21786 7449
rect 21456 7404 21508 7410
rect 21730 7375 21786 7384
rect 21456 7346 21508 7352
rect 21362 7304 21418 7313
rect 21362 7239 21418 7248
rect 21272 6928 21324 6934
rect 21272 6870 21324 6876
rect 21284 6497 21312 6870
rect 21270 6488 21326 6497
rect 21270 6423 21326 6432
rect 21376 5710 21404 7239
rect 21468 6769 21496 7346
rect 21548 6792 21600 6798
rect 21454 6760 21510 6769
rect 21548 6734 21600 6740
rect 21454 6695 21510 6704
rect 21468 6186 21496 6695
rect 21560 6458 21588 6734
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 21456 6180 21508 6186
rect 21456 6122 21508 6128
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21376 5370 21404 5646
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21468 4622 21496 6122
rect 21560 5642 21588 6394
rect 21836 5658 21864 13926
rect 22100 13874 22152 13880
rect 22112 13462 22140 13874
rect 22296 13870 22324 14214
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22204 13530 22232 13670
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 22020 12306 22048 13262
rect 22204 12986 22232 13466
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 22112 12442 22140 12582
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22008 12300 22060 12306
rect 22008 12242 22060 12248
rect 22296 11354 22324 13806
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22388 12850 22416 13330
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 22664 12442 22692 12786
rect 22848 12782 22876 20334
rect 22940 19378 22968 22374
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 23032 17513 23060 23462
rect 23110 20360 23166 20369
rect 23110 20295 23166 20304
rect 23018 17504 23074 17513
rect 23018 17439 23074 17448
rect 23124 17218 23152 20295
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23216 19514 23244 19858
rect 23296 19780 23348 19786
rect 23296 19722 23348 19728
rect 23204 19508 23256 19514
rect 23204 19450 23256 19456
rect 23308 19446 23336 19722
rect 23296 19440 23348 19446
rect 23296 19382 23348 19388
rect 23308 19310 23336 19382
rect 23204 19304 23256 19310
rect 23202 19272 23204 19281
rect 23296 19304 23348 19310
rect 23256 19272 23258 19281
rect 23296 19246 23348 19252
rect 23202 19207 23258 19216
rect 23400 18850 23428 24239
rect 23480 24210 23532 24216
rect 23492 23526 23520 24210
rect 23572 23588 23624 23594
rect 23572 23530 23624 23536
rect 23480 23520 23532 23526
rect 23480 23462 23532 23468
rect 23492 23254 23520 23462
rect 23584 23254 23612 23530
rect 23480 23248 23532 23254
rect 23480 23190 23532 23196
rect 23572 23248 23624 23254
rect 23572 23190 23624 23196
rect 23756 23180 23808 23186
rect 23756 23122 23808 23128
rect 23768 22778 23796 23122
rect 23860 22953 23888 24686
rect 23952 24614 23980 25298
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24780 24954 24808 25327
rect 24768 24948 24820 24954
rect 24768 24890 24820 24896
rect 24122 24848 24178 24857
rect 24122 24783 24178 24792
rect 23940 24608 23992 24614
rect 23940 24550 23992 24556
rect 23846 22944 23902 22953
rect 23846 22879 23902 22888
rect 23572 22772 23624 22778
rect 23572 22714 23624 22720
rect 23756 22772 23808 22778
rect 23756 22714 23808 22720
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23492 20466 23520 20742
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23492 19990 23520 20402
rect 23480 19984 23532 19990
rect 23480 19926 23532 19932
rect 23492 19242 23520 19926
rect 23480 19236 23532 19242
rect 23480 19178 23532 19184
rect 23492 18970 23520 19178
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23296 18828 23348 18834
rect 23400 18822 23520 18850
rect 23296 18770 23348 18776
rect 23308 18290 23336 18770
rect 23492 18766 23520 18822
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23296 18284 23348 18290
rect 23296 18226 23348 18232
rect 23296 18148 23348 18154
rect 23296 18090 23348 18096
rect 23308 18057 23336 18090
rect 23492 18086 23520 18702
rect 23480 18080 23532 18086
rect 23294 18048 23350 18057
rect 23294 17983 23350 17992
rect 23400 18040 23480 18068
rect 23400 17898 23428 18040
rect 23480 18022 23532 18028
rect 23308 17870 23428 17898
rect 23124 17190 23244 17218
rect 23020 16652 23072 16658
rect 23020 16594 23072 16600
rect 23032 16046 23060 16594
rect 23020 16040 23072 16046
rect 23020 15982 23072 15988
rect 23020 14952 23072 14958
rect 23020 14894 23072 14900
rect 22926 13832 22982 13841
rect 22926 13767 22982 13776
rect 22836 12776 22888 12782
rect 22836 12718 22888 12724
rect 22652 12436 22704 12442
rect 22652 12378 22704 12384
rect 22468 12300 22520 12306
rect 22468 12242 22520 12248
rect 22480 11898 22508 12242
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 21916 11008 21968 11014
rect 21916 10950 21968 10956
rect 21928 10470 21956 10950
rect 22204 10810 22232 11222
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22006 10704 22062 10713
rect 22006 10639 22062 10648
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 21928 7857 21956 10406
rect 22020 10033 22048 10639
rect 22480 10266 22508 11834
rect 22664 11150 22692 12378
rect 22940 12306 22968 13767
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22006 10024 22062 10033
rect 22006 9959 22062 9968
rect 22192 9920 22244 9926
rect 22020 9868 22192 9874
rect 22020 9862 22244 9868
rect 22020 9846 22232 9862
rect 22020 9654 22048 9846
rect 22008 9648 22060 9654
rect 22008 9590 22060 9596
rect 22190 9616 22246 9625
rect 22480 9586 22508 10202
rect 22572 9926 22600 11086
rect 22560 9920 22612 9926
rect 22560 9862 22612 9868
rect 22190 9551 22246 9560
rect 22468 9580 22520 9586
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 22112 8634 22140 8978
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 21914 7848 21970 7857
rect 21914 7783 21970 7792
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21928 5846 21956 7686
rect 22204 7342 22232 9551
rect 22468 9522 22520 9528
rect 23032 9466 23060 14894
rect 23112 14884 23164 14890
rect 23112 14826 23164 14832
rect 23124 14074 23152 14826
rect 23216 14346 23244 17190
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23202 13696 23258 13705
rect 23202 13631 23258 13640
rect 23112 11620 23164 11626
rect 23112 11562 23164 11568
rect 23124 9654 23152 11562
rect 23216 10849 23244 13631
rect 23202 10840 23258 10849
rect 23202 10775 23258 10784
rect 23112 9648 23164 9654
rect 23112 9590 23164 9596
rect 22572 9438 23060 9466
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 22006 6896 22062 6905
rect 22006 6831 22062 6840
rect 22020 6730 22048 6831
rect 22008 6724 22060 6730
rect 22008 6666 22060 6672
rect 22008 5908 22060 5914
rect 22008 5850 22060 5856
rect 21916 5840 21968 5846
rect 21916 5782 21968 5788
rect 22020 5658 22048 5850
rect 21548 5636 21600 5642
rect 21836 5630 21956 5658
rect 22020 5630 22140 5658
rect 21548 5578 21600 5584
rect 21928 4808 21956 5630
rect 22112 5370 22140 5630
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 21928 4780 22048 4808
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 21270 4312 21326 4321
rect 21270 4247 21326 4256
rect 21178 3632 21234 3641
rect 21178 3567 21234 3576
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 20732 2990 20760 3402
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20732 2650 20760 2926
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 20718 1864 20774 1873
rect 20718 1799 20774 1808
rect 19444 1414 20116 1442
rect 20088 480 20116 1414
rect 20732 480 20760 1799
rect 21284 610 21312 4247
rect 21468 3738 21496 4558
rect 21640 4208 21692 4214
rect 21638 4176 21640 4185
rect 21692 4176 21694 4185
rect 21638 4111 21694 4120
rect 21456 3732 21508 3738
rect 21456 3674 21508 3680
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 21272 604 21324 610
rect 21272 546 21324 552
rect 21376 480 21404 3062
rect 21928 2854 21956 3538
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 21928 2689 21956 2790
rect 21914 2680 21970 2689
rect 22020 2650 22048 4780
rect 22098 4584 22154 4593
rect 22098 4519 22154 4528
rect 21914 2615 21970 2624
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 22112 480 22140 4519
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 22296 3942 22324 4150
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 22388 3097 22416 7142
rect 22572 4826 22600 9438
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 23032 9081 23060 9318
rect 23018 9072 23074 9081
rect 23018 9007 23074 9016
rect 23308 8514 23336 17870
rect 23480 17604 23532 17610
rect 23480 17546 23532 17552
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 23400 17202 23428 17478
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 23492 17134 23520 17546
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23478 16416 23534 16425
rect 23478 16351 23534 16360
rect 23492 16250 23520 16351
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23492 15178 23520 15438
rect 23400 15162 23520 15178
rect 23388 15156 23520 15162
rect 23440 15150 23520 15156
rect 23388 15098 23440 15104
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23400 13546 23428 13874
rect 23400 13530 23520 13546
rect 23400 13524 23532 13530
rect 23400 13518 23480 13524
rect 23480 13466 23532 13472
rect 23492 12986 23520 13466
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23584 12866 23612 22714
rect 23952 22642 23980 24550
rect 24032 24268 24084 24274
rect 24032 24210 24084 24216
rect 24044 23526 24072 24210
rect 24032 23520 24084 23526
rect 24032 23462 24084 23468
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 23664 22568 23716 22574
rect 23662 22536 23664 22545
rect 23716 22536 23718 22545
rect 23662 22471 23718 22480
rect 24044 22098 24072 23462
rect 23756 22092 23808 22098
rect 23756 22034 23808 22040
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 23768 21350 23796 22034
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23676 18970 23704 20878
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23676 17377 23704 17614
rect 23662 17368 23718 17377
rect 23662 17303 23664 17312
rect 23716 17303 23718 17312
rect 23664 17274 23716 17280
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 23676 16250 23704 17138
rect 23768 16998 23796 21286
rect 23952 21146 23980 21422
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 23940 21004 23992 21010
rect 23940 20946 23992 20952
rect 23952 20602 23980 20946
rect 23940 20596 23992 20602
rect 23940 20538 23992 20544
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23860 19281 23888 20198
rect 23952 20058 23980 20538
rect 24032 20256 24084 20262
rect 24032 20198 24084 20204
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 24044 19961 24072 20198
rect 24030 19952 24086 19961
rect 24030 19887 24086 19896
rect 23846 19272 23902 19281
rect 23846 19207 23902 19216
rect 23846 17504 23902 17513
rect 23846 17439 23902 17448
rect 23756 16992 23808 16998
rect 23756 16934 23808 16940
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 23860 15978 23888 17439
rect 23848 15972 23900 15978
rect 23848 15914 23900 15920
rect 23860 15722 23888 15914
rect 23860 15706 23980 15722
rect 23848 15700 23980 15706
rect 23900 15694 23980 15700
rect 23848 15642 23900 15648
rect 23848 15564 23900 15570
rect 23848 15506 23900 15512
rect 23756 15428 23808 15434
rect 23756 15370 23808 15376
rect 23768 15337 23796 15370
rect 23754 15328 23810 15337
rect 23754 15263 23810 15272
rect 23768 15162 23796 15263
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23664 14952 23716 14958
rect 23664 14894 23716 14900
rect 23676 13938 23704 14894
rect 23860 14618 23888 15506
rect 23952 15026 23980 15694
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23938 14920 23994 14929
rect 23938 14855 23994 14864
rect 23848 14612 23900 14618
rect 23848 14554 23900 14560
rect 23848 14408 23900 14414
rect 23848 14350 23900 14356
rect 23860 14074 23888 14350
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23664 13932 23716 13938
rect 23664 13874 23716 13880
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23400 12838 23612 12866
rect 23400 12288 23428 12838
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23676 12374 23704 12718
rect 23754 12472 23810 12481
rect 23860 12442 23888 13874
rect 23754 12407 23810 12416
rect 23848 12436 23900 12442
rect 23664 12368 23716 12374
rect 23664 12310 23716 12316
rect 23400 12260 23520 12288
rect 23388 10056 23440 10062
rect 23386 10024 23388 10033
rect 23440 10024 23442 10033
rect 23386 9959 23442 9968
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 22756 8486 23336 8514
rect 22650 7576 22706 7585
rect 22650 7511 22706 7520
rect 22664 6866 22692 7511
rect 22652 6860 22704 6866
rect 22652 6802 22704 6808
rect 22664 6458 22692 6802
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 22756 5370 22784 8486
rect 23296 8424 23348 8430
rect 23296 8366 23348 8372
rect 23202 8256 23258 8265
rect 23202 8191 23258 8200
rect 23110 7848 23166 7857
rect 23110 7783 23166 7792
rect 23020 7200 23072 7206
rect 23020 7142 23072 7148
rect 23032 6798 23060 7142
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 22928 6656 22980 6662
rect 22928 6598 22980 6604
rect 22836 5840 22888 5846
rect 22836 5782 22888 5788
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22756 5273 22784 5306
rect 22742 5264 22798 5273
rect 22742 5199 22798 5208
rect 22756 5166 22784 5199
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22480 4214 22508 4422
rect 22468 4208 22520 4214
rect 22468 4150 22520 4156
rect 22572 4078 22600 4762
rect 22664 4185 22692 4966
rect 22848 4826 22876 5782
rect 22836 4820 22888 4826
rect 22836 4762 22888 4768
rect 22834 4720 22890 4729
rect 22834 4655 22890 4664
rect 22650 4176 22706 4185
rect 22650 4111 22706 4120
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22756 3398 22784 3538
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 22374 3088 22430 3097
rect 22374 3023 22430 3032
rect 22756 2446 22784 3334
rect 22744 2440 22796 2446
rect 22744 2382 22796 2388
rect 22848 1034 22876 4655
rect 22940 2990 22968 6598
rect 23032 5914 23060 6734
rect 23124 6458 23152 7783
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23124 6254 23152 6394
rect 23112 6248 23164 6254
rect 23112 6190 23164 6196
rect 23020 5908 23072 5914
rect 23020 5850 23072 5856
rect 23216 5273 23244 8191
rect 23308 7954 23336 8366
rect 23400 7954 23428 8774
rect 23296 7948 23348 7954
rect 23296 7890 23348 7896
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 23388 7268 23440 7274
rect 23388 7210 23440 7216
rect 23296 6996 23348 7002
rect 23296 6938 23348 6944
rect 23308 6662 23336 6938
rect 23400 6730 23428 7210
rect 23388 6724 23440 6730
rect 23388 6666 23440 6672
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 23202 5264 23258 5273
rect 23202 5199 23258 5208
rect 23296 4684 23348 4690
rect 23296 4626 23348 4632
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 23308 4146 23336 4626
rect 23400 4214 23428 4626
rect 23492 4282 23520 12260
rect 23676 11914 23704 12310
rect 23584 11886 23704 11914
rect 23584 11354 23612 11886
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23676 11558 23704 11698
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23572 11348 23624 11354
rect 23572 11290 23624 11296
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23584 10266 23612 11086
rect 23676 10810 23704 11494
rect 23768 11082 23796 12407
rect 23848 12378 23900 12384
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23860 11506 23888 12242
rect 23952 11665 23980 14855
rect 24032 14476 24084 14482
rect 24032 14418 24084 14424
rect 24044 13870 24072 14418
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 24044 11801 24072 13806
rect 24136 12714 24164 24783
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24676 24064 24728 24070
rect 24676 24006 24728 24012
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24216 23656 24268 23662
rect 24216 23598 24268 23604
rect 24228 21554 24256 23598
rect 24688 23089 24716 24006
rect 24780 23633 24808 24550
rect 24766 23624 24822 23633
rect 24766 23559 24822 23568
rect 24768 23520 24820 23526
rect 25516 23497 25544 27520
rect 25778 24168 25834 24177
rect 25778 24103 25834 24112
rect 24768 23462 24820 23468
rect 25502 23488 25558 23497
rect 24674 23080 24730 23089
rect 24674 23015 24730 23024
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24780 22545 24808 23462
rect 25502 23423 25558 23432
rect 25044 23180 25096 23186
rect 25044 23122 25096 23128
rect 25056 22778 25084 23122
rect 25320 22976 25372 22982
rect 25320 22918 25372 22924
rect 25044 22772 25096 22778
rect 25044 22714 25096 22720
rect 24950 22672 25006 22681
rect 24950 22607 25006 22616
rect 24964 22574 24992 22607
rect 24952 22568 25004 22574
rect 24766 22536 24822 22545
rect 24952 22510 25004 22516
rect 24766 22471 24822 22480
rect 24676 22432 24728 22438
rect 24676 22374 24728 22380
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24216 21548 24268 21554
rect 24216 21490 24268 21496
rect 24688 20777 24716 22374
rect 25044 22092 25096 22098
rect 25044 22034 25096 22040
rect 25056 22001 25084 22034
rect 25042 21992 25098 22001
rect 25042 21927 25098 21936
rect 24860 21888 24912 21894
rect 24780 21836 24860 21842
rect 24780 21830 24912 21836
rect 24780 21814 24900 21830
rect 24674 20768 24730 20777
rect 24289 20700 24585 20720
rect 24674 20703 24730 20712
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24780 20097 24808 21814
rect 25056 21690 25084 21927
rect 25044 21684 25096 21690
rect 25044 21626 25096 21632
rect 25228 21480 25280 21486
rect 25226 21448 25228 21457
rect 25280 21448 25282 21457
rect 25226 21383 25282 21392
rect 25332 21321 25360 22918
rect 25504 22772 25556 22778
rect 25504 22714 25556 22720
rect 25516 21554 25544 22714
rect 25504 21548 25556 21554
rect 25504 21490 25556 21496
rect 25318 21312 25374 21321
rect 25318 21247 25374 21256
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 24860 20936 24912 20942
rect 25148 20913 25176 20946
rect 24860 20878 24912 20884
rect 25134 20904 25190 20913
rect 24872 20602 24900 20878
rect 25134 20839 25190 20848
rect 25148 20602 25176 20839
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 24860 20596 24912 20602
rect 24860 20538 24912 20544
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 24766 20088 24822 20097
rect 24766 20023 24822 20032
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24872 19514 24900 20538
rect 25226 20496 25282 20505
rect 25226 20431 25282 20440
rect 25240 20398 25268 20431
rect 25228 20392 25280 20398
rect 25228 20334 25280 20340
rect 25240 20058 25268 20334
rect 25228 20052 25280 20058
rect 25228 19994 25280 20000
rect 25332 19553 25360 20742
rect 25318 19544 25374 19553
rect 24860 19508 24912 19514
rect 25318 19479 25374 19488
rect 24860 19450 24912 19456
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24766 18320 24822 18329
rect 24766 18255 24822 18264
rect 24492 18216 24544 18222
rect 24492 18158 24544 18164
rect 24504 17882 24532 18158
rect 24492 17876 24544 17882
rect 24492 17818 24544 17824
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24228 17105 24256 17138
rect 24214 17096 24270 17105
rect 24214 17031 24270 17040
rect 24228 16794 24256 17031
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16114 24716 17614
rect 24780 16697 24808 18255
rect 24872 18222 24900 19450
rect 25226 19408 25282 19417
rect 25226 19343 25282 19352
rect 24952 19304 25004 19310
rect 24952 19246 25004 19252
rect 24964 18630 24992 19246
rect 25240 18834 25268 19343
rect 25228 18828 25280 18834
rect 25228 18770 25280 18776
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 24964 18154 24992 18566
rect 25240 18426 25268 18770
rect 25412 18624 25464 18630
rect 25412 18566 25464 18572
rect 25424 18465 25452 18566
rect 25410 18456 25466 18465
rect 25228 18420 25280 18426
rect 25410 18391 25466 18400
rect 25228 18362 25280 18368
rect 24952 18148 25004 18154
rect 24952 18090 25004 18096
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24766 16688 24822 16697
rect 24766 16623 24822 16632
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24766 16008 24822 16017
rect 24766 15943 24822 15952
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24492 14884 24544 14890
rect 24492 14826 24544 14832
rect 24504 14414 24532 14826
rect 24492 14408 24544 14414
rect 24214 14376 24270 14385
rect 24492 14350 24544 14356
rect 24214 14311 24270 14320
rect 24124 12708 24176 12714
rect 24124 12650 24176 12656
rect 24122 12608 24178 12617
rect 24122 12543 24178 12552
rect 24030 11792 24086 11801
rect 24030 11727 24086 11736
rect 24136 11694 24164 12543
rect 24228 12345 24256 14311
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24400 13796 24452 13802
rect 24400 13738 24452 13744
rect 24412 13258 24440 13738
rect 24688 13530 24716 15506
rect 24676 13524 24728 13530
rect 24676 13466 24728 13472
rect 24400 13252 24452 13258
rect 24400 13194 24452 13200
rect 24780 13138 24808 15943
rect 24872 14618 24900 17682
rect 24964 17542 24992 18090
rect 25136 18080 25188 18086
rect 25042 18048 25098 18057
rect 25136 18022 25188 18028
rect 25042 17983 25098 17992
rect 25056 17746 25084 17983
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24964 16726 24992 17478
rect 25056 16794 25084 17682
rect 25148 17678 25176 18022
rect 25228 17876 25280 17882
rect 25228 17818 25280 17824
rect 25240 17785 25268 17818
rect 25226 17776 25282 17785
rect 25226 17711 25282 17720
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25226 17640 25282 17649
rect 25148 17338 25176 17614
rect 25226 17575 25282 17584
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25240 17134 25268 17575
rect 25410 17232 25466 17241
rect 25410 17167 25466 17176
rect 25228 17128 25280 17134
rect 25228 17070 25280 17076
rect 25424 16794 25452 17167
rect 25504 17060 25556 17066
rect 25504 17002 25556 17008
rect 25044 16788 25096 16794
rect 25044 16730 25096 16736
rect 25412 16788 25464 16794
rect 25412 16730 25464 16736
rect 24952 16720 25004 16726
rect 24952 16662 25004 16668
rect 24964 15978 24992 16662
rect 25516 16658 25544 17002
rect 25504 16652 25556 16658
rect 25504 16594 25556 16600
rect 25410 16144 25466 16153
rect 25410 16079 25412 16088
rect 25464 16079 25466 16088
rect 25412 16050 25464 16056
rect 24952 15972 25004 15978
rect 24952 15914 25004 15920
rect 24964 15366 24992 15914
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 25056 15706 25084 15846
rect 25044 15700 25096 15706
rect 25044 15642 25096 15648
rect 24952 15360 25004 15366
rect 24952 15302 25004 15308
rect 24964 14890 24992 15302
rect 24952 14884 25004 14890
rect 24952 14826 25004 14832
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24964 14550 24992 14826
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 24964 13870 24992 14486
rect 25504 14340 25556 14346
rect 25504 14282 25556 14288
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 25516 13734 25544 14282
rect 25504 13728 25556 13734
rect 25504 13670 25556 13676
rect 25134 13424 25190 13433
rect 24952 13388 25004 13394
rect 25134 13359 25190 13368
rect 24952 13330 25004 13336
rect 24688 13110 24808 13138
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12866 24716 13110
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24596 12838 24716 12866
rect 24214 12336 24270 12345
rect 24214 12271 24270 12280
rect 24596 12209 24624 12838
rect 24676 12708 24728 12714
rect 24676 12650 24728 12656
rect 24582 12200 24638 12209
rect 24582 12135 24638 12144
rect 24216 12096 24268 12102
rect 24216 12038 24268 12044
rect 24124 11688 24176 11694
rect 23938 11656 23994 11665
rect 24124 11630 24176 11636
rect 24228 11626 24256 12038
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24306 11656 24362 11665
rect 23938 11591 23994 11600
rect 24216 11620 24268 11626
rect 24306 11591 24362 11600
rect 24216 11562 24268 11568
rect 24032 11552 24084 11558
rect 23860 11478 23980 11506
rect 24032 11494 24084 11500
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23756 11076 23808 11082
rect 23756 11018 23808 11024
rect 23664 10804 23716 10810
rect 23664 10746 23716 10752
rect 23768 10538 23796 11018
rect 23860 10742 23888 11290
rect 23848 10736 23900 10742
rect 23848 10678 23900 10684
rect 23756 10532 23808 10538
rect 23756 10474 23808 10480
rect 23572 10260 23624 10266
rect 23572 10202 23624 10208
rect 23664 10124 23716 10130
rect 23664 10066 23716 10072
rect 23572 10056 23624 10062
rect 23572 9998 23624 10004
rect 23584 9450 23612 9998
rect 23676 9518 23704 10066
rect 23952 10010 23980 11478
rect 24044 11218 24072 11494
rect 24032 11212 24084 11218
rect 24032 11154 24084 11160
rect 24044 10198 24072 11154
rect 24320 11121 24348 11591
rect 24306 11112 24362 11121
rect 24306 11047 24362 11056
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24124 10804 24176 10810
rect 24124 10746 24176 10752
rect 24136 10606 24164 10746
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24032 10192 24084 10198
rect 24032 10134 24084 10140
rect 24136 10062 24164 10542
rect 24124 10056 24176 10062
rect 23952 9982 24072 10010
rect 24124 9998 24176 10004
rect 23756 9920 23808 9926
rect 23756 9862 23808 9868
rect 23846 9888 23902 9897
rect 23768 9586 23796 9862
rect 23846 9823 23902 9832
rect 23756 9580 23808 9586
rect 23756 9522 23808 9528
rect 23664 9512 23716 9518
rect 23664 9454 23716 9460
rect 23572 9444 23624 9450
rect 23572 9386 23624 9392
rect 23676 9382 23704 9454
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 23570 8936 23626 8945
rect 23570 8871 23626 8880
rect 23584 8242 23612 8871
rect 23676 8537 23704 9318
rect 23662 8528 23718 8537
rect 23662 8463 23718 8472
rect 23768 8430 23796 9522
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 23584 8214 23796 8242
rect 23662 8120 23718 8129
rect 23662 8055 23718 8064
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 23584 7206 23612 7890
rect 23572 7200 23624 7206
rect 23572 7142 23624 7148
rect 23676 6610 23704 8055
rect 23584 6582 23704 6610
rect 23584 6390 23612 6582
rect 23662 6488 23718 6497
rect 23662 6423 23664 6432
rect 23716 6423 23718 6432
rect 23664 6394 23716 6400
rect 23572 6384 23624 6390
rect 23572 6326 23624 6332
rect 23584 6186 23612 6326
rect 23572 6180 23624 6186
rect 23572 6122 23624 6128
rect 23572 5840 23624 5846
rect 23572 5782 23624 5788
rect 23584 5370 23612 5782
rect 23768 5681 23796 8214
rect 23860 7177 23888 9823
rect 23940 9444 23992 9450
rect 23940 9386 23992 9392
rect 23952 8974 23980 9386
rect 23940 8968 23992 8974
rect 23940 8910 23992 8916
rect 24044 8786 24072 9982
rect 24136 9382 24164 9998
rect 24124 9376 24176 9382
rect 24124 9318 24176 9324
rect 24136 9178 24164 9318
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 23952 8758 24072 8786
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 23846 7168 23902 7177
rect 23846 7103 23902 7112
rect 23754 5672 23810 5681
rect 23754 5607 23810 5616
rect 23572 5364 23624 5370
rect 23572 5306 23624 5312
rect 23584 4826 23612 5306
rect 23572 4820 23624 4826
rect 23572 4762 23624 4768
rect 23570 4448 23626 4457
rect 23570 4383 23626 4392
rect 23480 4276 23532 4282
rect 23480 4218 23532 4224
rect 23388 4208 23440 4214
rect 23388 4150 23440 4156
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23308 3738 23336 4082
rect 23388 4072 23440 4078
rect 23388 4014 23440 4020
rect 23400 3754 23428 4014
rect 23478 3768 23534 3777
rect 23296 3732 23348 3738
rect 23400 3726 23478 3754
rect 23478 3703 23534 3712
rect 23296 3674 23348 3680
rect 23308 3534 23336 3674
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23584 3194 23612 4383
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 23584 2990 23612 3130
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 22928 2984 22980 2990
rect 22928 2926 22980 2932
rect 23572 2984 23624 2990
rect 23860 2961 23888 2994
rect 23572 2926 23624 2932
rect 23846 2952 23902 2961
rect 23846 2887 23902 2896
rect 23756 2508 23808 2514
rect 23756 2450 23808 2456
rect 23768 2310 23796 2450
rect 23756 2304 23808 2310
rect 23756 2246 23808 2252
rect 23768 1737 23796 2246
rect 23754 1728 23810 1737
rect 23754 1663 23810 1672
rect 22756 1006 22876 1034
rect 22756 480 22784 1006
rect 23480 604 23532 610
rect 23480 546 23532 552
rect 23492 480 23520 546
rect 294 0 350 480
rect 938 0 994 480
rect 1582 0 1638 480
rect 2318 0 2374 480
rect 2962 0 3018 480
rect 3698 0 3754 480
rect 4342 0 4398 480
rect 4986 0 5042 480
rect 5722 0 5778 480
rect 6366 0 6422 480
rect 7102 0 7158 480
rect 7746 0 7802 480
rect 8390 0 8446 480
rect 9126 0 9182 480
rect 9770 0 9826 480
rect 10506 0 10562 480
rect 11150 0 11206 480
rect 11886 0 11942 480
rect 12530 0 12586 480
rect 13174 0 13230 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15290 0 15346 480
rect 15934 0 15990 480
rect 16578 0 16634 480
rect 17314 0 17370 480
rect 17958 0 18014 480
rect 18694 0 18750 480
rect 19338 0 19394 480
rect 20074 0 20130 480
rect 20718 0 20774 480
rect 21362 0 21418 480
rect 22098 0 22154 480
rect 22742 0 22798 480
rect 23478 0 23534 480
rect 23952 377 23980 8758
rect 24136 8616 24164 8774
rect 24044 8588 24164 8616
rect 24044 8022 24072 8588
rect 24228 8514 24256 10950
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24136 8486 24256 8514
rect 24032 8016 24084 8022
rect 24032 7958 24084 7964
rect 24044 7342 24072 7958
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 24032 7200 24084 7206
rect 24032 7142 24084 7148
rect 24044 5234 24072 7142
rect 24136 6905 24164 8486
rect 24216 8356 24268 8362
rect 24216 8298 24268 8304
rect 24228 7750 24256 8298
rect 24216 7744 24268 7750
rect 24688 7721 24716 12650
rect 24780 12442 24808 12922
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 24768 11620 24820 11626
rect 24768 11562 24820 11568
rect 24780 11506 24808 11562
rect 24780 11478 24900 11506
rect 24872 10266 24900 11478
rect 24860 10260 24912 10266
rect 24860 10202 24912 10208
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24780 8566 24808 8910
rect 24768 8560 24820 8566
rect 24768 8502 24820 8508
rect 24216 7686 24268 7692
rect 24674 7712 24730 7721
rect 24228 7410 24256 7686
rect 24289 7644 24585 7664
rect 24674 7647 24730 7656
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24780 7562 24808 8502
rect 24872 8430 24900 8978
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 24872 7954 24900 8366
rect 24860 7948 24912 7954
rect 24860 7890 24912 7896
rect 24688 7534 24808 7562
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24122 6896 24178 6905
rect 24122 6831 24178 6840
rect 24214 6760 24270 6769
rect 24214 6695 24216 6704
rect 24268 6695 24270 6704
rect 24216 6666 24268 6672
rect 24124 6656 24176 6662
rect 24124 6598 24176 6604
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 24136 5098 24164 6598
rect 24228 6322 24256 6666
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 24228 5914 24256 6258
rect 24216 5908 24268 5914
rect 24216 5850 24268 5856
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5234 24716 7534
rect 24766 7440 24822 7449
rect 24766 7375 24822 7384
rect 24780 6769 24808 7375
rect 24964 6798 24992 13330
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 25056 12986 25084 13262
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 25056 11694 25084 12242
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 25056 9110 25084 11630
rect 25148 11218 25176 13359
rect 25516 13326 25544 13670
rect 25688 13388 25740 13394
rect 25688 13330 25740 13336
rect 25504 13320 25556 13326
rect 25504 13262 25556 13268
rect 25228 13252 25280 13258
rect 25228 13194 25280 13200
rect 25240 12646 25268 13194
rect 25700 13161 25728 13330
rect 25686 13152 25742 13161
rect 25686 13087 25742 13096
rect 25700 12918 25728 13087
rect 25688 12912 25740 12918
rect 25688 12854 25740 12860
rect 25228 12640 25280 12646
rect 25228 12582 25280 12588
rect 25240 12238 25268 12582
rect 25504 12368 25556 12374
rect 25504 12310 25556 12316
rect 25320 12300 25372 12306
rect 25320 12242 25372 12248
rect 25228 12232 25280 12238
rect 25228 12174 25280 12180
rect 25240 11354 25268 12174
rect 25332 11558 25360 12242
rect 25320 11552 25372 11558
rect 25320 11494 25372 11500
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 25148 10810 25176 11154
rect 25136 10804 25188 10810
rect 25136 10746 25188 10752
rect 25134 10024 25190 10033
rect 25134 9959 25190 9968
rect 25044 9104 25096 9110
rect 25042 9072 25044 9081
rect 25096 9072 25098 9081
rect 25042 9007 25098 9016
rect 25056 8090 25084 9007
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 25148 7002 25176 9959
rect 25332 8906 25360 11494
rect 25516 11370 25544 12310
rect 25594 11792 25650 11801
rect 25594 11727 25596 11736
rect 25648 11727 25650 11736
rect 25596 11698 25648 11704
rect 25516 11342 25636 11370
rect 25792 11354 25820 24103
rect 26160 19825 26188 27520
rect 26896 25226 26924 27520
rect 26884 25220 26936 25226
rect 26884 25162 26936 25168
rect 27540 21049 27568 27520
rect 27526 21040 27582 21049
rect 27526 20975 27582 20984
rect 26146 19816 26202 19825
rect 26146 19751 26202 19760
rect 25964 16652 26016 16658
rect 25964 16594 26016 16600
rect 25976 16250 26004 16594
rect 25964 16244 26016 16250
rect 25964 16186 26016 16192
rect 25964 13320 26016 13326
rect 25964 13262 26016 13268
rect 25976 12918 26004 13262
rect 25964 12912 26016 12918
rect 25964 12854 26016 12860
rect 25320 8900 25372 8906
rect 25320 8842 25372 8848
rect 25410 7712 25466 7721
rect 25410 7647 25466 7656
rect 25424 7546 25452 7647
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25228 7336 25280 7342
rect 25226 7304 25228 7313
rect 25280 7304 25282 7313
rect 25226 7239 25282 7248
rect 25412 7200 25464 7206
rect 25412 7142 25464 7148
rect 25136 6996 25188 7002
rect 25136 6938 25188 6944
rect 25042 6896 25098 6905
rect 25042 6831 25098 6840
rect 24952 6792 25004 6798
rect 24766 6760 24822 6769
rect 24952 6734 25004 6740
rect 24766 6695 24822 6704
rect 24964 6458 24992 6734
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 24860 6248 24912 6254
rect 24780 6196 24860 6202
rect 24780 6190 24912 6196
rect 24780 6174 24900 6190
rect 24780 5370 24808 6174
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24124 5092 24176 5098
rect 24124 5034 24176 5040
rect 24136 4758 24164 5034
rect 24216 4820 24268 4826
rect 24216 4762 24268 4768
rect 24124 4752 24176 4758
rect 24124 4694 24176 4700
rect 24228 4128 24256 4762
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 25056 4162 25084 6831
rect 25148 5914 25176 6938
rect 25320 6860 25372 6866
rect 25320 6802 25372 6808
rect 25136 5908 25188 5914
rect 25136 5850 25188 5856
rect 25226 5264 25282 5273
rect 25226 5199 25282 5208
rect 25240 5166 25268 5199
rect 25228 5160 25280 5166
rect 25228 5102 25280 5108
rect 24308 4140 24360 4146
rect 24228 4100 24308 4128
rect 24032 4072 24084 4078
rect 24032 4014 24084 4020
rect 24044 3942 24072 4014
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 24228 3738 24256 4100
rect 24308 4082 24360 4088
rect 24952 4140 25004 4146
rect 25056 4134 25176 4162
rect 24952 4082 25004 4088
rect 24768 3936 24820 3942
rect 24820 3884 24900 3890
rect 24768 3878 24900 3884
rect 24780 3862 24900 3878
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 24674 3632 24730 3641
rect 24124 3596 24176 3602
rect 24674 3567 24730 3576
rect 24124 3538 24176 3544
rect 24136 3194 24164 3538
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 24122 3088 24178 3097
rect 24122 3023 24178 3032
rect 24136 480 24164 3023
rect 24582 2952 24638 2961
rect 24582 2887 24638 2896
rect 24490 2680 24546 2689
rect 24596 2650 24624 2887
rect 24688 2689 24716 3567
rect 24766 2816 24822 2825
rect 24766 2751 24822 2760
rect 24674 2680 24730 2689
rect 24490 2615 24546 2624
rect 24584 2644 24636 2650
rect 24504 2446 24532 2615
rect 24674 2615 24730 2624
rect 24584 2586 24636 2592
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24780 480 24808 2751
rect 24872 2650 24900 3862
rect 24964 3738 24992 4082
rect 25044 4072 25096 4078
rect 25044 4014 25096 4020
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 25056 3194 25084 4014
rect 25044 3188 25096 3194
rect 25044 3130 25096 3136
rect 25148 2990 25176 4134
rect 25332 4078 25360 6802
rect 25424 6798 25452 7142
rect 25412 6792 25464 6798
rect 25412 6734 25464 6740
rect 25424 5914 25452 6734
rect 25504 6180 25556 6186
rect 25504 6122 25556 6128
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 25516 5817 25544 6122
rect 25502 5808 25558 5817
rect 25502 5743 25558 5752
rect 25608 4457 25636 11342
rect 25780 11348 25832 11354
rect 25780 11290 25832 11296
rect 25688 8900 25740 8906
rect 25688 8842 25740 8848
rect 25700 8362 25728 8842
rect 25688 8356 25740 8362
rect 25688 8298 25740 8304
rect 25700 5001 25728 8298
rect 26884 5296 26936 5302
rect 26884 5238 26936 5244
rect 25686 4992 25742 5001
rect 25686 4927 25742 4936
rect 25594 4448 25650 4457
rect 25594 4383 25650 4392
rect 26146 4176 26202 4185
rect 26146 4111 26202 4120
rect 25320 4072 25372 4078
rect 25320 4014 25372 4020
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 25424 3505 25452 3878
rect 25410 3496 25466 3505
rect 25410 3431 25466 3440
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 25228 2916 25280 2922
rect 25228 2858 25280 2864
rect 24860 2644 24912 2650
rect 24860 2586 24912 2592
rect 25240 2553 25268 2858
rect 25226 2544 25282 2553
rect 25226 2479 25282 2488
rect 25502 1592 25558 1601
rect 25502 1527 25558 1536
rect 25516 480 25544 1527
rect 26160 480 26188 4111
rect 26896 480 26924 5238
rect 27526 3496 27582 3505
rect 27526 3431 27582 3440
rect 27540 480 27568 3431
rect 23938 368 23994 377
rect 23938 303 23994 312
rect 24122 0 24178 480
rect 24766 0 24822 480
rect 25502 0 25558 480
rect 26146 0 26202 480
rect 26882 0 26938 480
rect 27526 0 27582 480
<< via2 >>
rect 23110 27648 23166 27704
rect 938 24112 994 24168
rect 1582 22616 1638 22672
rect 1582 13912 1638 13968
rect 386 12824 442 12880
rect 1490 12416 1546 12472
rect 2962 21392 3018 21448
rect 4342 24248 4398 24304
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 4986 23296 5042 23352
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 3698 20440 3754 20496
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 6366 24656 6422 24712
rect 7746 22752 7802 22808
rect 9126 24792 9182 24848
rect 9678 24656 9734 24712
rect 9586 23296 9642 23352
rect 9586 21936 9642 21992
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 9770 23568 9826 23624
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10598 22772 10654 22808
rect 10598 22752 10600 22772
rect 10600 22752 10652 22772
rect 10652 22752 10654 22772
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10782 22888 10838 22944
rect 10874 22752 10930 22808
rect 10138 21664 10194 21720
rect 9678 20848 9734 20904
rect 5998 17856 6054 17912
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 9954 20712 10010 20768
rect 9586 19352 9642 19408
rect 9494 18828 9550 18864
rect 9494 18808 9496 18828
rect 9496 18808 9548 18828
rect 9548 18808 9550 18828
rect 9770 19216 9826 19272
rect 8298 15952 8354 16008
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 11334 24520 11390 24576
rect 11150 21548 11206 21584
rect 11150 21528 11152 21548
rect 11152 21528 11204 21548
rect 11204 21528 11206 21548
rect 10966 20576 11022 20632
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10874 20032 10930 20088
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 9954 13912 10010 13968
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 9126 12824 9182 12880
rect 2318 12416 2374 12472
rect 2042 11056 2098 11112
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 9494 12724 9496 12744
rect 9496 12724 9548 12744
rect 9548 12724 9550 12744
rect 9494 12688 9550 12724
rect 9586 11600 9642 11656
rect 9218 11192 9274 11248
rect 8942 11056 8998 11112
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 2778 10648 2834 10704
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10138 18264 10194 18320
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10138 17856 10194 17912
rect 11886 24384 11942 24440
rect 12162 24248 12218 24304
rect 11518 20884 11520 20904
rect 11520 20884 11572 20904
rect 11572 20884 11574 20904
rect 11518 20848 11574 20884
rect 10782 17212 10784 17232
rect 10784 17212 10836 17232
rect 10836 17212 10838 17232
rect 10782 17176 10838 17212
rect 11334 17584 11390 17640
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 12806 24656 12862 24712
rect 13726 24404 13782 24440
rect 13726 24384 13728 24404
rect 13728 24384 13780 24404
rect 13780 24384 13782 24404
rect 14186 24792 14242 24848
rect 14370 24792 14426 24848
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14554 24656 14610 24712
rect 12530 23296 12586 23352
rect 12254 22480 12310 22536
rect 12714 22924 12716 22944
rect 12716 22924 12768 22944
rect 12768 22924 12770 22944
rect 12714 22888 12770 22924
rect 12714 21684 12770 21720
rect 12714 21664 12716 21684
rect 12716 21664 12768 21684
rect 12768 21664 12770 21684
rect 12346 20304 12402 20360
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 9862 11056 9918 11112
rect 9310 10668 9366 10704
rect 9310 10648 9312 10668
rect 9312 10648 9364 10668
rect 9364 10648 9366 10668
rect 9586 10648 9642 10704
rect 4986 10104 5042 10160
rect 2318 8880 2374 8936
rect 294 4392 350 4448
rect 938 4120 994 4176
rect 1582 2488 1638 2544
rect 3790 7928 3846 7984
rect 3698 6840 3754 6896
rect 2962 5208 3018 5264
rect 3698 4664 3754 4720
rect 4342 7384 4398 7440
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 7102 8472 7158 8528
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 6366 6704 6422 6760
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5722 1808 5778 1864
rect 7746 7792 7802 7848
rect 9586 6296 9642 6352
rect 9770 9016 9826 9072
rect 8390 3304 8446 3360
rect 8758 1536 8814 1592
rect 9218 2372 9274 2408
rect 9218 2352 9220 2372
rect 9220 2352 9272 2372
rect 9272 2352 9274 2372
rect 9862 6296 9918 6352
rect 10046 3460 10102 3496
rect 10046 3440 10048 3460
rect 10048 3440 10100 3460
rect 10100 3440 10102 3460
rect 9954 2488 10010 2544
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 11058 13368 11114 13424
rect 10966 12008 11022 12064
rect 10782 8916 10784 8936
rect 10784 8916 10836 8936
rect 10836 8916 10838 8936
rect 10782 8880 10838 8916
rect 11794 17176 11850 17232
rect 11886 16244 11942 16280
rect 11886 16224 11888 16244
rect 11888 16224 11940 16244
rect 11940 16224 11942 16244
rect 11242 9560 11298 9616
rect 11150 7384 11206 7440
rect 11518 11872 11574 11928
rect 11702 10920 11758 10976
rect 11518 9016 11574 9072
rect 11242 6704 11298 6760
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 11334 5652 11336 5672
rect 11336 5652 11388 5672
rect 11388 5652 11390 5672
rect 11334 5616 11390 5652
rect 11334 4972 11336 4992
rect 11336 4972 11388 4992
rect 11388 4972 11390 4992
rect 11334 4936 11390 4972
rect 11150 3576 11206 3632
rect 11426 3884 11428 3904
rect 11428 3884 11480 3904
rect 11480 3884 11482 3904
rect 11426 3848 11482 3884
rect 11426 3712 11482 3768
rect 10322 3068 10324 3088
rect 10324 3068 10376 3088
rect 10376 3068 10378 3088
rect 10322 3032 10378 3068
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10966 1400 11022 1456
rect 12070 17876 12126 17912
rect 12070 17856 12072 17876
rect 12072 17856 12124 17876
rect 12124 17856 12126 17876
rect 12070 15680 12126 15736
rect 12530 20168 12586 20224
rect 13726 23568 13782 23624
rect 13358 22616 13414 22672
rect 12622 19896 12678 19952
rect 12438 18264 12494 18320
rect 12714 18148 12770 18184
rect 12714 18128 12716 18148
rect 12716 18128 12768 18148
rect 12768 18128 12770 18148
rect 11978 9288 12034 9344
rect 12714 12824 12770 12880
rect 12622 12008 12678 12064
rect 12346 11228 12348 11248
rect 12348 11228 12400 11248
rect 12400 11228 12402 11248
rect 12346 11192 12402 11228
rect 13174 17060 13230 17096
rect 13174 17040 13176 17060
rect 13176 17040 13228 17060
rect 13228 17040 13230 17060
rect 13726 23024 13782 23080
rect 14278 24112 14334 24168
rect 14094 22752 14150 22808
rect 14002 20440 14058 20496
rect 13358 19352 13414 19408
rect 13818 20032 13874 20088
rect 13818 17856 13874 17912
rect 13450 16904 13506 16960
rect 13266 14320 13322 14376
rect 13358 13948 13360 13968
rect 13360 13948 13412 13968
rect 13412 13948 13414 13968
rect 13358 13912 13414 13948
rect 13174 13232 13230 13288
rect 12898 12552 12954 12608
rect 11978 6840 12034 6896
rect 12070 6704 12126 6760
rect 11886 5344 11942 5400
rect 11794 3304 11850 3360
rect 13174 12552 13230 12608
rect 13174 12300 13230 12336
rect 13174 12280 13176 12300
rect 13176 12280 13228 12300
rect 13228 12280 13230 12300
rect 12806 7792 12862 7848
rect 11610 1808 11666 1864
rect 11978 2760 12034 2816
rect 12714 3712 12770 3768
rect 12714 2796 12716 2816
rect 12716 2796 12768 2816
rect 12768 2796 12770 2816
rect 12714 2760 12770 2796
rect 12898 3712 12954 3768
rect 13174 9444 13230 9480
rect 13174 9424 13176 9444
rect 13176 9424 13228 9444
rect 13228 9424 13230 9444
rect 13082 7656 13138 7712
rect 13358 12552 13414 12608
rect 14370 23296 14426 23352
rect 14278 19760 14334 19816
rect 13726 15544 13782 15600
rect 14462 18264 14518 18320
rect 14094 16496 14150 16552
rect 14186 16224 14242 16280
rect 13818 15000 13874 15056
rect 14002 14456 14058 14512
rect 13818 13912 13874 13968
rect 13542 12144 13598 12200
rect 13910 11872 13966 11928
rect 14002 11756 14058 11792
rect 14002 11736 14004 11756
rect 14004 11736 14056 11756
rect 14056 11736 14058 11756
rect 13358 10104 13414 10160
rect 13634 9968 13690 10024
rect 14002 10376 14058 10432
rect 14002 9968 14058 10024
rect 13910 9560 13966 9616
rect 13450 7928 13506 7984
rect 13634 7792 13690 7848
rect 13818 5072 13874 5128
rect 13634 4528 13690 4584
rect 13266 3712 13322 3768
rect 13542 3712 13598 3768
rect 15934 24792 15990 24848
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15290 23296 15346 23352
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14738 21936 14794 21992
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14646 21412 14702 21448
rect 14646 21392 14648 21412
rect 14648 21392 14700 21412
rect 14700 21392 14702 21412
rect 14554 16632 14610 16688
rect 14186 11328 14242 11384
rect 14370 11328 14426 11384
rect 14370 9052 14372 9072
rect 14372 9052 14424 9072
rect 14424 9052 14426 9072
rect 14370 9016 14426 9052
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14738 19352 14794 19408
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14830 19216 14886 19272
rect 15566 21972 15568 21992
rect 15568 21972 15620 21992
rect 15620 21972 15622 21992
rect 15566 21936 15622 21972
rect 15658 20440 15714 20496
rect 15474 19760 15530 19816
rect 14830 18808 14886 18864
rect 15290 18692 15346 18728
rect 15290 18672 15292 18692
rect 15292 18672 15344 18692
rect 15344 18672 15346 18692
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14830 17992 14886 18048
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15934 22752 15990 22808
rect 15750 19352 15806 19408
rect 15474 15680 15530 15736
rect 15474 15544 15530 15600
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15290 12688 15346 12744
rect 15382 12416 15438 12472
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14738 11056 14794 11112
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14830 10512 14886 10568
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14738 9560 14794 9616
rect 14278 6704 14334 6760
rect 14462 6840 14518 6896
rect 14554 5344 14610 5400
rect 14554 4800 14610 4856
rect 13174 2916 13230 2952
rect 13174 2896 13176 2916
rect 13176 2896 13228 2916
rect 13228 2896 13230 2916
rect 12898 2624 12954 2680
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14922 6704 14978 6760
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14830 6160 14886 6216
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15382 10376 15438 10432
rect 15382 9696 15438 9752
rect 15382 9288 15438 9344
rect 15474 9152 15530 9208
rect 16118 22888 16174 22944
rect 16026 17584 16082 17640
rect 16026 12824 16082 12880
rect 16762 19216 16818 19272
rect 17130 20304 17186 20360
rect 16394 16632 16450 16688
rect 16302 15816 16358 15872
rect 15934 12552 15990 12608
rect 15934 12416 15990 12472
rect 15750 12280 15806 12336
rect 15658 9832 15714 9888
rect 15290 4528 15346 4584
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15566 4256 15622 4312
rect 15474 3984 15530 4040
rect 15474 3440 15530 3496
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14278 2488 14334 2544
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15382 1672 15438 1728
rect 14554 1536 14610 1592
rect 15842 9832 15898 9888
rect 16210 12280 16266 12336
rect 16854 16496 16910 16552
rect 16670 15680 16726 15736
rect 16486 15408 16542 15464
rect 16486 14728 16542 14784
rect 16394 12824 16450 12880
rect 16394 12724 16396 12744
rect 16396 12724 16448 12744
rect 16448 12724 16450 12744
rect 16394 12688 16450 12724
rect 16302 11600 16358 11656
rect 16578 12280 16634 12336
rect 16302 10240 16358 10296
rect 17682 20168 17738 20224
rect 17222 17584 17278 17640
rect 17038 14728 17094 14784
rect 17958 24404 18014 24440
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 17958 24384 17960 24404
rect 17960 24384 18012 24404
rect 18012 24384 18014 24404
rect 18970 24112 19026 24168
rect 19154 23296 19210 23352
rect 17406 13912 17462 13968
rect 16762 12144 16818 12200
rect 16946 11056 17002 11112
rect 15934 7656 15990 7712
rect 15842 5616 15898 5672
rect 15934 4548 15990 4584
rect 15934 4528 15936 4548
rect 15936 4528 15988 4548
rect 15988 4528 15990 4548
rect 16486 9832 16542 9888
rect 16394 9696 16450 9752
rect 16486 8472 16542 8528
rect 17314 12180 17316 12200
rect 17316 12180 17368 12200
rect 17368 12180 17370 12200
rect 17314 12144 17370 12180
rect 17314 11600 17370 11656
rect 18050 15952 18106 16008
rect 17682 15544 17738 15600
rect 19246 21392 19302 21448
rect 18602 17448 18658 17504
rect 18970 19488 19026 19544
rect 18878 18264 18934 18320
rect 18786 17992 18842 18048
rect 18878 17196 18934 17232
rect 18878 17176 18880 17196
rect 18880 17176 18932 17196
rect 18932 17176 18934 17196
rect 18326 15816 18382 15872
rect 17406 11464 17462 11520
rect 17314 11192 17370 11248
rect 17406 10648 17462 10704
rect 17774 13776 17830 13832
rect 17774 10784 17830 10840
rect 17222 8064 17278 8120
rect 16302 7520 16358 7576
rect 16486 7404 16542 7440
rect 16486 7384 16488 7404
rect 16488 7384 16540 7404
rect 16540 7384 16542 7404
rect 16210 5616 16266 5672
rect 15934 3848 15990 3904
rect 15750 992 15806 1048
rect 16578 3032 16634 3088
rect 16394 2080 16450 2136
rect 17222 7248 17278 7304
rect 18418 14884 18474 14920
rect 18418 14864 18420 14884
rect 18420 14864 18472 14884
rect 18472 14864 18474 14884
rect 18510 14764 18512 14784
rect 18512 14764 18564 14784
rect 18564 14764 18566 14784
rect 18510 14728 18566 14764
rect 18694 13912 18750 13968
rect 18694 12280 18750 12336
rect 18510 12144 18566 12200
rect 18326 10920 18382 10976
rect 18142 6840 18198 6896
rect 16854 5752 16910 5808
rect 17038 4664 17094 4720
rect 17682 5208 17738 5264
rect 17498 5072 17554 5128
rect 18878 10920 18934 10976
rect 18878 8336 18934 8392
rect 18418 5208 18474 5264
rect 18050 4820 18106 4856
rect 18050 4800 18052 4820
rect 18052 4800 18104 4820
rect 18104 4800 18106 4820
rect 17314 3984 17370 4040
rect 17222 1944 17278 2000
rect 17222 1672 17278 1728
rect 17958 3576 18014 3632
rect 17774 3476 17776 3496
rect 17776 3476 17828 3496
rect 17828 3476 17830 3496
rect 17774 3440 17830 3476
rect 17774 2508 17830 2544
rect 17774 2488 17776 2508
rect 17776 2488 17828 2508
rect 17828 2488 17830 2508
rect 17590 1536 17646 1592
rect 18418 3440 18474 3496
rect 18694 3576 18750 3632
rect 19246 18400 19302 18456
rect 19246 16940 19248 16960
rect 19248 16940 19300 16960
rect 19300 16940 19302 16960
rect 19246 16904 19302 16940
rect 19154 16652 19210 16688
rect 19154 16632 19156 16652
rect 19156 16632 19208 16652
rect 19208 16632 19210 16652
rect 20258 24692 20260 24712
rect 20260 24692 20312 24712
rect 20312 24692 20314 24712
rect 20258 24656 20314 24692
rect 20074 24520 20130 24576
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19982 24112 20038 24168
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19890 23024 19946 23080
rect 19798 22616 19854 22672
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19798 19896 19854 19952
rect 19614 19352 19670 19408
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 21638 23432 21694 23488
rect 20166 22752 20222 22808
rect 20810 22500 20866 22536
rect 20810 22480 20812 22500
rect 20812 22480 20864 22500
rect 20864 22480 20866 22500
rect 20442 22072 20498 22128
rect 20994 22772 21050 22808
rect 20994 22752 20996 22772
rect 20996 22752 21048 22772
rect 21048 22752 21050 22772
rect 19982 17312 20038 17368
rect 20166 17312 20222 17368
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 20074 16360 20130 16416
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19522 12688 19578 12744
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19062 10532 19118 10568
rect 19062 10512 19064 10532
rect 19064 10512 19116 10532
rect 19116 10512 19118 10532
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19338 9968 19394 10024
rect 19338 7812 19394 7848
rect 19338 7792 19340 7812
rect 19340 7792 19392 7812
rect 19392 7792 19394 7812
rect 19154 6332 19156 6352
rect 19156 6332 19208 6352
rect 19208 6332 19210 6352
rect 19154 6296 19210 6332
rect 19246 5072 19302 5128
rect 19338 4936 19394 4992
rect 19154 3712 19210 3768
rect 18970 2624 19026 2680
rect 18602 2352 18658 2408
rect 19982 10648 20038 10704
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19706 9968 19762 10024
rect 19706 9696 19762 9752
rect 20350 15544 20406 15600
rect 20902 20440 20958 20496
rect 20902 20324 20958 20360
rect 20902 20304 20904 20324
rect 20904 20304 20956 20324
rect 20956 20304 20958 20324
rect 21178 20304 21234 20360
rect 21454 21528 21510 21584
rect 21178 19760 21234 19816
rect 20718 18420 20774 18456
rect 20718 18400 20720 18420
rect 20720 18400 20772 18420
rect 20772 18400 20774 18420
rect 20718 15580 20720 15600
rect 20720 15580 20772 15600
rect 20772 15580 20774 15600
rect 20718 15544 20774 15580
rect 20534 12416 20590 12472
rect 21362 18300 21364 18320
rect 21364 18300 21416 18320
rect 21416 18300 21418 18320
rect 21362 18264 21418 18300
rect 21822 22480 21878 22536
rect 21730 21800 21786 21856
rect 22190 20304 22246 20360
rect 21822 19488 21878 19544
rect 21086 16088 21142 16144
rect 20902 13232 20958 13288
rect 20810 12144 20866 12200
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 20258 9560 20314 9616
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 20166 8200 20222 8256
rect 20350 7928 20406 7984
rect 21086 10124 21142 10160
rect 21086 10104 21088 10124
rect 21088 10104 21140 10124
rect 21140 10104 21142 10124
rect 21086 9696 21142 9752
rect 20994 8336 21050 8392
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19614 6196 19616 6216
rect 19616 6196 19668 6216
rect 19668 6196 19670 6216
rect 19614 6160 19670 6196
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19982 5616 20038 5672
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19522 3440 19578 3496
rect 19890 3460 19946 3496
rect 19890 3440 19892 3460
rect 19892 3440 19944 3460
rect 19944 3440 19946 3460
rect 19430 2760 19486 2816
rect 18970 2080 19026 2136
rect 18694 1400 18750 1456
rect 20074 2760 20130 2816
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20902 5072 20958 5128
rect 21086 6432 21142 6488
rect 20810 4392 20866 4448
rect 20994 4392 21050 4448
rect 21362 14492 21364 14512
rect 21364 14492 21416 14512
rect 21416 14492 21418 14512
rect 21362 14456 21418 14492
rect 21730 15272 21786 15328
rect 22098 18672 22154 18728
rect 21822 15000 21878 15056
rect 21270 14320 21326 14376
rect 21362 13812 21364 13832
rect 21364 13812 21416 13832
rect 21416 13812 21418 13832
rect 21362 13776 21418 13812
rect 22282 17176 22338 17232
rect 22006 14864 22062 14920
rect 22466 24520 22522 24576
rect 23202 27104 23258 27160
rect 23662 26560 23718 26616
rect 24766 25880 24822 25936
rect 24766 25336 24822 25392
rect 23386 24248 23442 24304
rect 22650 21528 22706 21584
rect 22650 20984 22706 21040
rect 22650 19760 22706 19816
rect 22742 18964 22798 19000
rect 22742 18944 22744 18964
rect 22744 18944 22796 18964
rect 22796 18944 22798 18964
rect 22558 18128 22614 18184
rect 21454 10920 21510 10976
rect 21362 10804 21418 10840
rect 21362 10784 21364 10804
rect 21364 10784 21416 10804
rect 21416 10784 21418 10804
rect 21454 10240 21510 10296
rect 21362 9444 21418 9480
rect 21362 9424 21364 9444
rect 21364 9424 21416 9444
rect 21416 9424 21418 9444
rect 21730 10920 21786 10976
rect 21638 9832 21694 9888
rect 21362 8880 21418 8936
rect 21730 7656 21786 7712
rect 21730 7384 21786 7440
rect 21362 7248 21418 7304
rect 21270 6432 21326 6488
rect 21454 6704 21510 6760
rect 23110 20304 23166 20360
rect 23018 17448 23074 17504
rect 23202 19252 23204 19272
rect 23204 19252 23256 19272
rect 23256 19252 23258 19272
rect 23202 19216 23258 19252
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24122 24792 24178 24848
rect 23846 22888 23902 22944
rect 23294 17992 23350 18048
rect 22926 13776 22982 13832
rect 22006 10648 22062 10704
rect 22006 9968 22062 10024
rect 22190 9560 22246 9616
rect 21914 7792 21970 7848
rect 23202 13640 23258 13696
rect 23202 10784 23258 10840
rect 22006 6840 22062 6896
rect 21270 4256 21326 4312
rect 21178 3576 21234 3632
rect 20718 1808 20774 1864
rect 21638 4156 21640 4176
rect 21640 4156 21692 4176
rect 21692 4156 21694 4176
rect 21638 4120 21694 4156
rect 21914 2624 21970 2680
rect 22098 4528 22154 4584
rect 23018 9016 23074 9072
rect 23478 16360 23534 16416
rect 23662 22516 23664 22536
rect 23664 22516 23716 22536
rect 23716 22516 23718 22536
rect 23662 22480 23718 22516
rect 23662 17332 23718 17368
rect 23662 17312 23664 17332
rect 23664 17312 23716 17332
rect 23716 17312 23718 17332
rect 24030 19896 24086 19952
rect 23846 19216 23902 19272
rect 23846 17448 23902 17504
rect 23754 15272 23810 15328
rect 23938 14864 23994 14920
rect 23754 12416 23810 12472
rect 23386 10004 23388 10024
rect 23388 10004 23440 10024
rect 23440 10004 23442 10024
rect 23386 9968 23442 10004
rect 22650 7520 22706 7576
rect 23202 8200 23258 8256
rect 23110 7792 23166 7848
rect 22742 5208 22798 5264
rect 22834 4664 22890 4720
rect 22650 4120 22706 4176
rect 22374 3032 22430 3088
rect 23202 5208 23258 5264
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 23568 24822 23624
rect 25778 24112 25834 24168
rect 24674 23024 24730 23080
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 25502 23432 25558 23488
rect 24950 22616 25006 22672
rect 24766 22480 24822 22536
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 25042 21936 25098 21992
rect 24674 20712 24730 20768
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 25226 21428 25228 21448
rect 25228 21428 25280 21448
rect 25280 21428 25282 21448
rect 25226 21392 25282 21428
rect 25318 21256 25374 21312
rect 25134 20848 25190 20904
rect 24766 20032 24822 20088
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 25226 20440 25282 20496
rect 25318 19488 25374 19544
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24766 18264 24822 18320
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24214 17040 24270 17096
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 25226 19352 25282 19408
rect 25410 18400 25466 18456
rect 24766 16632 24822 16688
rect 24766 15952 24822 16008
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24214 14320 24270 14376
rect 24122 12552 24178 12608
rect 24030 11736 24086 11792
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 25042 17992 25098 18048
rect 25226 17720 25282 17776
rect 25226 17584 25282 17640
rect 25410 17176 25466 17232
rect 25410 16108 25466 16144
rect 25410 16088 25412 16108
rect 25412 16088 25464 16108
rect 25464 16088 25466 16108
rect 25134 13368 25190 13424
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24214 12280 24270 12336
rect 24582 12144 24638 12200
rect 23938 11600 23994 11656
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24306 11600 24362 11656
rect 24306 11056 24362 11112
rect 23846 9832 23902 9888
rect 23570 8880 23626 8936
rect 23662 8472 23718 8528
rect 23662 8064 23718 8120
rect 23662 6452 23718 6488
rect 23662 6432 23664 6452
rect 23664 6432 23716 6452
rect 23716 6432 23718 6452
rect 23846 7112 23902 7168
rect 23754 5616 23810 5672
rect 23570 4392 23626 4448
rect 23478 3712 23534 3768
rect 23846 2896 23902 2952
rect 23754 1672 23810 1728
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24674 7656 24730 7712
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24122 6840 24178 6896
rect 24214 6724 24270 6760
rect 24214 6704 24216 6724
rect 24216 6704 24268 6724
rect 24268 6704 24270 6724
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24766 7384 24822 7440
rect 25686 13096 25742 13152
rect 25134 9968 25190 10024
rect 25042 9052 25044 9072
rect 25044 9052 25096 9072
rect 25096 9052 25098 9072
rect 25042 9016 25098 9052
rect 25594 11756 25650 11792
rect 25594 11736 25596 11756
rect 25596 11736 25648 11756
rect 25648 11736 25650 11756
rect 27526 20984 27582 21040
rect 26146 19760 26202 19816
rect 25410 7656 25466 7712
rect 25226 7284 25228 7304
rect 25228 7284 25280 7304
rect 25280 7284 25282 7304
rect 25226 7248 25282 7284
rect 25042 6840 25098 6896
rect 24766 6704 24822 6760
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 25226 5208 25282 5264
rect 24674 3576 24730 3632
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24122 3032 24178 3088
rect 24582 2896 24638 2952
rect 24490 2624 24546 2680
rect 24766 2760 24822 2816
rect 24674 2624 24730 2680
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25502 5752 25558 5808
rect 25686 4936 25742 4992
rect 25594 4392 25650 4448
rect 26146 4120 26202 4176
rect 25410 3440 25466 3496
rect 25226 2488 25282 2544
rect 25502 1536 25558 1592
rect 27526 3440 27582 3496
rect 23938 312 23994 368
<< metal3 >>
rect 23105 27706 23171 27709
rect 27520 27706 28000 27736
rect 23105 27704 28000 27706
rect 23105 27648 23110 27704
rect 23166 27648 28000 27704
rect 23105 27646 28000 27648
rect 23105 27643 23171 27646
rect 27520 27616 28000 27646
rect 23197 27162 23263 27165
rect 27520 27162 28000 27192
rect 23197 27160 28000 27162
rect 23197 27104 23202 27160
rect 23258 27104 28000 27160
rect 23197 27102 28000 27104
rect 23197 27099 23263 27102
rect 27520 27072 28000 27102
rect 23657 26618 23723 26621
rect 27520 26618 28000 26648
rect 23657 26616 28000 26618
rect 23657 26560 23662 26616
rect 23718 26560 28000 26616
rect 23657 26558 28000 26560
rect 23657 26555 23723 26558
rect 27520 26528 28000 26558
rect 24761 25938 24827 25941
rect 27520 25938 28000 25968
rect 24761 25936 28000 25938
rect 24761 25880 24766 25936
rect 24822 25880 28000 25936
rect 24761 25878 28000 25880
rect 24761 25875 24827 25878
rect 27520 25848 28000 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 24761 25394 24827 25397
rect 27520 25394 28000 25424
rect 24761 25392 28000 25394
rect 24761 25336 24766 25392
rect 24822 25336 28000 25392
rect 24761 25334 28000 25336
rect 24761 25331 24827 25334
rect 27520 25304 28000 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 9121 24850 9187 24853
rect 14181 24850 14247 24853
rect 9121 24848 14247 24850
rect 9121 24792 9126 24848
rect 9182 24792 14186 24848
rect 14242 24792 14247 24848
rect 9121 24790 14247 24792
rect 9121 24787 9187 24790
rect 14181 24787 14247 24790
rect 14365 24850 14431 24853
rect 15929 24850 15995 24853
rect 14365 24848 15995 24850
rect 14365 24792 14370 24848
rect 14426 24792 15934 24848
rect 15990 24792 15995 24848
rect 14365 24790 15995 24792
rect 14365 24787 14431 24790
rect 15929 24787 15995 24790
rect 24117 24850 24183 24853
rect 27520 24850 28000 24880
rect 24117 24848 28000 24850
rect 24117 24792 24122 24848
rect 24178 24792 28000 24848
rect 24117 24790 28000 24792
rect 24117 24787 24183 24790
rect 27520 24760 28000 24790
rect 6361 24714 6427 24717
rect 9673 24714 9739 24717
rect 6361 24712 9739 24714
rect 6361 24656 6366 24712
rect 6422 24656 9678 24712
rect 9734 24656 9739 24712
rect 6361 24654 9739 24656
rect 6361 24651 6427 24654
rect 9673 24651 9739 24654
rect 12801 24714 12867 24717
rect 14549 24714 14615 24717
rect 20253 24714 20319 24717
rect 12801 24712 14615 24714
rect 12801 24656 12806 24712
rect 12862 24656 14554 24712
rect 14610 24656 14615 24712
rect 12801 24654 14615 24656
rect 12801 24651 12867 24654
rect 14549 24651 14615 24654
rect 19382 24712 20319 24714
rect 19382 24656 20258 24712
rect 20314 24656 20319 24712
rect 19382 24654 20319 24656
rect 11329 24578 11395 24581
rect 19382 24578 19442 24654
rect 20253 24651 20319 24654
rect 11329 24576 19442 24578
rect 11329 24520 11334 24576
rect 11390 24520 19442 24576
rect 11329 24518 19442 24520
rect 20069 24578 20135 24581
rect 22461 24578 22527 24581
rect 20069 24576 22527 24578
rect 20069 24520 20074 24576
rect 20130 24520 22466 24576
rect 22522 24520 22527 24576
rect 20069 24518 22527 24520
rect 11329 24515 11395 24518
rect 20069 24515 20135 24518
rect 22461 24515 22527 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 11881 24442 11947 24445
rect 13721 24442 13787 24445
rect 17953 24442 18019 24445
rect 11881 24440 13554 24442
rect 11881 24384 11886 24440
rect 11942 24384 13554 24440
rect 11881 24382 13554 24384
rect 11881 24379 11947 24382
rect 4337 24306 4403 24309
rect 12157 24306 12223 24309
rect 4337 24304 12223 24306
rect 4337 24248 4342 24304
rect 4398 24248 12162 24304
rect 12218 24248 12223 24304
rect 4337 24246 12223 24248
rect 13494 24306 13554 24382
rect 13721 24440 18019 24442
rect 13721 24384 13726 24440
rect 13782 24384 17958 24440
rect 18014 24384 18019 24440
rect 13721 24382 18019 24384
rect 13721 24379 13787 24382
rect 17953 24379 18019 24382
rect 23381 24306 23447 24309
rect 13494 24304 23447 24306
rect 13494 24248 23386 24304
rect 23442 24248 23447 24304
rect 13494 24246 23447 24248
rect 4337 24243 4403 24246
rect 12157 24243 12223 24246
rect 23381 24243 23447 24246
rect 933 24170 999 24173
rect 14273 24170 14339 24173
rect 933 24168 14339 24170
rect 933 24112 938 24168
rect 994 24112 14278 24168
rect 14334 24112 14339 24168
rect 933 24110 14339 24112
rect 933 24107 999 24110
rect 14273 24107 14339 24110
rect 18965 24170 19031 24173
rect 19977 24170 20043 24173
rect 18965 24168 20043 24170
rect 18965 24112 18970 24168
rect 19026 24112 19982 24168
rect 20038 24112 20043 24168
rect 18965 24110 20043 24112
rect 18965 24107 19031 24110
rect 19977 24107 20043 24110
rect 25773 24170 25839 24173
rect 27520 24170 28000 24200
rect 25773 24168 28000 24170
rect 25773 24112 25778 24168
rect 25834 24112 28000 24168
rect 25773 24110 28000 24112
rect 25773 24107 25839 24110
rect 27520 24080 28000 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 9765 23626 9831 23629
rect 13721 23626 13787 23629
rect 9765 23624 13787 23626
rect 9765 23568 9770 23624
rect 9826 23568 13726 23624
rect 13782 23568 13787 23624
rect 9765 23566 13787 23568
rect 9765 23563 9831 23566
rect 13721 23563 13787 23566
rect 24761 23626 24827 23629
rect 27520 23626 28000 23656
rect 24761 23624 28000 23626
rect 24761 23568 24766 23624
rect 24822 23568 28000 23624
rect 24761 23566 28000 23568
rect 24761 23563 24827 23566
rect 27520 23536 28000 23566
rect 21633 23490 21699 23493
rect 25497 23490 25563 23493
rect 21633 23488 25563 23490
rect 21633 23432 21638 23488
rect 21694 23432 25502 23488
rect 25558 23432 25563 23488
rect 21633 23430 25563 23432
rect 21633 23427 21699 23430
rect 25497 23427 25563 23430
rect 10277 23424 10597 23425
rect 0 23354 480 23384
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 4981 23354 5047 23357
rect 9581 23354 9647 23357
rect 0 23294 1226 23354
rect 0 23264 480 23294
rect 1166 22130 1226 23294
rect 4981 23352 9647 23354
rect 4981 23296 4986 23352
rect 5042 23296 9586 23352
rect 9642 23296 9647 23352
rect 4981 23294 9647 23296
rect 4981 23291 5047 23294
rect 9581 23291 9647 23294
rect 12525 23354 12591 23357
rect 14365 23354 14431 23357
rect 12525 23352 14431 23354
rect 12525 23296 12530 23352
rect 12586 23296 14370 23352
rect 14426 23296 14431 23352
rect 12525 23294 14431 23296
rect 12525 23291 12591 23294
rect 14365 23291 14431 23294
rect 15285 23354 15351 23357
rect 19149 23354 19215 23357
rect 15285 23352 19215 23354
rect 15285 23296 15290 23352
rect 15346 23296 19154 23352
rect 19210 23296 19215 23352
rect 15285 23294 19215 23296
rect 15285 23291 15351 23294
rect 19149 23291 19215 23294
rect 13721 23082 13787 23085
rect 19885 23082 19951 23085
rect 13721 23080 19951 23082
rect 13721 23024 13726 23080
rect 13782 23024 19890 23080
rect 19946 23024 19951 23080
rect 13721 23022 19951 23024
rect 13721 23019 13787 23022
rect 19885 23019 19951 23022
rect 24669 23082 24735 23085
rect 27520 23082 28000 23112
rect 24669 23080 28000 23082
rect 24669 23024 24674 23080
rect 24730 23024 28000 23080
rect 24669 23022 28000 23024
rect 24669 23019 24735 23022
rect 27520 22992 28000 23022
rect 10777 22946 10843 22949
rect 12709 22946 12775 22949
rect 10777 22944 12775 22946
rect 10777 22888 10782 22944
rect 10838 22888 12714 22944
rect 12770 22888 12775 22944
rect 10777 22886 12775 22888
rect 10777 22883 10843 22886
rect 12709 22883 12775 22886
rect 16113 22946 16179 22949
rect 23841 22946 23907 22949
rect 16113 22944 23907 22946
rect 16113 22888 16118 22944
rect 16174 22888 23846 22944
rect 23902 22888 23907 22944
rect 16113 22886 23907 22888
rect 16113 22883 16179 22886
rect 23841 22883 23907 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 7741 22810 7807 22813
rect 10593 22810 10659 22813
rect 7741 22808 10659 22810
rect 7741 22752 7746 22808
rect 7802 22752 10598 22808
rect 10654 22752 10659 22808
rect 7741 22750 10659 22752
rect 7741 22747 7807 22750
rect 10593 22747 10659 22750
rect 10869 22810 10935 22813
rect 14089 22810 14155 22813
rect 10869 22808 14155 22810
rect 10869 22752 10874 22808
rect 10930 22752 14094 22808
rect 14150 22752 14155 22808
rect 10869 22750 14155 22752
rect 10869 22747 10935 22750
rect 14089 22747 14155 22750
rect 15929 22810 15995 22813
rect 20161 22810 20227 22813
rect 20989 22810 21055 22813
rect 15929 22808 21055 22810
rect 15929 22752 15934 22808
rect 15990 22752 20166 22808
rect 20222 22752 20994 22808
rect 21050 22752 21055 22808
rect 15929 22750 21055 22752
rect 15929 22747 15995 22750
rect 20161 22747 20227 22750
rect 20989 22747 21055 22750
rect 1577 22674 1643 22677
rect 13353 22674 13419 22677
rect 1577 22672 13419 22674
rect 1577 22616 1582 22672
rect 1638 22616 13358 22672
rect 13414 22616 13419 22672
rect 1577 22614 13419 22616
rect 1577 22611 1643 22614
rect 13353 22611 13419 22614
rect 19793 22674 19859 22677
rect 24945 22674 25011 22677
rect 19793 22672 25011 22674
rect 19793 22616 19798 22672
rect 19854 22616 24950 22672
rect 25006 22616 25011 22672
rect 19793 22614 25011 22616
rect 19793 22611 19859 22614
rect 24945 22611 25011 22614
rect 12249 22538 12315 22541
rect 20805 22538 20871 22541
rect 12249 22536 20871 22538
rect 12249 22480 12254 22536
rect 12310 22480 20810 22536
rect 20866 22480 20871 22536
rect 12249 22478 20871 22480
rect 12249 22475 12315 22478
rect 20805 22475 20871 22478
rect 21817 22538 21883 22541
rect 23657 22538 23723 22541
rect 21817 22536 23723 22538
rect 21817 22480 21822 22536
rect 21878 22480 23662 22536
rect 23718 22480 23723 22536
rect 21817 22478 23723 22480
rect 21817 22475 21883 22478
rect 23657 22475 23723 22478
rect 24761 22538 24827 22541
rect 27520 22538 28000 22568
rect 24761 22536 28000 22538
rect 24761 22480 24766 22536
rect 24822 22480 28000 22536
rect 24761 22478 28000 22480
rect 24761 22475 24827 22478
rect 27520 22448 28000 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 20437 22130 20503 22133
rect 1166 22128 20503 22130
rect 1166 22072 20442 22128
rect 20498 22072 20503 22128
rect 1166 22070 20503 22072
rect 20437 22067 20503 22070
rect 9581 21994 9647 21997
rect 14733 21994 14799 21997
rect 9581 21992 14799 21994
rect 9581 21936 9586 21992
rect 9642 21936 14738 21992
rect 14794 21936 14799 21992
rect 9581 21934 14799 21936
rect 9581 21931 9647 21934
rect 14733 21931 14799 21934
rect 15561 21994 15627 21997
rect 25037 21994 25103 21997
rect 15561 21992 25103 21994
rect 15561 21936 15566 21992
rect 15622 21936 25042 21992
rect 25098 21936 25103 21992
rect 15561 21934 25103 21936
rect 15561 21931 15627 21934
rect 25037 21931 25103 21934
rect 21725 21858 21791 21861
rect 27520 21858 28000 21888
rect 21590 21856 21791 21858
rect 21590 21800 21730 21856
rect 21786 21800 21791 21856
rect 21590 21798 21791 21800
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 10133 21722 10199 21725
rect 12709 21722 12775 21725
rect 10133 21720 12775 21722
rect 10133 21664 10138 21720
rect 10194 21664 12714 21720
rect 12770 21664 12775 21720
rect 10133 21662 12775 21664
rect 10133 21659 10199 21662
rect 12709 21659 12775 21662
rect 11145 21586 11211 21589
rect 21449 21586 21515 21589
rect 21590 21586 21650 21798
rect 21725 21795 21791 21798
rect 24764 21798 28000 21858
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 11145 21584 21650 21586
rect 11145 21528 11150 21584
rect 11206 21528 21454 21584
rect 21510 21528 21650 21584
rect 11145 21526 21650 21528
rect 22645 21586 22711 21589
rect 24764 21586 24824 21798
rect 27520 21768 28000 21798
rect 22645 21584 24824 21586
rect 22645 21528 22650 21584
rect 22706 21528 24824 21584
rect 22645 21526 24824 21528
rect 11145 21523 11211 21526
rect 21449 21523 21515 21526
rect 22645 21523 22711 21526
rect 2957 21450 3023 21453
rect 14641 21450 14707 21453
rect 2957 21448 14707 21450
rect 2957 21392 2962 21448
rect 3018 21392 14646 21448
rect 14702 21392 14707 21448
rect 2957 21390 14707 21392
rect 2957 21387 3023 21390
rect 14641 21387 14707 21390
rect 19241 21450 19307 21453
rect 25221 21450 25287 21453
rect 19241 21448 25287 21450
rect 19241 21392 19246 21448
rect 19302 21392 25226 21448
rect 25282 21392 25287 21448
rect 19241 21390 25287 21392
rect 19241 21387 19307 21390
rect 25221 21387 25287 21390
rect 25313 21314 25379 21317
rect 27520 21314 28000 21344
rect 25313 21312 28000 21314
rect 25313 21256 25318 21312
rect 25374 21256 28000 21312
rect 25313 21254 28000 21256
rect 25313 21251 25379 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 27520 21224 28000 21254
rect 19610 21183 19930 21184
rect 22645 21042 22711 21045
rect 27521 21042 27587 21045
rect 22645 21040 27587 21042
rect 22645 20984 22650 21040
rect 22706 20984 27526 21040
rect 27582 20984 27587 21040
rect 22645 20982 27587 20984
rect 22645 20979 22711 20982
rect 27521 20979 27587 20982
rect 9673 20906 9739 20909
rect 11513 20906 11579 20909
rect 25129 20906 25195 20909
rect 9673 20904 9874 20906
rect 9673 20848 9678 20904
rect 9734 20848 9874 20904
rect 9673 20846 9874 20848
rect 9673 20843 9739 20846
rect 9814 20770 9874 20846
rect 11513 20904 25195 20906
rect 11513 20848 11518 20904
rect 11574 20848 25134 20904
rect 25190 20848 25195 20904
rect 11513 20846 25195 20848
rect 11513 20843 11579 20846
rect 25129 20843 25195 20846
rect 9949 20770 10015 20773
rect 9814 20768 10015 20770
rect 9814 20712 9954 20768
rect 10010 20712 10015 20768
rect 9814 20710 10015 20712
rect 9949 20707 10015 20710
rect 24669 20770 24735 20773
rect 27520 20770 28000 20800
rect 24669 20768 28000 20770
rect 24669 20712 24674 20768
rect 24730 20712 28000 20768
rect 24669 20710 28000 20712
rect 24669 20707 24735 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 27520 20680 28000 20710
rect 24277 20639 24597 20640
rect 10961 20634 11027 20637
rect 10961 20632 14842 20634
rect 10961 20576 10966 20632
rect 11022 20576 14842 20632
rect 10961 20574 14842 20576
rect 10961 20571 11027 20574
rect 3693 20498 3759 20501
rect 13997 20498 14063 20501
rect 3693 20496 14063 20498
rect 3693 20440 3698 20496
rect 3754 20440 14002 20496
rect 14058 20440 14063 20496
rect 3693 20438 14063 20440
rect 14782 20498 14842 20574
rect 15653 20498 15719 20501
rect 20897 20498 20963 20501
rect 25221 20498 25287 20501
rect 14782 20496 17602 20498
rect 14782 20440 15658 20496
rect 15714 20440 17602 20496
rect 14782 20438 17602 20440
rect 3693 20435 3759 20438
rect 13997 20435 14063 20438
rect 15653 20435 15719 20438
rect 12341 20362 12407 20365
rect 17125 20362 17191 20365
rect 12341 20360 17191 20362
rect 12341 20304 12346 20360
rect 12402 20304 17130 20360
rect 17186 20304 17191 20360
rect 12341 20302 17191 20304
rect 17542 20362 17602 20438
rect 20897 20496 25287 20498
rect 20897 20440 20902 20496
rect 20958 20440 25226 20496
rect 25282 20440 25287 20496
rect 20897 20438 25287 20440
rect 20897 20435 20963 20438
rect 25221 20435 25287 20438
rect 20897 20362 20963 20365
rect 17542 20360 20963 20362
rect 17542 20304 20902 20360
rect 20958 20304 20963 20360
rect 17542 20302 20963 20304
rect 12341 20299 12407 20302
rect 17125 20299 17191 20302
rect 20897 20299 20963 20302
rect 21173 20362 21239 20365
rect 22185 20362 22251 20365
rect 23105 20362 23171 20365
rect 21173 20360 23171 20362
rect 21173 20304 21178 20360
rect 21234 20304 22190 20360
rect 22246 20304 23110 20360
rect 23166 20304 23171 20360
rect 21173 20302 23171 20304
rect 21173 20299 21239 20302
rect 22185 20299 22251 20302
rect 23105 20299 23171 20302
rect 12525 20226 12591 20229
rect 17677 20226 17743 20229
rect 12525 20224 17743 20226
rect 12525 20168 12530 20224
rect 12586 20168 17682 20224
rect 17738 20168 17743 20224
rect 12525 20166 17743 20168
rect 12525 20163 12591 20166
rect 17677 20163 17743 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 10869 20090 10935 20093
rect 13813 20090 13879 20093
rect 10869 20088 13879 20090
rect 10869 20032 10874 20088
rect 10930 20032 13818 20088
rect 13874 20032 13879 20088
rect 10869 20030 13879 20032
rect 10869 20027 10935 20030
rect 13813 20027 13879 20030
rect 24761 20090 24827 20093
rect 27520 20090 28000 20120
rect 24761 20088 28000 20090
rect 24761 20032 24766 20088
rect 24822 20032 28000 20088
rect 24761 20030 28000 20032
rect 24761 20027 24827 20030
rect 27520 20000 28000 20030
rect 12617 19954 12683 19957
rect 19793 19954 19859 19957
rect 24025 19954 24091 19957
rect 12617 19952 19626 19954
rect 12617 19896 12622 19952
rect 12678 19896 19626 19952
rect 12617 19894 19626 19896
rect 12617 19891 12683 19894
rect 14273 19818 14339 19821
rect 15469 19818 15535 19821
rect 14273 19816 15535 19818
rect 14273 19760 14278 19816
rect 14334 19760 15474 19816
rect 15530 19760 15535 19816
rect 14273 19758 15535 19760
rect 19566 19818 19626 19894
rect 19793 19952 24091 19954
rect 19793 19896 19798 19952
rect 19854 19896 24030 19952
rect 24086 19896 24091 19952
rect 19793 19894 24091 19896
rect 19793 19891 19859 19894
rect 24025 19891 24091 19894
rect 21173 19818 21239 19821
rect 19566 19816 21239 19818
rect 19566 19760 21178 19816
rect 21234 19760 21239 19816
rect 19566 19758 21239 19760
rect 14273 19755 14339 19758
rect 15469 19755 15535 19758
rect 21173 19755 21239 19758
rect 22645 19818 22711 19821
rect 26141 19818 26207 19821
rect 22645 19816 26207 19818
rect 22645 19760 22650 19816
rect 22706 19760 26146 19816
rect 26202 19760 26207 19816
rect 22645 19758 26207 19760
rect 22645 19755 22711 19758
rect 26141 19755 26207 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 18965 19546 19031 19549
rect 21817 19546 21883 19549
rect 18965 19544 21883 19546
rect 18965 19488 18970 19544
rect 19026 19488 21822 19544
rect 21878 19488 21883 19544
rect 18965 19486 21883 19488
rect 18965 19483 19031 19486
rect 21817 19483 21883 19486
rect 25313 19546 25379 19549
rect 27520 19546 28000 19576
rect 25313 19544 28000 19546
rect 25313 19488 25318 19544
rect 25374 19488 28000 19544
rect 25313 19486 28000 19488
rect 25313 19483 25379 19486
rect 27520 19456 28000 19486
rect 9581 19410 9647 19413
rect 13353 19410 13419 19413
rect 14733 19410 14799 19413
rect 15745 19410 15811 19413
rect 9500 19408 9690 19410
rect 9500 19352 9586 19408
rect 9642 19352 9690 19408
rect 9500 19350 9690 19352
rect 9581 19347 9690 19350
rect 13353 19408 15811 19410
rect 13353 19352 13358 19408
rect 13414 19352 14738 19408
rect 14794 19352 15750 19408
rect 15806 19352 15811 19408
rect 13353 19350 15811 19352
rect 13353 19347 13419 19350
rect 14733 19347 14799 19350
rect 15745 19347 15811 19350
rect 19609 19410 19675 19413
rect 25221 19410 25287 19413
rect 19609 19408 25287 19410
rect 19609 19352 19614 19408
rect 19670 19352 25226 19408
rect 25282 19352 25287 19408
rect 19609 19350 25287 19352
rect 19609 19347 19675 19350
rect 25221 19347 25287 19350
rect 9630 19274 9690 19347
rect 9765 19274 9831 19277
rect 9630 19272 9831 19274
rect 9630 19216 9770 19272
rect 9826 19216 9831 19272
rect 9630 19214 9831 19216
rect 9765 19211 9831 19214
rect 14825 19274 14891 19277
rect 16757 19274 16823 19277
rect 14825 19272 16823 19274
rect 14825 19216 14830 19272
rect 14886 19216 16762 19272
rect 16818 19216 16823 19272
rect 14825 19214 16823 19216
rect 14825 19211 14891 19214
rect 16757 19211 16823 19214
rect 23197 19274 23263 19277
rect 23841 19274 23907 19277
rect 23197 19272 23907 19274
rect 23197 19216 23202 19272
rect 23258 19216 23846 19272
rect 23902 19216 23907 19272
rect 23197 19214 23907 19216
rect 23197 19211 23263 19214
rect 23841 19211 23907 19214
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 22737 19002 22803 19005
rect 27520 19002 28000 19032
rect 22737 19000 28000 19002
rect 22737 18944 22742 19000
rect 22798 18944 28000 19000
rect 22737 18942 28000 18944
rect 22737 18939 22803 18942
rect 27520 18912 28000 18942
rect 9489 18866 9555 18869
rect 14825 18866 14891 18869
rect 9489 18864 14891 18866
rect 9489 18808 9494 18864
rect 9550 18808 14830 18864
rect 14886 18808 14891 18864
rect 9489 18806 14891 18808
rect 9489 18803 9555 18806
rect 14825 18803 14891 18806
rect 15285 18730 15351 18733
rect 22093 18730 22159 18733
rect 15285 18728 22159 18730
rect 15285 18672 15290 18728
rect 15346 18672 22098 18728
rect 22154 18672 22159 18728
rect 15285 18670 22159 18672
rect 15285 18667 15351 18670
rect 22093 18667 22159 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 19241 18458 19307 18461
rect 20713 18458 20779 18461
rect 19241 18456 20779 18458
rect 19241 18400 19246 18456
rect 19302 18400 20718 18456
rect 20774 18400 20779 18456
rect 19241 18398 20779 18400
rect 19241 18395 19307 18398
rect 20713 18395 20779 18398
rect 25405 18458 25471 18461
rect 27520 18458 28000 18488
rect 25405 18456 28000 18458
rect 25405 18400 25410 18456
rect 25466 18400 28000 18456
rect 25405 18398 28000 18400
rect 25405 18395 25471 18398
rect 27520 18368 28000 18398
rect 10133 18322 10199 18325
rect 12433 18322 12499 18325
rect 10133 18320 12499 18322
rect 10133 18264 10138 18320
rect 10194 18264 12438 18320
rect 12494 18264 12499 18320
rect 10133 18262 12499 18264
rect 10133 18259 10199 18262
rect 12433 18259 12499 18262
rect 14457 18322 14523 18325
rect 18873 18322 18939 18325
rect 14457 18320 18939 18322
rect 14457 18264 14462 18320
rect 14518 18264 18878 18320
rect 18934 18264 18939 18320
rect 14457 18262 18939 18264
rect 14457 18259 14523 18262
rect 18873 18259 18939 18262
rect 21357 18322 21423 18325
rect 24761 18322 24827 18325
rect 21357 18320 24827 18322
rect 21357 18264 21362 18320
rect 21418 18264 24766 18320
rect 24822 18264 24827 18320
rect 21357 18262 24827 18264
rect 21357 18259 21423 18262
rect 24761 18259 24827 18262
rect 12709 18186 12775 18189
rect 22553 18186 22619 18189
rect 12709 18184 22619 18186
rect 12709 18128 12714 18184
rect 12770 18128 22558 18184
rect 22614 18128 22619 18184
rect 12709 18126 22619 18128
rect 12709 18123 12775 18126
rect 22553 18123 22619 18126
rect 14825 18050 14891 18053
rect 18781 18050 18847 18053
rect 14825 18048 18847 18050
rect 14825 17992 14830 18048
rect 14886 17992 18786 18048
rect 18842 17992 18847 18048
rect 14825 17990 18847 17992
rect 14825 17987 14891 17990
rect 18781 17987 18847 17990
rect 23289 18050 23355 18053
rect 25037 18050 25103 18053
rect 23289 18048 25103 18050
rect 23289 17992 23294 18048
rect 23350 17992 25042 18048
rect 25098 17992 25103 18048
rect 23289 17990 25103 17992
rect 23289 17987 23355 17990
rect 25037 17987 25103 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 5993 17914 6059 17917
rect 10133 17914 10199 17917
rect 5993 17912 10199 17914
rect 5993 17856 5998 17912
rect 6054 17856 10138 17912
rect 10194 17856 10199 17912
rect 5993 17854 10199 17856
rect 5993 17851 6059 17854
rect 10133 17851 10199 17854
rect 12065 17914 12131 17917
rect 13813 17914 13879 17917
rect 12065 17912 13879 17914
rect 12065 17856 12070 17912
rect 12126 17856 13818 17912
rect 13874 17856 13879 17912
rect 12065 17854 13879 17856
rect 12065 17851 12131 17854
rect 13813 17851 13879 17854
rect 25221 17778 25287 17781
rect 27520 17778 28000 17808
rect 25221 17776 28000 17778
rect 25221 17720 25226 17776
rect 25282 17720 28000 17776
rect 25221 17718 28000 17720
rect 25221 17715 25287 17718
rect 27520 17688 28000 17718
rect 11329 17642 11395 17645
rect 16021 17642 16087 17645
rect 11329 17640 16087 17642
rect 11329 17584 11334 17640
rect 11390 17584 16026 17640
rect 16082 17584 16087 17640
rect 11329 17582 16087 17584
rect 11329 17579 11395 17582
rect 16021 17579 16087 17582
rect 17217 17642 17283 17645
rect 25221 17642 25287 17645
rect 17217 17640 25287 17642
rect 17217 17584 17222 17640
rect 17278 17584 25226 17640
rect 25282 17584 25287 17640
rect 17217 17582 25287 17584
rect 17217 17579 17283 17582
rect 25221 17579 25287 17582
rect 18597 17506 18663 17509
rect 23013 17506 23079 17509
rect 23841 17506 23907 17509
rect 18597 17504 23907 17506
rect 18597 17448 18602 17504
rect 18658 17448 23018 17504
rect 23074 17448 23846 17504
rect 23902 17448 23907 17504
rect 18597 17446 23907 17448
rect 18597 17443 18663 17446
rect 23013 17443 23079 17446
rect 23841 17443 23907 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 19977 17370 20043 17373
rect 20161 17370 20227 17373
rect 23657 17370 23723 17373
rect 19977 17368 23723 17370
rect 19977 17312 19982 17368
rect 20038 17312 20166 17368
rect 20222 17312 23662 17368
rect 23718 17312 23723 17368
rect 19977 17310 23723 17312
rect 19977 17307 20043 17310
rect 20161 17307 20227 17310
rect 23657 17307 23723 17310
rect 10777 17234 10843 17237
rect 11789 17234 11855 17237
rect 10777 17232 11855 17234
rect 10777 17176 10782 17232
rect 10838 17176 11794 17232
rect 11850 17176 11855 17232
rect 10777 17174 11855 17176
rect 10777 17171 10843 17174
rect 11789 17171 11855 17174
rect 18873 17234 18939 17237
rect 22277 17234 22343 17237
rect 18873 17232 22343 17234
rect 18873 17176 18878 17232
rect 18934 17176 22282 17232
rect 22338 17176 22343 17232
rect 18873 17174 22343 17176
rect 18873 17171 18939 17174
rect 22277 17171 22343 17174
rect 25405 17234 25471 17237
rect 27520 17234 28000 17264
rect 25405 17232 28000 17234
rect 25405 17176 25410 17232
rect 25466 17176 28000 17232
rect 25405 17174 28000 17176
rect 25405 17171 25471 17174
rect 27520 17144 28000 17174
rect 13169 17098 13235 17101
rect 24209 17098 24275 17101
rect 13169 17096 24275 17098
rect 13169 17040 13174 17096
rect 13230 17040 24214 17096
rect 24270 17040 24275 17096
rect 13169 17038 24275 17040
rect 13169 17035 13235 17038
rect 24209 17035 24275 17038
rect 13445 16962 13511 16965
rect 19241 16962 19307 16965
rect 13445 16960 19307 16962
rect 13445 16904 13450 16960
rect 13506 16904 19246 16960
rect 19302 16904 19307 16960
rect 13445 16902 19307 16904
rect 13445 16899 13511 16902
rect 19241 16899 19307 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 14549 16690 14615 16693
rect 16389 16690 16455 16693
rect 19149 16690 19215 16693
rect 14549 16688 16314 16690
rect 14549 16632 14554 16688
rect 14610 16632 16314 16688
rect 14549 16630 16314 16632
rect 14549 16627 14615 16630
rect 14089 16554 14155 16557
rect 16254 16554 16314 16630
rect 16389 16688 19215 16690
rect 16389 16632 16394 16688
rect 16450 16632 19154 16688
rect 19210 16632 19215 16688
rect 16389 16630 19215 16632
rect 16389 16627 16455 16630
rect 19149 16627 19215 16630
rect 24761 16690 24827 16693
rect 27520 16690 28000 16720
rect 24761 16688 28000 16690
rect 24761 16632 24766 16688
rect 24822 16632 28000 16688
rect 24761 16630 28000 16632
rect 24761 16627 24827 16630
rect 27520 16600 28000 16630
rect 16849 16554 16915 16557
rect 14089 16552 16130 16554
rect 14089 16496 14094 16552
rect 14150 16496 16130 16552
rect 14089 16494 16130 16496
rect 16254 16552 16915 16554
rect 16254 16496 16854 16552
rect 16910 16496 16915 16552
rect 16254 16494 16915 16496
rect 14089 16491 14155 16494
rect 16070 16418 16130 16494
rect 16849 16491 16915 16494
rect 20069 16418 20135 16421
rect 23473 16418 23539 16421
rect 16070 16416 23539 16418
rect 16070 16360 20074 16416
rect 20130 16360 23478 16416
rect 23534 16360 23539 16416
rect 16070 16358 23539 16360
rect 20069 16355 20135 16358
rect 23473 16355 23539 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 11881 16282 11947 16285
rect 14181 16282 14247 16285
rect 11881 16280 14247 16282
rect 11881 16224 11886 16280
rect 11942 16224 14186 16280
rect 14242 16224 14247 16280
rect 11881 16222 14247 16224
rect 11881 16219 11947 16222
rect 14181 16219 14247 16222
rect 21081 16146 21147 16149
rect 25405 16146 25471 16149
rect 21081 16144 25471 16146
rect 21081 16088 21086 16144
rect 21142 16088 25410 16144
rect 25466 16088 25471 16144
rect 21081 16086 25471 16088
rect 21081 16083 21147 16086
rect 25405 16083 25471 16086
rect 8293 16010 8359 16013
rect 18045 16010 18111 16013
rect 8293 16008 18111 16010
rect 8293 15952 8298 16008
rect 8354 15952 18050 16008
rect 18106 15952 18111 16008
rect 8293 15950 18111 15952
rect 8293 15947 8359 15950
rect 18045 15947 18111 15950
rect 24761 16010 24827 16013
rect 27520 16010 28000 16040
rect 24761 16008 28000 16010
rect 24761 15952 24766 16008
rect 24822 15952 28000 16008
rect 24761 15950 28000 15952
rect 24761 15947 24827 15950
rect 27520 15920 28000 15950
rect 16297 15874 16363 15877
rect 18321 15874 18387 15877
rect 16297 15872 18387 15874
rect 16297 15816 16302 15872
rect 16358 15816 18326 15872
rect 18382 15816 18387 15872
rect 16297 15814 18387 15816
rect 16297 15811 16363 15814
rect 18321 15811 18387 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 12065 15738 12131 15741
rect 15469 15738 15535 15741
rect 16665 15738 16731 15741
rect 12065 15736 16731 15738
rect 12065 15680 12070 15736
rect 12126 15680 15474 15736
rect 15530 15680 16670 15736
rect 16726 15680 16731 15736
rect 12065 15678 16731 15680
rect 12065 15675 12131 15678
rect 15469 15675 15535 15678
rect 16665 15675 16731 15678
rect 13721 15602 13787 15605
rect 15469 15602 15535 15605
rect 13721 15600 15535 15602
rect 13721 15544 13726 15600
rect 13782 15544 15474 15600
rect 15530 15544 15535 15600
rect 13721 15542 15535 15544
rect 13721 15539 13787 15542
rect 15469 15539 15535 15542
rect 17677 15602 17743 15605
rect 20345 15602 20411 15605
rect 20713 15602 20779 15605
rect 17677 15600 20779 15602
rect 17677 15544 17682 15600
rect 17738 15544 20350 15600
rect 20406 15544 20718 15600
rect 20774 15544 20779 15600
rect 17677 15542 20779 15544
rect 17677 15539 17743 15542
rect 20345 15539 20411 15542
rect 20713 15539 20779 15542
rect 16481 15466 16547 15469
rect 27520 15466 28000 15496
rect 16481 15464 28000 15466
rect 16481 15408 16486 15464
rect 16542 15408 28000 15464
rect 16481 15406 28000 15408
rect 16481 15403 16547 15406
rect 27520 15376 28000 15406
rect 21725 15330 21791 15333
rect 23749 15330 23815 15333
rect 21725 15328 23815 15330
rect 21725 15272 21730 15328
rect 21786 15272 23754 15328
rect 23810 15272 23815 15328
rect 21725 15270 23815 15272
rect 21725 15267 21791 15270
rect 23749 15267 23815 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 13813 15058 13879 15061
rect 21817 15058 21883 15061
rect 13813 15056 21883 15058
rect 13813 15000 13818 15056
rect 13874 15000 21822 15056
rect 21878 15000 21883 15056
rect 13813 14998 21883 15000
rect 13813 14995 13879 14998
rect 21817 14995 21883 14998
rect 18413 14922 18479 14925
rect 22001 14922 22067 14925
rect 18413 14920 22067 14922
rect 18413 14864 18418 14920
rect 18474 14864 22006 14920
rect 22062 14864 22067 14920
rect 18413 14862 22067 14864
rect 18413 14859 18479 14862
rect 22001 14859 22067 14862
rect 23933 14922 23999 14925
rect 27520 14922 28000 14952
rect 23933 14920 28000 14922
rect 23933 14864 23938 14920
rect 23994 14864 28000 14920
rect 23933 14862 28000 14864
rect 23933 14859 23999 14862
rect 27520 14832 28000 14862
rect 16481 14786 16547 14789
rect 17033 14786 17099 14789
rect 18505 14786 18571 14789
rect 16481 14784 18571 14786
rect 16481 14728 16486 14784
rect 16542 14728 17038 14784
rect 17094 14728 18510 14784
rect 18566 14728 18571 14784
rect 16481 14726 18571 14728
rect 16481 14723 16547 14726
rect 17033 14723 17099 14726
rect 18505 14723 18571 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 13997 14514 14063 14517
rect 21357 14514 21423 14517
rect 13997 14512 21423 14514
rect 13997 14456 14002 14512
rect 14058 14456 21362 14512
rect 21418 14456 21423 14512
rect 13997 14454 21423 14456
rect 13997 14451 14063 14454
rect 21357 14451 21423 14454
rect 13261 14378 13327 14381
rect 21265 14378 21331 14381
rect 13261 14376 21331 14378
rect 13261 14320 13266 14376
rect 13322 14320 21270 14376
rect 21326 14320 21331 14376
rect 13261 14318 21331 14320
rect 13261 14315 13327 14318
rect 21265 14315 21331 14318
rect 24209 14378 24275 14381
rect 27520 14378 28000 14408
rect 24209 14376 28000 14378
rect 24209 14320 24214 14376
rect 24270 14320 28000 14376
rect 24209 14318 28000 14320
rect 24209 14315 24275 14318
rect 27520 14288 28000 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13970 480 14000
rect 1577 13970 1643 13973
rect 0 13968 1643 13970
rect 0 13912 1582 13968
rect 1638 13912 1643 13968
rect 0 13910 1643 13912
rect 0 13880 480 13910
rect 1577 13907 1643 13910
rect 9949 13970 10015 13973
rect 13353 13970 13419 13973
rect 9949 13968 13419 13970
rect 9949 13912 9954 13968
rect 10010 13912 13358 13968
rect 13414 13912 13419 13968
rect 9949 13910 13419 13912
rect 9949 13907 10015 13910
rect 13353 13907 13419 13910
rect 13813 13970 13879 13973
rect 17401 13970 17467 13973
rect 13813 13968 17467 13970
rect 13813 13912 13818 13968
rect 13874 13912 17406 13968
rect 17462 13912 17467 13968
rect 13813 13910 17467 13912
rect 13813 13907 13879 13910
rect 17401 13907 17467 13910
rect 18689 13970 18755 13973
rect 24710 13970 24716 13972
rect 18689 13968 24716 13970
rect 18689 13912 18694 13968
rect 18750 13912 24716 13968
rect 18689 13910 24716 13912
rect 18689 13907 18755 13910
rect 24710 13908 24716 13910
rect 24780 13908 24786 13972
rect 14774 13772 14780 13836
rect 14844 13834 14850 13836
rect 17769 13834 17835 13837
rect 14844 13832 17835 13834
rect 14844 13776 17774 13832
rect 17830 13776 17835 13832
rect 14844 13774 17835 13776
rect 14844 13772 14850 13774
rect 17769 13771 17835 13774
rect 21357 13834 21423 13837
rect 22921 13834 22987 13837
rect 21357 13832 22987 13834
rect 21357 13776 21362 13832
rect 21418 13776 22926 13832
rect 22982 13776 22987 13832
rect 21357 13774 22987 13776
rect 21357 13771 21423 13774
rect 22921 13771 22987 13774
rect 23197 13698 23263 13701
rect 27520 13698 28000 13728
rect 23197 13696 28000 13698
rect 23197 13640 23202 13696
rect 23258 13640 28000 13696
rect 23197 13638 28000 13640
rect 23197 13635 23263 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 27520 13608 28000 13638
rect 19610 13567 19930 13568
rect 11053 13426 11119 13429
rect 25129 13426 25195 13429
rect 11053 13424 25195 13426
rect 11053 13368 11058 13424
rect 11114 13368 25134 13424
rect 25190 13368 25195 13424
rect 11053 13366 25195 13368
rect 11053 13363 11119 13366
rect 25129 13363 25195 13366
rect 13169 13290 13235 13293
rect 20897 13290 20963 13293
rect 13169 13288 20963 13290
rect 13169 13232 13174 13288
rect 13230 13232 20902 13288
rect 20958 13232 20963 13288
rect 13169 13230 20963 13232
rect 13169 13227 13235 13230
rect 20897 13227 20963 13230
rect 25681 13154 25747 13157
rect 27520 13154 28000 13184
rect 25681 13152 28000 13154
rect 25681 13096 25686 13152
rect 25742 13096 28000 13152
rect 25681 13094 28000 13096
rect 25681 13091 25747 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13094
rect 24277 13023 24597 13024
rect 381 12882 447 12885
rect 9121 12882 9187 12885
rect 12709 12882 12775 12885
rect 16021 12882 16087 12885
rect 16389 12882 16455 12885
rect 381 12880 16087 12882
rect 381 12824 386 12880
rect 442 12824 9126 12880
rect 9182 12824 12714 12880
rect 12770 12824 16026 12880
rect 16082 12824 16087 12880
rect 381 12822 16087 12824
rect 381 12819 447 12822
rect 9121 12819 9187 12822
rect 12709 12819 12775 12822
rect 16021 12819 16087 12822
rect 16254 12880 16455 12882
rect 16254 12824 16394 12880
rect 16450 12824 16455 12880
rect 16254 12822 16455 12824
rect 9489 12746 9555 12749
rect 15285 12746 15351 12749
rect 16254 12746 16314 12822
rect 16389 12819 16455 12822
rect 9489 12744 15351 12746
rect 9489 12688 9494 12744
rect 9550 12688 15290 12744
rect 15346 12688 15351 12744
rect 9489 12686 15351 12688
rect 9489 12683 9555 12686
rect 15285 12683 15351 12686
rect 15748 12686 16314 12746
rect 16389 12746 16455 12749
rect 19517 12746 19583 12749
rect 16389 12744 19583 12746
rect 16389 12688 16394 12744
rect 16450 12688 19522 12744
rect 19578 12688 19583 12744
rect 16389 12686 19583 12688
rect 12893 12610 12959 12613
rect 13169 12610 13235 12613
rect 12893 12608 13235 12610
rect 12893 12552 12898 12608
rect 12954 12552 13174 12608
rect 13230 12552 13235 12608
rect 12893 12550 13235 12552
rect 12893 12547 12959 12550
rect 13169 12547 13235 12550
rect 13353 12610 13419 12613
rect 15748 12610 15808 12686
rect 16389 12683 16455 12686
rect 19517 12683 19583 12686
rect 13353 12608 15808 12610
rect 13353 12552 13358 12608
rect 13414 12552 15808 12608
rect 13353 12550 15808 12552
rect 15929 12610 15995 12613
rect 16246 12610 16252 12612
rect 15929 12608 16252 12610
rect 15929 12552 15934 12608
rect 15990 12552 16252 12608
rect 15929 12550 16252 12552
rect 13353 12547 13419 12550
rect 15929 12547 15995 12550
rect 16246 12548 16252 12550
rect 16316 12548 16322 12612
rect 24117 12610 24183 12613
rect 27520 12610 28000 12640
rect 24117 12608 28000 12610
rect 24117 12552 24122 12608
rect 24178 12552 28000 12608
rect 24117 12550 28000 12552
rect 24117 12547 24183 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 27520 12520 28000 12550
rect 19610 12479 19930 12480
rect 1485 12474 1551 12477
rect 2313 12474 2379 12477
rect 1485 12472 2379 12474
rect 1485 12416 1490 12472
rect 1546 12416 2318 12472
rect 2374 12416 2379 12472
rect 1485 12414 2379 12416
rect 1485 12411 1551 12414
rect 2313 12411 2379 12414
rect 15377 12474 15443 12477
rect 15929 12474 15995 12477
rect 15377 12472 15995 12474
rect 15377 12416 15382 12472
rect 15438 12416 15934 12472
rect 15990 12416 15995 12472
rect 15377 12414 15995 12416
rect 15377 12411 15443 12414
rect 15929 12411 15995 12414
rect 20529 12474 20595 12477
rect 23749 12474 23815 12477
rect 20529 12472 23815 12474
rect 20529 12416 20534 12472
rect 20590 12416 23754 12472
rect 23810 12416 23815 12472
rect 20529 12414 23815 12416
rect 20529 12411 20595 12414
rect 23749 12411 23815 12414
rect 13169 12338 13235 12341
rect 15745 12338 15811 12341
rect 13169 12336 15811 12338
rect 13169 12280 13174 12336
rect 13230 12280 15750 12336
rect 15806 12280 15811 12336
rect 13169 12278 15811 12280
rect 13169 12275 13235 12278
rect 15745 12275 15811 12278
rect 16205 12340 16271 12341
rect 16205 12336 16252 12340
rect 16316 12338 16322 12340
rect 16573 12338 16639 12341
rect 18689 12338 18755 12341
rect 24209 12338 24275 12341
rect 16205 12280 16210 12336
rect 16205 12276 16252 12280
rect 16316 12278 16362 12338
rect 16573 12336 18755 12338
rect 16573 12280 16578 12336
rect 16634 12280 18694 12336
rect 18750 12280 18755 12336
rect 16573 12278 18755 12280
rect 16316 12276 16322 12278
rect 16205 12275 16271 12276
rect 16573 12275 16639 12278
rect 18689 12275 18755 12278
rect 18830 12336 24275 12338
rect 18830 12280 24214 12336
rect 24270 12280 24275 12336
rect 18830 12278 24275 12280
rect 13537 12202 13603 12205
rect 16757 12202 16823 12205
rect 13537 12200 16823 12202
rect 13537 12144 13542 12200
rect 13598 12144 16762 12200
rect 16818 12144 16823 12200
rect 13537 12142 16823 12144
rect 13537 12139 13603 12142
rect 16757 12139 16823 12142
rect 17309 12202 17375 12205
rect 18505 12202 18571 12205
rect 18830 12202 18890 12278
rect 24209 12275 24275 12278
rect 20805 12202 20871 12205
rect 24577 12202 24643 12205
rect 17309 12200 18890 12202
rect 17309 12144 17314 12200
rect 17370 12144 18510 12200
rect 18566 12144 18890 12200
rect 17309 12142 18890 12144
rect 18968 12200 24643 12202
rect 18968 12144 20810 12200
rect 20866 12144 24582 12200
rect 24638 12144 24643 12200
rect 18968 12142 24643 12144
rect 17309 12139 17375 12142
rect 18505 12139 18571 12142
rect 10961 12066 11027 12069
rect 12617 12066 12683 12069
rect 10961 12064 12683 12066
rect 10961 12008 10966 12064
rect 11022 12008 12622 12064
rect 12678 12008 12683 12064
rect 10961 12006 12683 12008
rect 10961 12003 11027 12006
rect 12617 12003 12683 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 11513 11930 11579 11933
rect 13905 11930 13971 11933
rect 11513 11928 13971 11930
rect 11513 11872 11518 11928
rect 11574 11872 13910 11928
rect 13966 11872 13971 11928
rect 11513 11870 13971 11872
rect 11513 11867 11579 11870
rect 13905 11867 13971 11870
rect 13997 11794 14063 11797
rect 18968 11794 19028 12142
rect 20805 12139 20871 12142
rect 24577 12139 24643 12142
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 27520 11930 28000 11960
rect 25822 11870 28000 11930
rect 13997 11792 19028 11794
rect 13997 11736 14002 11792
rect 14058 11736 19028 11792
rect 13997 11734 19028 11736
rect 24025 11794 24091 11797
rect 25589 11794 25655 11797
rect 24025 11792 25655 11794
rect 24025 11736 24030 11792
rect 24086 11736 25594 11792
rect 25650 11736 25655 11792
rect 24025 11734 25655 11736
rect 13997 11731 14063 11734
rect 24025 11731 24091 11734
rect 25589 11731 25655 11734
rect 9581 11658 9647 11661
rect 16297 11658 16363 11661
rect 17309 11658 17375 11661
rect 23933 11658 23999 11661
rect 9581 11656 10794 11658
rect 9581 11600 9586 11656
rect 9642 11600 10794 11656
rect 9581 11598 10794 11600
rect 9581 11595 9647 11598
rect 10734 11522 10794 11598
rect 16297 11656 17375 11658
rect 16297 11600 16302 11656
rect 16358 11600 17314 11656
rect 17370 11600 17375 11656
rect 16297 11598 17375 11600
rect 16297 11595 16363 11598
rect 17309 11595 17375 11598
rect 17542 11656 23999 11658
rect 17542 11600 23938 11656
rect 23994 11600 23999 11656
rect 17542 11598 23999 11600
rect 17401 11522 17467 11525
rect 10734 11520 17467 11522
rect 10734 11464 17406 11520
rect 17462 11464 17467 11520
rect 10734 11462 17467 11464
rect 17401 11459 17467 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 14181 11386 14247 11389
rect 14365 11386 14431 11389
rect 17542 11386 17602 11598
rect 23933 11595 23999 11598
rect 24301 11658 24367 11661
rect 25822 11658 25882 11870
rect 27520 11840 28000 11870
rect 24301 11656 25882 11658
rect 24301 11600 24306 11656
rect 24362 11600 25882 11656
rect 24301 11598 25882 11600
rect 24301 11595 24367 11598
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 27520 11386 28000 11416
rect 14181 11384 17602 11386
rect 14181 11328 14186 11384
rect 14242 11328 14370 11384
rect 14426 11328 17602 11384
rect 14181 11326 17602 11328
rect 23016 11326 28000 11386
rect 14181 11323 14247 11326
rect 14365 11323 14431 11326
rect 9213 11250 9279 11253
rect 12341 11250 12407 11253
rect 9213 11248 12407 11250
rect 9213 11192 9218 11248
rect 9274 11192 12346 11248
rect 12402 11192 12407 11248
rect 9213 11190 12407 11192
rect 9213 11187 9279 11190
rect 12341 11187 12407 11190
rect 17309 11250 17375 11253
rect 23016 11250 23076 11326
rect 27520 11296 28000 11326
rect 17309 11248 23076 11250
rect 17309 11192 17314 11248
rect 17370 11192 23076 11248
rect 17309 11190 23076 11192
rect 17309 11187 17375 11190
rect 2037 11114 2103 11117
rect 8937 11114 9003 11117
rect 9857 11114 9923 11117
rect 2037 11112 9923 11114
rect 2037 11056 2042 11112
rect 2098 11056 8942 11112
rect 8998 11056 9862 11112
rect 9918 11056 9923 11112
rect 2037 11054 9923 11056
rect 2037 11051 2103 11054
rect 8937 11051 9003 11054
rect 9857 11051 9923 11054
rect 14733 11114 14799 11117
rect 16941 11114 17007 11117
rect 24301 11114 24367 11117
rect 14733 11112 17007 11114
rect 14733 11056 14738 11112
rect 14794 11056 16946 11112
rect 17002 11056 17007 11112
rect 14733 11054 17007 11056
rect 14733 11051 14799 11054
rect 16941 11051 17007 11054
rect 24120 11112 24367 11114
rect 24120 11056 24306 11112
rect 24362 11056 24367 11112
rect 24120 11054 24367 11056
rect 11697 10978 11763 10981
rect 14774 10978 14780 10980
rect 11697 10976 14780 10978
rect 11697 10920 11702 10976
rect 11758 10920 14780 10976
rect 11697 10918 14780 10920
rect 11697 10915 11763 10918
rect 14774 10916 14780 10918
rect 14844 10916 14850 10980
rect 18321 10978 18387 10981
rect 18873 10978 18939 10981
rect 21449 10978 21515 10981
rect 18321 10976 21515 10978
rect 18321 10920 18326 10976
rect 18382 10920 18878 10976
rect 18934 10920 21454 10976
rect 21510 10920 21515 10976
rect 18321 10918 21515 10920
rect 18321 10915 18387 10918
rect 18873 10915 18939 10918
rect 21449 10915 21515 10918
rect 21725 10978 21791 10981
rect 23606 10978 23612 10980
rect 21725 10976 23612 10978
rect 21725 10920 21730 10976
rect 21786 10920 23612 10976
rect 21725 10918 23612 10920
rect 21725 10915 21791 10918
rect 23606 10916 23612 10918
rect 23676 10978 23682 10980
rect 24120 10978 24180 11054
rect 24301 11051 24367 11054
rect 23676 10918 24180 10978
rect 23676 10916 23682 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 17769 10842 17835 10845
rect 21357 10842 21423 10845
rect 23197 10842 23263 10845
rect 27520 10842 28000 10872
rect 17769 10840 21423 10842
rect 17769 10784 17774 10840
rect 17830 10784 21362 10840
rect 21418 10784 21423 10840
rect 17769 10782 21423 10784
rect 17769 10779 17835 10782
rect 21357 10779 21423 10782
rect 21590 10840 23263 10842
rect 21590 10784 23202 10840
rect 23258 10784 23263 10840
rect 21590 10782 23263 10784
rect 2773 10706 2839 10709
rect 9305 10706 9371 10709
rect 2773 10704 9371 10706
rect 2773 10648 2778 10704
rect 2834 10648 9310 10704
rect 9366 10648 9371 10704
rect 2773 10646 9371 10648
rect 2773 10643 2839 10646
rect 9305 10643 9371 10646
rect 9581 10706 9647 10709
rect 17401 10706 17467 10709
rect 19977 10706 20043 10709
rect 21590 10706 21650 10782
rect 23197 10779 23263 10782
rect 24902 10782 28000 10842
rect 9581 10704 19810 10706
rect 9581 10648 9586 10704
rect 9642 10648 17406 10704
rect 17462 10648 19810 10704
rect 9581 10646 19810 10648
rect 9581 10643 9647 10646
rect 17401 10643 17467 10646
rect 14825 10570 14891 10573
rect 19057 10570 19123 10573
rect 14825 10568 19123 10570
rect 14825 10512 14830 10568
rect 14886 10512 19062 10568
rect 19118 10512 19123 10568
rect 14825 10510 19123 10512
rect 19750 10570 19810 10646
rect 19977 10704 21650 10706
rect 19977 10648 19982 10704
rect 20038 10648 21650 10704
rect 19977 10646 21650 10648
rect 22001 10706 22067 10709
rect 24902 10706 24962 10782
rect 27520 10752 28000 10782
rect 22001 10704 24962 10706
rect 22001 10648 22006 10704
rect 22062 10648 24962 10704
rect 22001 10646 24962 10648
rect 19977 10643 20043 10646
rect 22001 10643 22067 10646
rect 19750 10510 21282 10570
rect 14825 10507 14891 10510
rect 19057 10507 19123 10510
rect 13997 10434 14063 10437
rect 15377 10434 15443 10437
rect 13997 10432 15443 10434
rect 13997 10376 14002 10432
rect 14058 10376 15382 10432
rect 15438 10376 15443 10432
rect 13997 10374 15443 10376
rect 13997 10371 14063 10374
rect 15377 10371 15443 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 16297 10298 16363 10301
rect 10734 10296 16363 10298
rect 10734 10240 16302 10296
rect 16358 10240 16363 10296
rect 10734 10238 16363 10240
rect 4981 10162 5047 10165
rect 10734 10162 10794 10238
rect 16297 10235 16363 10238
rect 4981 10160 10794 10162
rect 4981 10104 4986 10160
rect 5042 10104 10794 10160
rect 4981 10102 10794 10104
rect 13353 10162 13419 10165
rect 21081 10162 21147 10165
rect 13353 10160 21147 10162
rect 13353 10104 13358 10160
rect 13414 10104 21086 10160
rect 21142 10104 21147 10160
rect 13353 10102 21147 10104
rect 21222 10162 21282 10510
rect 21449 10298 21515 10301
rect 21449 10296 23812 10298
rect 21449 10240 21454 10296
rect 21510 10240 23812 10296
rect 21449 10238 23812 10240
rect 21449 10235 21515 10238
rect 23752 10162 23812 10238
rect 27520 10162 28000 10192
rect 21222 10102 23306 10162
rect 23752 10102 28000 10162
rect 4981 10099 5047 10102
rect 13353 10099 13419 10102
rect 21081 10099 21147 10102
rect 13629 10026 13695 10029
rect 13997 10026 14063 10029
rect 19333 10026 19399 10029
rect 13629 10024 19399 10026
rect 13629 9968 13634 10024
rect 13690 9968 14002 10024
rect 14058 9968 19338 10024
rect 19394 9968 19399 10024
rect 13629 9966 19399 9968
rect 13629 9963 13695 9966
rect 13997 9963 14063 9966
rect 19333 9963 19399 9966
rect 19701 10026 19767 10029
rect 22001 10026 22067 10029
rect 19701 10024 22067 10026
rect 19701 9968 19706 10024
rect 19762 9968 22006 10024
rect 22062 9968 22067 10024
rect 19701 9966 22067 9968
rect 19701 9963 19767 9966
rect 22001 9963 22067 9966
rect 15653 9890 15719 9893
rect 15837 9890 15903 9893
rect 15653 9888 15903 9890
rect 15653 9832 15658 9888
rect 15714 9832 15842 9888
rect 15898 9832 15903 9888
rect 15653 9830 15903 9832
rect 15653 9827 15719 9830
rect 15837 9827 15903 9830
rect 16481 9890 16547 9893
rect 21633 9890 21699 9893
rect 16481 9888 21699 9890
rect 16481 9832 16486 9888
rect 16542 9832 21638 9888
rect 21694 9832 21699 9888
rect 16481 9830 21699 9832
rect 23246 9890 23306 10102
rect 27520 10072 28000 10102
rect 23381 10026 23447 10029
rect 25129 10026 25195 10029
rect 23381 10024 25195 10026
rect 23381 9968 23386 10024
rect 23442 9968 25134 10024
rect 25190 9968 25195 10024
rect 23381 9966 25195 9968
rect 23381 9963 23447 9966
rect 25129 9963 25195 9966
rect 23841 9890 23907 9893
rect 23246 9888 23907 9890
rect 23246 9832 23846 9888
rect 23902 9832 23907 9888
rect 23246 9830 23907 9832
rect 16481 9827 16547 9830
rect 21633 9827 21699 9830
rect 23841 9827 23907 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 15377 9754 15443 9757
rect 16389 9754 16455 9757
rect 19701 9754 19767 9757
rect 15377 9752 19767 9754
rect 15377 9696 15382 9752
rect 15438 9696 16394 9752
rect 16450 9696 19706 9752
rect 19762 9696 19767 9752
rect 15377 9694 19767 9696
rect 15377 9691 15443 9694
rect 16389 9691 16455 9694
rect 19701 9691 19767 9694
rect 21081 9754 21147 9757
rect 21081 9752 24180 9754
rect 21081 9696 21086 9752
rect 21142 9696 24180 9752
rect 21081 9694 24180 9696
rect 21081 9691 21147 9694
rect 11237 9618 11303 9621
rect 13905 9618 13971 9621
rect 11237 9616 13971 9618
rect 11237 9560 11242 9616
rect 11298 9560 13910 9616
rect 13966 9560 13971 9616
rect 11237 9558 13971 9560
rect 11237 9555 11303 9558
rect 13905 9555 13971 9558
rect 14733 9618 14799 9621
rect 20253 9618 20319 9621
rect 22185 9618 22251 9621
rect 14733 9616 22251 9618
rect 14733 9560 14738 9616
rect 14794 9560 20258 9616
rect 20314 9560 22190 9616
rect 22246 9560 22251 9616
rect 14733 9558 22251 9560
rect 24120 9618 24180 9694
rect 27520 9618 28000 9648
rect 24120 9558 28000 9618
rect 14733 9555 14799 9558
rect 20253 9555 20319 9558
rect 22185 9555 22251 9558
rect 27520 9528 28000 9558
rect 13169 9482 13235 9485
rect 21357 9482 21423 9485
rect 13169 9480 21423 9482
rect 13169 9424 13174 9480
rect 13230 9424 21362 9480
rect 21418 9424 21423 9480
rect 13169 9422 21423 9424
rect 13169 9419 13235 9422
rect 21357 9419 21423 9422
rect 11973 9346 12039 9349
rect 15377 9346 15443 9349
rect 11973 9344 16498 9346
rect 11973 9288 11978 9344
rect 12034 9288 15382 9344
rect 15438 9288 16498 9344
rect 11973 9286 16498 9288
rect 11973 9283 12039 9286
rect 15377 9283 15443 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 15469 9210 15535 9213
rect 10734 9208 15535 9210
rect 10734 9152 15474 9208
rect 15530 9152 15535 9208
rect 10734 9150 15535 9152
rect 9765 9074 9831 9077
rect 10734 9074 10794 9150
rect 15469 9147 15535 9150
rect 9765 9072 10794 9074
rect 9765 9016 9770 9072
rect 9826 9016 10794 9072
rect 9765 9014 10794 9016
rect 11513 9074 11579 9077
rect 14365 9074 14431 9077
rect 11513 9072 14431 9074
rect 11513 9016 11518 9072
rect 11574 9016 14370 9072
rect 14426 9016 14431 9072
rect 11513 9014 14431 9016
rect 16438 9074 16498 9286
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 23013 9074 23079 9077
rect 16438 9072 23079 9074
rect 16438 9016 23018 9072
rect 23074 9016 23079 9072
rect 16438 9014 23079 9016
rect 9765 9011 9831 9014
rect 11513 9011 11579 9014
rect 14365 9011 14431 9014
rect 23013 9011 23079 9014
rect 25037 9074 25103 9077
rect 27520 9074 28000 9104
rect 25037 9072 28000 9074
rect 25037 9016 25042 9072
rect 25098 9016 28000 9072
rect 25037 9014 28000 9016
rect 25037 9011 25103 9014
rect 27520 8984 28000 9014
rect 2313 8938 2379 8941
rect 10777 8938 10843 8941
rect 2313 8936 10843 8938
rect 2313 8880 2318 8936
rect 2374 8880 10782 8936
rect 10838 8880 10843 8936
rect 2313 8878 10843 8880
rect 2313 8875 2379 8878
rect 10777 8875 10843 8878
rect 21357 8938 21423 8941
rect 23565 8938 23631 8941
rect 21357 8936 23631 8938
rect 21357 8880 21362 8936
rect 21418 8880 23570 8936
rect 23626 8880 23631 8936
rect 21357 8878 23631 8880
rect 21357 8875 21423 8878
rect 23565 8875 23631 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 7097 8530 7163 8533
rect 16481 8530 16547 8533
rect 7097 8528 16547 8530
rect 7097 8472 7102 8528
rect 7158 8472 16486 8528
rect 16542 8472 16547 8528
rect 7097 8470 16547 8472
rect 7097 8467 7163 8470
rect 16481 8467 16547 8470
rect 23657 8530 23723 8533
rect 27520 8530 28000 8560
rect 23657 8528 28000 8530
rect 23657 8472 23662 8528
rect 23718 8472 28000 8528
rect 23657 8470 28000 8472
rect 23657 8467 23723 8470
rect 27520 8440 28000 8470
rect 18873 8394 18939 8397
rect 20989 8394 21055 8397
rect 18873 8392 21055 8394
rect 18873 8336 18878 8392
rect 18934 8336 20994 8392
rect 21050 8336 21055 8392
rect 18873 8334 21055 8336
rect 18873 8331 18939 8334
rect 20989 8331 21055 8334
rect 20161 8258 20227 8261
rect 23197 8258 23263 8261
rect 20161 8256 23263 8258
rect 20161 8200 20166 8256
rect 20222 8200 23202 8256
rect 23258 8200 23263 8256
rect 20161 8198 23263 8200
rect 20161 8195 20227 8198
rect 23197 8195 23263 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 17217 8122 17283 8125
rect 23657 8124 23723 8125
rect 13310 8120 17283 8122
rect 13310 8064 17222 8120
rect 17278 8064 17283 8120
rect 13310 8062 17283 8064
rect 3785 7986 3851 7989
rect 13310 7986 13370 8062
rect 17217 8059 17283 8062
rect 23606 8060 23612 8124
rect 23676 8122 23723 8124
rect 23676 8120 23768 8122
rect 23718 8064 23768 8120
rect 23676 8062 23768 8064
rect 23676 8060 23723 8062
rect 23657 8059 23723 8060
rect 3785 7984 13370 7986
rect 3785 7928 3790 7984
rect 3846 7928 13370 7984
rect 3785 7926 13370 7928
rect 13445 7986 13511 7989
rect 20345 7986 20411 7989
rect 13445 7984 20411 7986
rect 13445 7928 13450 7984
rect 13506 7928 20350 7984
rect 20406 7928 20411 7984
rect 13445 7926 20411 7928
rect 3785 7923 3851 7926
rect 13445 7923 13511 7926
rect 20345 7923 20411 7926
rect 7741 7850 7807 7853
rect 12801 7850 12867 7853
rect 7741 7848 12867 7850
rect 7741 7792 7746 7848
rect 7802 7792 12806 7848
rect 12862 7792 12867 7848
rect 7741 7790 12867 7792
rect 7741 7787 7807 7790
rect 12801 7787 12867 7790
rect 13629 7850 13695 7853
rect 19333 7850 19399 7853
rect 13629 7848 19399 7850
rect 13629 7792 13634 7848
rect 13690 7792 19338 7848
rect 19394 7792 19399 7848
rect 13629 7790 19399 7792
rect 13629 7787 13695 7790
rect 19333 7787 19399 7790
rect 21909 7850 21975 7853
rect 23105 7850 23171 7853
rect 27520 7850 28000 7880
rect 21909 7848 28000 7850
rect 21909 7792 21914 7848
rect 21970 7792 23110 7848
rect 23166 7792 28000 7848
rect 21909 7790 28000 7792
rect 21909 7787 21975 7790
rect 23105 7787 23171 7790
rect 27520 7760 28000 7790
rect 13077 7714 13143 7717
rect 6134 7712 13143 7714
rect 6134 7656 13082 7712
rect 13138 7656 13143 7712
rect 6134 7654 13143 7656
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 4337 7442 4403 7445
rect 6134 7442 6194 7654
rect 13077 7651 13143 7654
rect 15929 7714 15995 7717
rect 21725 7714 21791 7717
rect 15929 7712 21791 7714
rect 15929 7656 15934 7712
rect 15990 7656 21730 7712
rect 21786 7656 21791 7712
rect 15929 7654 21791 7656
rect 15929 7651 15995 7654
rect 21725 7651 21791 7654
rect 24669 7714 24735 7717
rect 25405 7714 25471 7717
rect 24669 7712 25471 7714
rect 24669 7656 24674 7712
rect 24730 7656 25410 7712
rect 25466 7656 25471 7712
rect 24669 7654 25471 7656
rect 24669 7651 24735 7654
rect 25405 7651 25471 7654
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 16297 7578 16363 7581
rect 22645 7578 22711 7581
rect 16297 7576 22711 7578
rect 16297 7520 16302 7576
rect 16358 7520 22650 7576
rect 22706 7520 22711 7576
rect 16297 7518 22711 7520
rect 16297 7515 16363 7518
rect 22645 7515 22711 7518
rect 4337 7440 6194 7442
rect 4337 7384 4342 7440
rect 4398 7384 6194 7440
rect 4337 7382 6194 7384
rect 11145 7442 11211 7445
rect 16481 7442 16547 7445
rect 21725 7442 21791 7445
rect 24761 7442 24827 7445
rect 11145 7440 16547 7442
rect 11145 7384 11150 7440
rect 11206 7384 16486 7440
rect 16542 7384 16547 7440
rect 11145 7382 16547 7384
rect 4337 7379 4403 7382
rect 11145 7379 11211 7382
rect 16481 7379 16547 7382
rect 16622 7382 21650 7442
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 16622 7034 16682 7382
rect 17217 7306 17283 7309
rect 21357 7306 21423 7309
rect 17217 7304 21423 7306
rect 17217 7248 17222 7304
rect 17278 7248 21362 7304
rect 21418 7248 21423 7304
rect 17217 7246 21423 7248
rect 21590 7306 21650 7382
rect 21725 7440 24827 7442
rect 21725 7384 21730 7440
rect 21786 7384 24766 7440
rect 24822 7384 24827 7440
rect 21725 7382 24827 7384
rect 21725 7379 21791 7382
rect 24761 7379 24827 7382
rect 25221 7306 25287 7309
rect 27520 7306 28000 7336
rect 21590 7304 25287 7306
rect 21590 7248 25226 7304
rect 25282 7248 25287 7304
rect 21590 7246 25287 7248
rect 17217 7243 17283 7246
rect 21357 7243 21423 7246
rect 25221 7243 25287 7246
rect 25454 7246 28000 7306
rect 23841 7170 23907 7173
rect 25454 7170 25514 7246
rect 27520 7216 28000 7246
rect 23841 7168 25514 7170
rect 23841 7112 23846 7168
rect 23902 7112 25514 7168
rect 23841 7110 25514 7112
rect 23841 7107 23907 7110
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 15150 6974 16682 7034
rect 3693 6898 3759 6901
rect 11973 6898 12039 6901
rect 3693 6896 12039 6898
rect 3693 6840 3698 6896
rect 3754 6840 11978 6896
rect 12034 6840 12039 6896
rect 3693 6838 12039 6840
rect 3693 6835 3759 6838
rect 11973 6835 12039 6838
rect 14457 6898 14523 6901
rect 15150 6898 15210 6974
rect 14457 6896 15210 6898
rect 14457 6840 14462 6896
rect 14518 6840 15210 6896
rect 14457 6838 15210 6840
rect 18137 6898 18203 6901
rect 22001 6898 22067 6901
rect 18137 6896 22067 6898
rect 18137 6840 18142 6896
rect 18198 6840 22006 6896
rect 22062 6840 22067 6896
rect 18137 6838 22067 6840
rect 14457 6835 14523 6838
rect 18137 6835 18203 6838
rect 22001 6835 22067 6838
rect 24117 6898 24183 6901
rect 25037 6898 25103 6901
rect 24117 6896 25103 6898
rect 24117 6840 24122 6896
rect 24178 6840 25042 6896
rect 25098 6840 25103 6896
rect 24117 6838 25103 6840
rect 24117 6835 24183 6838
rect 25037 6835 25103 6838
rect 6361 6762 6427 6765
rect 11237 6762 11303 6765
rect 6361 6760 11303 6762
rect 6361 6704 6366 6760
rect 6422 6704 11242 6760
rect 11298 6704 11303 6760
rect 6361 6702 11303 6704
rect 6361 6699 6427 6702
rect 11237 6699 11303 6702
rect 12065 6762 12131 6765
rect 14273 6762 14339 6765
rect 14917 6762 14983 6765
rect 12065 6760 14983 6762
rect 12065 6704 12070 6760
rect 12126 6704 14278 6760
rect 14334 6704 14922 6760
rect 14978 6704 14983 6760
rect 12065 6702 14983 6704
rect 12065 6699 12131 6702
rect 14273 6699 14339 6702
rect 14917 6699 14983 6702
rect 21449 6762 21515 6765
rect 24209 6762 24275 6765
rect 21449 6760 24275 6762
rect 21449 6704 21454 6760
rect 21510 6704 24214 6760
rect 24270 6704 24275 6760
rect 21449 6702 24275 6704
rect 21449 6699 21515 6702
rect 24209 6699 24275 6702
rect 24761 6762 24827 6765
rect 27520 6762 28000 6792
rect 24761 6760 28000 6762
rect 24761 6704 24766 6760
rect 24822 6704 28000 6760
rect 24761 6702 28000 6704
rect 24761 6699 24827 6702
rect 27520 6672 28000 6702
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 21081 6490 21147 6493
rect 19014 6488 21147 6490
rect 19014 6432 21086 6488
rect 21142 6432 21147 6488
rect 19014 6430 21147 6432
rect 9581 6354 9647 6357
rect 9857 6354 9923 6357
rect 19014 6354 19074 6430
rect 21081 6427 21147 6430
rect 21265 6490 21331 6493
rect 23657 6490 23723 6493
rect 21265 6488 23723 6490
rect 21265 6432 21270 6488
rect 21326 6432 23662 6488
rect 23718 6432 23723 6488
rect 21265 6430 23723 6432
rect 21265 6427 21331 6430
rect 23657 6427 23723 6430
rect 9581 6352 19074 6354
rect 9581 6296 9586 6352
rect 9642 6296 9862 6352
rect 9918 6296 19074 6352
rect 9581 6294 19074 6296
rect 19149 6354 19215 6357
rect 19149 6352 22018 6354
rect 19149 6296 19154 6352
rect 19210 6296 22018 6352
rect 19149 6294 22018 6296
rect 9581 6291 9647 6294
rect 9857 6291 9923 6294
rect 19149 6291 19215 6294
rect 14825 6218 14891 6221
rect 19609 6218 19675 6221
rect 14825 6216 19675 6218
rect 14825 6160 14830 6216
rect 14886 6160 19614 6216
rect 19670 6160 19675 6216
rect 14825 6158 19675 6160
rect 21958 6218 22018 6294
rect 21958 6158 22202 6218
rect 14825 6155 14891 6158
rect 19609 6155 19675 6158
rect 22142 6082 22202 6158
rect 27520 6082 28000 6112
rect 22142 6022 28000 6082
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 16849 5810 16915 5813
rect 25497 5810 25563 5813
rect 16849 5808 25563 5810
rect 16849 5752 16854 5808
rect 16910 5752 25502 5808
rect 25558 5752 25563 5808
rect 16849 5750 25563 5752
rect 16849 5747 16915 5750
rect 25497 5747 25563 5750
rect 11329 5674 11395 5677
rect 15837 5674 15903 5677
rect 11329 5672 15903 5674
rect 11329 5616 11334 5672
rect 11390 5616 15842 5672
rect 15898 5616 15903 5672
rect 11329 5614 15903 5616
rect 11329 5611 11395 5614
rect 15837 5611 15903 5614
rect 16205 5674 16271 5677
rect 19977 5674 20043 5677
rect 16205 5672 20043 5674
rect 16205 5616 16210 5672
rect 16266 5616 19982 5672
rect 20038 5616 20043 5672
rect 16205 5614 20043 5616
rect 16205 5611 16271 5614
rect 19977 5611 20043 5614
rect 23749 5674 23815 5677
rect 23749 5672 24778 5674
rect 23749 5616 23754 5672
rect 23810 5616 24778 5672
rect 23749 5614 24778 5616
rect 23749 5611 23815 5614
rect 24718 5538 24778 5614
rect 27520 5538 28000 5568
rect 24718 5478 28000 5538
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 27520 5448 28000 5478
rect 24277 5407 24597 5408
rect 11881 5402 11947 5405
rect 14549 5402 14615 5405
rect 11881 5400 14615 5402
rect 11881 5344 11886 5400
rect 11942 5344 14554 5400
rect 14610 5344 14615 5400
rect 11881 5342 14615 5344
rect 11881 5339 11947 5342
rect 14549 5339 14615 5342
rect 2957 5266 3023 5269
rect 17677 5266 17743 5269
rect 2957 5264 17743 5266
rect 2957 5208 2962 5264
rect 3018 5208 17682 5264
rect 17738 5208 17743 5264
rect 2957 5206 17743 5208
rect 2957 5203 3023 5206
rect 17677 5203 17743 5206
rect 18413 5266 18479 5269
rect 22737 5266 22803 5269
rect 18413 5264 22803 5266
rect 18413 5208 18418 5264
rect 18474 5208 22742 5264
rect 22798 5208 22803 5264
rect 18413 5206 22803 5208
rect 18413 5203 18479 5206
rect 22737 5203 22803 5206
rect 23197 5266 23263 5269
rect 25221 5266 25287 5269
rect 23197 5264 25287 5266
rect 23197 5208 23202 5264
rect 23258 5208 25226 5264
rect 25282 5208 25287 5264
rect 23197 5206 25287 5208
rect 23197 5203 23263 5206
rect 25221 5203 25287 5206
rect 13813 5130 13879 5133
rect 17493 5130 17559 5133
rect 13813 5128 17559 5130
rect 13813 5072 13818 5128
rect 13874 5072 17498 5128
rect 17554 5072 17559 5128
rect 13813 5070 17559 5072
rect 13813 5067 13879 5070
rect 17493 5067 17559 5070
rect 19241 5130 19307 5133
rect 20897 5130 20963 5133
rect 19241 5128 20963 5130
rect 19241 5072 19246 5128
rect 19302 5072 20902 5128
rect 20958 5072 20963 5128
rect 19241 5070 20963 5072
rect 19241 5067 19307 5070
rect 20897 5067 20963 5070
rect 11329 4994 11395 4997
rect 19333 4994 19399 4997
rect 11329 4992 19399 4994
rect 11329 4936 11334 4992
rect 11390 4936 19338 4992
rect 19394 4936 19399 4992
rect 11329 4934 19399 4936
rect 11329 4931 11395 4934
rect 19333 4931 19399 4934
rect 25681 4994 25747 4997
rect 27520 4994 28000 5024
rect 25681 4992 28000 4994
rect 25681 4936 25686 4992
rect 25742 4936 28000 4992
rect 25681 4934 28000 4936
rect 25681 4931 25747 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 27520 4904 28000 4934
rect 19610 4863 19930 4864
rect 14549 4858 14615 4861
rect 18045 4858 18111 4861
rect 14549 4856 18111 4858
rect 14549 4800 14554 4856
rect 14610 4800 18050 4856
rect 18106 4800 18111 4856
rect 14549 4798 18111 4800
rect 14549 4795 14615 4798
rect 18045 4795 18111 4798
rect 0 4722 480 4752
rect 3693 4722 3759 4725
rect 0 4720 3759 4722
rect 0 4664 3698 4720
rect 3754 4664 3759 4720
rect 0 4662 3759 4664
rect 0 4632 480 4662
rect 3693 4659 3759 4662
rect 17033 4722 17099 4725
rect 22829 4722 22895 4725
rect 17033 4720 22895 4722
rect 17033 4664 17038 4720
rect 17094 4664 22834 4720
rect 22890 4664 22895 4720
rect 17033 4662 22895 4664
rect 17033 4659 17099 4662
rect 22829 4659 22895 4662
rect 13629 4586 13695 4589
rect 614 4584 13695 4586
rect 614 4528 13634 4584
rect 13690 4528 13695 4584
rect 614 4526 13695 4528
rect 289 4450 355 4453
rect 614 4450 674 4526
rect 13629 4523 13695 4526
rect 15285 4586 15351 4589
rect 15929 4586 15995 4589
rect 22093 4586 22159 4589
rect 15285 4584 15808 4586
rect 15285 4528 15290 4584
rect 15346 4528 15808 4584
rect 15285 4526 15808 4528
rect 15285 4523 15351 4526
rect 289 4448 674 4450
rect 289 4392 294 4448
rect 350 4392 674 4448
rect 289 4390 674 4392
rect 15748 4450 15808 4526
rect 15929 4584 22159 4586
rect 15929 4528 15934 4584
rect 15990 4528 22098 4584
rect 22154 4528 22159 4584
rect 15929 4526 22159 4528
rect 15929 4523 15995 4526
rect 22093 4523 22159 4526
rect 20805 4450 20871 4453
rect 15748 4448 20871 4450
rect 15748 4392 20810 4448
rect 20866 4392 20871 4448
rect 15748 4390 20871 4392
rect 289 4387 355 4390
rect 20805 4387 20871 4390
rect 20989 4450 21055 4453
rect 23565 4450 23631 4453
rect 20989 4448 23631 4450
rect 20989 4392 20994 4448
rect 21050 4392 23570 4448
rect 23626 4392 23631 4448
rect 20989 4390 23631 4392
rect 20989 4387 21055 4390
rect 23565 4387 23631 4390
rect 25589 4450 25655 4453
rect 27520 4450 28000 4480
rect 25589 4448 28000 4450
rect 25589 4392 25594 4448
rect 25650 4392 28000 4448
rect 25589 4390 28000 4392
rect 25589 4387 25655 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4390
rect 24277 4319 24597 4320
rect 15561 4314 15627 4317
rect 21265 4314 21331 4317
rect 15561 4312 21331 4314
rect 15561 4256 15566 4312
rect 15622 4256 21270 4312
rect 21326 4256 21331 4312
rect 15561 4254 21331 4256
rect 15561 4251 15627 4254
rect 21265 4251 21331 4254
rect 933 4178 999 4181
rect 21633 4178 21699 4181
rect 933 4176 21699 4178
rect 933 4120 938 4176
rect 994 4120 21638 4176
rect 21694 4120 21699 4176
rect 933 4118 21699 4120
rect 933 4115 999 4118
rect 21633 4115 21699 4118
rect 22645 4178 22711 4181
rect 26141 4178 26207 4181
rect 22645 4176 26207 4178
rect 22645 4120 22650 4176
rect 22706 4120 26146 4176
rect 26202 4120 26207 4176
rect 22645 4118 26207 4120
rect 22645 4115 22711 4118
rect 26141 4115 26207 4118
rect 15469 4042 15535 4045
rect 17309 4042 17375 4045
rect 15469 4040 17375 4042
rect 15469 3984 15474 4040
rect 15530 3984 17314 4040
rect 17370 3984 17375 4040
rect 15469 3982 17375 3984
rect 15469 3979 15535 3982
rect 17309 3979 17375 3982
rect 11421 3906 11487 3909
rect 15929 3906 15995 3909
rect 11421 3904 15995 3906
rect 11421 3848 11426 3904
rect 11482 3848 15934 3904
rect 15990 3848 15995 3904
rect 11421 3846 15995 3848
rect 11421 3843 11487 3846
rect 15929 3843 15995 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 11421 3770 11487 3773
rect 12709 3770 12775 3773
rect 11421 3768 12775 3770
rect 11421 3712 11426 3768
rect 11482 3712 12714 3768
rect 12770 3712 12775 3768
rect 11421 3710 12775 3712
rect 11421 3707 11487 3710
rect 12709 3707 12775 3710
rect 12893 3770 12959 3773
rect 13261 3770 13327 3773
rect 12893 3768 13327 3770
rect 12893 3712 12898 3768
rect 12954 3712 13266 3768
rect 13322 3712 13327 3768
rect 12893 3710 13327 3712
rect 12893 3707 12959 3710
rect 13261 3707 13327 3710
rect 13537 3770 13603 3773
rect 19149 3770 19215 3773
rect 13537 3768 19215 3770
rect 13537 3712 13542 3768
rect 13598 3712 19154 3768
rect 19210 3712 19215 3768
rect 13537 3710 19215 3712
rect 13537 3707 13603 3710
rect 19149 3707 19215 3710
rect 23473 3770 23539 3773
rect 27520 3770 28000 3800
rect 23473 3768 28000 3770
rect 23473 3712 23478 3768
rect 23534 3712 28000 3768
rect 23473 3710 28000 3712
rect 23473 3707 23539 3710
rect 27520 3680 28000 3710
rect 11145 3634 11211 3637
rect 17953 3634 18019 3637
rect 11145 3632 18019 3634
rect 11145 3576 11150 3632
rect 11206 3576 17958 3632
rect 18014 3576 18019 3632
rect 11145 3574 18019 3576
rect 11145 3571 11211 3574
rect 17953 3571 18019 3574
rect 18689 3634 18755 3637
rect 21173 3634 21239 3637
rect 24669 3634 24735 3637
rect 18689 3632 24735 3634
rect 18689 3576 18694 3632
rect 18750 3576 21178 3632
rect 21234 3576 24674 3632
rect 24730 3576 24735 3632
rect 18689 3574 24735 3576
rect 18689 3571 18755 3574
rect 21173 3571 21239 3574
rect 24669 3571 24735 3574
rect 10041 3498 10107 3501
rect 15469 3498 15535 3501
rect 10041 3496 15535 3498
rect 10041 3440 10046 3496
rect 10102 3440 15474 3496
rect 15530 3440 15535 3496
rect 10041 3438 15535 3440
rect 10041 3435 10107 3438
rect 15469 3435 15535 3438
rect 17769 3498 17835 3501
rect 18413 3498 18479 3501
rect 19517 3498 19583 3501
rect 19885 3498 19951 3501
rect 17769 3496 19951 3498
rect 17769 3440 17774 3496
rect 17830 3440 18418 3496
rect 18474 3440 19522 3496
rect 19578 3440 19890 3496
rect 19946 3440 19951 3496
rect 17769 3438 19951 3440
rect 17769 3435 17835 3438
rect 18413 3435 18479 3438
rect 19517 3435 19583 3438
rect 19885 3435 19951 3438
rect 25405 3498 25471 3501
rect 27521 3498 27587 3501
rect 25405 3496 27587 3498
rect 25405 3440 25410 3496
rect 25466 3440 27526 3496
rect 27582 3440 27587 3496
rect 25405 3438 27587 3440
rect 25405 3435 25471 3438
rect 27521 3435 27587 3438
rect 8385 3362 8451 3365
rect 11789 3362 11855 3365
rect 8385 3360 11855 3362
rect 8385 3304 8390 3360
rect 8446 3304 11794 3360
rect 11850 3304 11855 3360
rect 8385 3302 11855 3304
rect 8385 3299 8451 3302
rect 11789 3299 11855 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 24710 3164 24716 3228
rect 24780 3226 24786 3228
rect 27520 3226 28000 3256
rect 24780 3166 28000 3226
rect 24780 3164 24786 3166
rect 27520 3136 28000 3166
rect 10317 3090 10383 3093
rect 16573 3090 16639 3093
rect 10317 3088 16639 3090
rect 10317 3032 10322 3088
rect 10378 3032 16578 3088
rect 16634 3032 16639 3088
rect 10317 3030 16639 3032
rect 10317 3027 10383 3030
rect 16573 3027 16639 3030
rect 22369 3090 22435 3093
rect 24117 3090 24183 3093
rect 22369 3088 24183 3090
rect 22369 3032 22374 3088
rect 22430 3032 24122 3088
rect 24178 3032 24183 3088
rect 22369 3030 24183 3032
rect 22369 3027 22435 3030
rect 24117 3027 24183 3030
rect 13169 2954 13235 2957
rect 23841 2954 23907 2957
rect 13169 2952 23907 2954
rect 13169 2896 13174 2952
rect 13230 2896 23846 2952
rect 23902 2896 23907 2952
rect 13169 2894 23907 2896
rect 13169 2891 13235 2894
rect 23841 2891 23907 2894
rect 24577 2954 24643 2957
rect 24710 2954 24716 2956
rect 24577 2952 24716 2954
rect 24577 2896 24582 2952
rect 24638 2896 24716 2952
rect 24577 2894 24716 2896
rect 24577 2891 24643 2894
rect 24710 2892 24716 2894
rect 24780 2892 24786 2956
rect 11973 2818 12039 2821
rect 12709 2818 12775 2821
rect 19425 2818 19491 2821
rect 11973 2816 12450 2818
rect 11973 2760 11978 2816
rect 12034 2760 12450 2816
rect 11973 2758 12450 2760
rect 11973 2755 12039 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 12390 2682 12450 2758
rect 12709 2816 19491 2818
rect 12709 2760 12714 2816
rect 12770 2760 19430 2816
rect 19486 2760 19491 2816
rect 12709 2758 19491 2760
rect 12709 2755 12775 2758
rect 19425 2755 19491 2758
rect 20069 2818 20135 2821
rect 24761 2818 24827 2821
rect 20069 2816 24827 2818
rect 20069 2760 20074 2816
rect 20130 2760 24766 2816
rect 24822 2760 24827 2816
rect 20069 2758 24827 2760
rect 20069 2755 20135 2758
rect 24761 2755 24827 2758
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 12893 2682 12959 2685
rect 18965 2682 19031 2685
rect 12390 2680 19031 2682
rect 12390 2624 12898 2680
rect 12954 2624 18970 2680
rect 19026 2624 19031 2680
rect 12390 2622 19031 2624
rect 12893 2619 12959 2622
rect 18965 2619 19031 2622
rect 21909 2682 21975 2685
rect 24485 2682 24551 2685
rect 21909 2680 24551 2682
rect 21909 2624 21914 2680
rect 21970 2624 24490 2680
rect 24546 2624 24551 2680
rect 21909 2622 24551 2624
rect 21909 2619 21975 2622
rect 24485 2619 24551 2622
rect 24669 2682 24735 2685
rect 27520 2682 28000 2712
rect 24669 2680 28000 2682
rect 24669 2624 24674 2680
rect 24730 2624 28000 2680
rect 24669 2622 28000 2624
rect 24669 2619 24735 2622
rect 27520 2592 28000 2622
rect 1577 2546 1643 2549
rect 9949 2546 10015 2549
rect 14273 2546 14339 2549
rect 1577 2544 6194 2546
rect 1577 2488 1582 2544
rect 1638 2488 6194 2544
rect 1577 2486 6194 2488
rect 1577 2483 1643 2486
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 6134 2138 6194 2486
rect 9949 2544 14339 2546
rect 9949 2488 9954 2544
rect 10010 2488 14278 2544
rect 14334 2488 14339 2544
rect 9949 2486 14339 2488
rect 9949 2483 10015 2486
rect 14273 2483 14339 2486
rect 17769 2546 17835 2549
rect 25221 2546 25287 2549
rect 17769 2544 25287 2546
rect 17769 2488 17774 2544
rect 17830 2488 25226 2544
rect 25282 2488 25287 2544
rect 17769 2486 25287 2488
rect 17769 2483 17835 2486
rect 25221 2483 25287 2486
rect 9213 2410 9279 2413
rect 18597 2410 18663 2413
rect 9213 2408 18663 2410
rect 9213 2352 9218 2408
rect 9274 2352 18602 2408
rect 18658 2352 18663 2408
rect 9213 2350 18663 2352
rect 9213 2347 9279 2350
rect 18597 2347 18663 2350
rect 18830 2350 27538 2410
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 16389 2138 16455 2141
rect 18830 2138 18890 2350
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 6134 2078 11714 2138
rect 11654 2002 11714 2078
rect 16389 2136 18890 2138
rect 16389 2080 16394 2136
rect 16450 2080 18890 2136
rect 16389 2078 18890 2080
rect 18965 2138 19031 2141
rect 18965 2136 20914 2138
rect 18965 2080 18970 2136
rect 19026 2080 20914 2136
rect 18965 2078 20914 2080
rect 16389 2075 16455 2078
rect 18965 2075 19031 2078
rect 17217 2002 17283 2005
rect 11654 2000 17283 2002
rect 11654 1944 17222 2000
rect 17278 1944 17283 2000
rect 11654 1942 17283 1944
rect 17217 1939 17283 1942
rect 5717 1866 5783 1869
rect 11605 1866 11671 1869
rect 20713 1866 20779 1869
rect 5717 1864 11530 1866
rect 5717 1808 5722 1864
rect 5778 1808 11530 1864
rect 5717 1806 11530 1808
rect 5717 1803 5783 1806
rect 11470 1730 11530 1806
rect 11605 1864 20779 1866
rect 11605 1808 11610 1864
rect 11666 1808 20718 1864
rect 20774 1808 20779 1864
rect 11605 1806 20779 1808
rect 20854 1866 20914 2078
rect 27478 2032 27538 2350
rect 27478 1942 28000 2032
rect 27520 1912 28000 1942
rect 20854 1806 25698 1866
rect 11605 1803 11671 1806
rect 20713 1803 20779 1806
rect 15377 1730 15443 1733
rect 11470 1728 15443 1730
rect 11470 1672 15382 1728
rect 15438 1672 15443 1728
rect 11470 1670 15443 1672
rect 15377 1667 15443 1670
rect 17217 1730 17283 1733
rect 23749 1730 23815 1733
rect 17217 1728 23815 1730
rect 17217 1672 17222 1728
rect 17278 1672 23754 1728
rect 23810 1672 23815 1728
rect 17217 1670 23815 1672
rect 17217 1667 17283 1670
rect 23749 1667 23815 1670
rect 8753 1594 8819 1597
rect 14549 1594 14615 1597
rect 8753 1592 14615 1594
rect 8753 1536 8758 1592
rect 8814 1536 14554 1592
rect 14610 1536 14615 1592
rect 8753 1534 14615 1536
rect 8753 1531 8819 1534
rect 14549 1531 14615 1534
rect 17585 1594 17651 1597
rect 25497 1594 25563 1597
rect 17585 1592 25563 1594
rect 17585 1536 17590 1592
rect 17646 1536 25502 1592
rect 25558 1536 25563 1592
rect 17585 1534 25563 1536
rect 17585 1531 17651 1534
rect 25497 1531 25563 1534
rect 10961 1458 11027 1461
rect 18689 1458 18755 1461
rect 10961 1456 18755 1458
rect 10961 1400 10966 1456
rect 11022 1400 18694 1456
rect 18750 1400 18755 1456
rect 10961 1398 18755 1400
rect 25638 1458 25698 1806
rect 27520 1458 28000 1488
rect 25638 1398 28000 1458
rect 10961 1395 11027 1398
rect 18689 1395 18755 1398
rect 27520 1368 28000 1398
rect 15745 1050 15811 1053
rect 15745 1048 27538 1050
rect 15745 992 15750 1048
rect 15806 992 27538 1048
rect 15745 990 27538 992
rect 15745 987 15811 990
rect 27478 944 27538 990
rect 27478 854 28000 944
rect 27520 824 28000 854
rect 23933 370 23999 373
rect 27520 370 28000 400
rect 23933 368 28000 370
rect 23933 312 23938 368
rect 23994 312 28000 368
rect 23933 310 28000 312
rect 23933 307 23999 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 24716 13908 24780 13972
rect 14780 13772 14844 13836
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 16252 12548 16316 12612
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 16252 12336 16316 12340
rect 16252 12280 16266 12336
rect 16266 12280 16316 12336
rect 16252 12276 16316 12280
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 14780 10916 14844 10980
rect 23612 10916 23676 10980
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 23612 8120 23676 8124
rect 23612 8064 23662 8120
rect 23662 8064 23676 8120
rect 23612 8060 23676 8064
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 24716 3164 24780 3228
rect 24716 2892 24780 2956
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14779 13836 14845 13837
rect 14779 13772 14780 13836
rect 14844 13772 14845 13836
rect 14779 13771 14845 13772
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 14782 10981 14842 13771
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 16251 12612 16317 12613
rect 16251 12548 16252 12612
rect 16316 12548 16317 12612
rect 16251 12547 16317 12548
rect 16254 12341 16314 12547
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 16251 12340 16317 12341
rect 16251 12276 16252 12340
rect 16316 12276 16317 12340
rect 16251 12275 16317 12276
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14779 10980 14845 10981
rect 14779 10916 14780 10980
rect 14844 10916 14845 10980
rect 14779 10915 14845 10916
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24715 13972 24781 13973
rect 24715 13908 24716 13972
rect 24780 13908 24781 13972
rect 24715 13907 24781 13908
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 23611 10980 23677 10981
rect 23611 10916 23612 10980
rect 23676 10916 23677 10980
rect 23611 10915 23677 10916
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 23614 8125 23674 10915
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 23611 8124 23677 8125
rect 23611 8060 23612 8124
rect 23676 8060 23677 8124
rect 23611 8059 23677 8060
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24718 3229 24778 13907
rect 24715 3228 24781 3229
rect 24715 3164 24716 3228
rect 24780 3164 24781 3228
rect 24715 3163 24781 3164
rect 24718 2957 24778 3163
rect 24715 2956 24781 2957
rect 24715 2892 24716 2956
rect 24780 2892 24781 2956
rect 24715 2891 24781 2892
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _105_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_97 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10028 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_94
timestamp 1604681595
transform 1 0 9752 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 10304 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_104
timestamp 1604681595
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_106
timestamp 1604681595
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1604681595
transform 1 0 11040 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 12512 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1604681595
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_128
timestamp 1604681595
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_133
timestamp 1604681595
transform 1 0 13340 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12788 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14076 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13616 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1604681595
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604681595
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 16100 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_176
timestamp 1604681595
transform 1 0 17296 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1604681595
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1604681595
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1604681595
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16836 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1604681595
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1604681595
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1604681595
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18308 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18400 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19872 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19688 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_207
timestamp 1604681595
transform 1 0 20148 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_196
timestamp 1604681595
transform 1 0 19136 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_200
timestamp 1604681595
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_227
timestamp 1604681595
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_223
timestamp 1604681595
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_223
timestamp 1604681595
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_239
timestamp 1604681595
transform 1 0 23092 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_235
timestamp 1604681595
transform 1 0 22724 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_236
timestamp 1604681595
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 22908 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 22356 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1604681595
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_240
timestamp 1604681595
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_255
timestamp 1604681595
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_251
timestamp 1604681595
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1604681595
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_265
timestamp 1604681595
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1604681595
transform 1 0 25208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24932 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _042_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269
timestamp 1604681595
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 9844 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_99
timestamp 1604681595
transform 1 0 10212 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 10948 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12052 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1604681595
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_115
timestamp 1604681595
transform 1 0 11684 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1604681595
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_142
timestamp 1604681595
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_146
timestamp 1604681595
transform 1 0 14536 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_150
timestamp 1604681595
transform 1 0 14904 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 17756 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17204 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 1604681595
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_177
timestamp 1604681595
transform 1 0 17388 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_200
timestamp 1604681595
transform 1 0 19504 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_205
timestamp 1604681595
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 21344 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21068 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20516 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_209
timestamp 1604681595
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1604681595
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1604681595
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23828 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23276 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_243
timestamp 1604681595
transform 1 0 23460 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_266
timestamp 1604681595
transform 1 0 25576 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_274
timestamp 1604681595
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12052 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1604681595
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_114
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_118
timestamp 1604681595
transform 1 0 11960 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1604681595
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13984 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_138
timestamp 1604681595
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 15364 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16284 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_146
timestamp 1604681595
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_150
timestamp 1604681595
transform 1 0 14904 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_163
timestamp 1604681595
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16468 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18216 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_173
timestamp 1604681595
transform 1 0 17020 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604681595
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19780 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_195
timestamp 1604681595
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_199
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_212
timestamp 1604681595
transform 1 0 20608 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_217
timestamp 1604681595
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_221
timestamp 1604681595
transform 1 0 21436 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_236
timestamp 1604681595
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_240
timestamp 1604681595
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 25208 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_254
timestamp 1604681595
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_258
timestamp 1604681595
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_266
timestamp 1604681595
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_270
timestamp 1604681595
transform 1 0 25944 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1604681595
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_109
timestamp 1604681595
transform 1 0 11132 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_112
timestamp 1604681595
transform 1 0 11408 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_116
timestamp 1604681595
transform 1 0 11776 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_128
timestamp 1604681595
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_132
timestamp 1604681595
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 15732 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 15548 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1604681595
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1604681595
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_167
timestamp 1604681595
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_180
timestamp 1604681595
transform 1 0 17664 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_186
timestamp 1604681595
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18400 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19136 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 19504 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1604681595
transform 1 0 18952 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_198
timestamp 1604681595
transform 1 0 19320 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_210
timestamp 1604681595
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_224
timestamp 1604681595
transform 1 0 21712 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_229
timestamp 1604681595
transform 1 0 22172 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23276 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22356 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22724 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_233
timestamp 1604681595
transform 1 0 22540 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_237
timestamp 1604681595
transform 1 0 22908 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_260
timestamp 1604681595
transform 1 0 25024 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_272
timestamp 1604681595
transform 1 0 26128 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14260 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12696 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_139
timestamp 1604681595
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_162
timestamp 1604681595
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_166
timestamp 1604681595
transform 1 0 16376 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 19872 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1604681595
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1604681595
transform 1 0 19228 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_201
timestamp 1604681595
transform 1 0 19596 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21804 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_223
timestamp 1604681595
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_227
timestamp 1604681595
transform 1 0 21988 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_231
timestamp 1604681595
transform 1 0 22356 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1604681595
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_240
timestamp 1604681595
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 25208 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_254
timestamp 1604681595
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_258
timestamp 1604681595
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_266
timestamp 1604681595
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_270
timestamp 1604681595
transform 1 0 25944 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_276
timestamp 1604681595
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604681595
transform 1 0 11316 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604681595
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_114
timestamp 1604681595
transform 1 0 11592 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 12328 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_125
timestamp 1604681595
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12696 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13340 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_129
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_142
timestamp 1604681595
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_145
timestamp 1604681595
transform 1 0 14444 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_150
timestamp 1604681595
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1604681595
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_146
timestamp 1604681595
transform 1 0 14536 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 15272 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_162
timestamp 1604681595
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 1604681595
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15732 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_182
timestamp 1604681595
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18216 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 19596 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_205
timestamp 1604681595
transform 1 0 19964 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604681595
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_204
timestamp 1604681595
transform 1 0 19872 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20516 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_210
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_224
timestamp 1604681595
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_228
timestamp 1604681595
transform 1 0 22080 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_236
timestamp 1604681595
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_230
timestamp 1604681595
transform 1 0 22264 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_236
timestamp 1604681595
transform 1 0 22816 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22908 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1604681595
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_7_254
timestamp 1604681595
transform 1 0 24472 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_258
timestamp 1604681595
transform 1 0 24840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_259
timestamp 1604681595
transform 1 0 24932 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_266
timestamp 1604681595
transform 1 0 25576 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_262
timestamp 1604681595
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 25392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 25024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_268
timestamp 1604681595
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1604681595
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_272
timestamp 1604681595
transform 1 0 26128 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_276
timestamp 1604681595
transform 1 0 26496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11776 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_8_105
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_113
timestamp 1604681595
transform 1 0 11500 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_139
timestamp 1604681595
transform 1 0 13892 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_143
timestamp 1604681595
transform 1 0 14260 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 15640 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_149
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_161
timestamp 1604681595
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_165
timestamp 1604681595
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18216 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16652 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17664 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_182
timestamp 1604681595
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 19780 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19228 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_195
timestamp 1604681595
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_199
timestamp 1604681595
transform 1 0 19412 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1604681595
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_210
timestamp 1604681595
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_224
timestamp 1604681595
transform 1 0 21712 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23184 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_236
timestamp 1604681595
transform 1 0 22816 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_249
timestamp 1604681595
transform 1 0 24012 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 24748 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1604681595
transform 1 0 24380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_266
timestamp 1604681595
transform 1 0 25576 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp 1604681595
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1604681595
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604681595
transform 1 0 12512 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1604681595
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_127
timestamp 1604681595
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_131
timestamp 1604681595
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_154
timestamp 1604681595
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_158
timestamp 1604681595
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18124 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_171
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1604681595
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1604681595
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_204
timestamp 1604681595
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 22172 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 20608 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1604681595
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1604681595
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23276 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_233
timestamp 1604681595
transform 1 0 22540 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1604681595
transform 1 0 22908 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1604681595
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 25208 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604681595
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_254
timestamp 1604681595
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_258
timestamp 1604681595
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_266
timestamp 1604681595
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_270
timestamp 1604681595
transform 1 0 25944 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_276
timestamp 1604681595
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604681595
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13340 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_129
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_142
timestamp 1604681595
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_146
timestamp 1604681595
transform 1 0 14536 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1604681595
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_163
timestamp 1604681595
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16928 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_167
timestamp 1604681595
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_171
timestamp 1604681595
transform 1 0 16836 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 19412 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_191
timestamp 1604681595
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_195
timestamp 1604681595
transform 1 0 19044 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_202
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_210
timestamp 1604681595
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_224
timestamp 1604681595
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_228
timestamp 1604681595
transform 1 0 22080 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23276 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22724 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_234
timestamp 1604681595
transform 1 0 22632 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_237
timestamp 1604681595
transform 1 0 22908 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 25208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_260
timestamp 1604681595
transform 1 0 25024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_264
timestamp 1604681595
transform 1 0 25392 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_272
timestamp 1604681595
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_110
timestamp 1604681595
transform 1 0 11224 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1604681595
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1604681595
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1604681595
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13708 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13156 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_133
timestamp 1604681595
transform 1 0 13340 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_156
timestamp 1604681595
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_160
timestamp 1604681595
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_173
timestamp 1604681595
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp 1604681595
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1604681595
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18860 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_189
timestamp 1604681595
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_202
timestamp 1604681595
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_206
timestamp 1604681595
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20424 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_11_229
timestamp 1604681595
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_233
timestamp 1604681595
transform 1 0 22540 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_237
timestamp 1604681595
transform 1 0 22908 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 25576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1604681595
transform 1 0 25392 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_268
timestamp 1604681595
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_272
timestamp 1604681595
transform 1 0 26128 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_276
timestamp 1604681595
transform 1 0 26496 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11316 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_107
timestamp 1604681595
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_130
timestamp 1604681595
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_134
timestamp 1604681595
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_142
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16284 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15916 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_146
timestamp 1604681595
transform 1 0 14536 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_150
timestamp 1604681595
transform 1 0 14904 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp 1604681595
transform 1 0 15548 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1604681595
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_184
timestamp 1604681595
transform 1 0 18032 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1604681595
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1604681595
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21804 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_210
timestamp 1604681595
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_219
timestamp 1604681595
transform 1 0 21252 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_223
timestamp 1604681595
transform 1 0 21620 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23736 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24104 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_244
timestamp 1604681595
transform 1 0 23552 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_248
timestamp 1604681595
transform 1 0 23920 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24564 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_252
timestamp 1604681595
transform 1 0 24288 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_264
timestamp 1604681595
transform 1 0 25392 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_272
timestamp 1604681595
transform 1 0 26128 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_101
timestamp 1604681595
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1604681595
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_97
timestamp 1604681595
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_94
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_124
timestamp 1604681595
transform 1 0 12512 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604681595
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_14_129
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12788 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_141
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_140
timestamp 1604681595
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_136
timestamp 1604681595
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14352 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_150
timestamp 1604681595
transform 1 0 14904 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_146
timestamp 1604681595
transform 1 0 14536 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_153
timestamp 1604681595
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_157
timestamp 1604681595
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15916 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15640 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_171
timestamp 1604681595
transform 1 0 16836 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_167
timestamp 1604681595
transform 1 0 16468 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_174
timestamp 1604681595
transform 1 0 17112 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_170
timestamp 1604681595
transform 1 0 16744 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17020 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17204 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_184
timestamp 1604681595
transform 1 0 18032 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_177
timestamp 1604681595
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 18400 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 18492 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_191
timestamp 1604681595
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_188
timestamp 1604681595
transform 1 0 18400 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_191
timestamp 1604681595
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_195
timestamp 1604681595
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_195
timestamp 1604681595
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1604681595
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19412 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1604681595
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1604681595
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_224
timestamp 1604681595
transform 1 0 21712 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_222
timestamp 1604681595
transform 1 0 21528 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_229
timestamp 1604681595
transform 1 0 22172 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_236
timestamp 1604681595
transform 1 0 22816 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1604681595
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22356 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 22540 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_240
timestamp 1604681595
transform 1 0 23184 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604681595
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23552 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23736 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604681595
transform 1 0 25116 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_265
timestamp 1604681595
transform 1 0 25484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1604681595
transform 1 0 24380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_257
timestamp 1604681595
transform 1 0 24748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_264
timestamp 1604681595
transform 1 0 25392 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_272
timestamp 1604681595
transform 1 0 26128 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1604681595
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_82
timestamp 1604681595
transform 1 0 8648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9476 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_87
timestamp 1604681595
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14444 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_140
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_164
timestamp 1604681595
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_168
timestamp 1604681595
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18860 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_188
timestamp 1604681595
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_192
timestamp 1604681595
transform 1 0 18768 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1604681595
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_216
timestamp 1604681595
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_229
timestamp 1604681595
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23828 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_233
timestamp 1604681595
transform 1 0 22540 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_237
timestamp 1604681595
transform 1 0 22908 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604681595
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604681595
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_266
timestamp 1604681595
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_270
timestamp 1604681595
transform 1 0 25944 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_276
timestamp 1604681595
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 9936 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10396 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_99
timestamp 1604681595
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_103
timestamp 1604681595
transform 1 0 10580 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12512 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10948 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_116
timestamp 1604681595
transform 1 0 11776 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_120
timestamp 1604681595
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_143
timestamp 1604681595
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15456 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_147
timestamp 1604681595
transform 1 0 14628 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_165
timestamp 1604681595
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17020 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_169
timestamp 1604681595
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_182
timestamp 1604681595
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_186
timestamp 1604681595
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_199
timestamp 1604681595
transform 1 0 19412 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_203
timestamp 1604681595
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_207
timestamp 1604681595
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 22080 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21344 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20332 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_211
timestamp 1604681595
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_218
timestamp 1604681595
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_222
timestamp 1604681595
transform 1 0 21528 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23460 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_237
timestamp 1604681595
transform 1 0 22908 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_241
timestamp 1604681595
transform 1 0 23276 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 25208 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_254
timestamp 1604681595
transform 1 0 24472 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_258
timestamp 1604681595
transform 1 0 24840 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_266
timestamp 1604681595
transform 1 0 25576 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1604681595
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_11
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_23
timestamp 1604681595
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_35
timestamp 1604681595
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_47
timestamp 1604681595
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9200 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_97
timestamp 1604681595
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1604681595
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_127
timestamp 1604681595
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_131
timestamp 1604681595
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_144
timestamp 1604681595
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15088 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_148
timestamp 1604681595
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 17572 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_171
timestamp 1604681595
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1604681595
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18584 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21068 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_209
timestamp 1604681595
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_213
timestamp 1604681595
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24012 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23828 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604681595
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604681595
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 25576 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_258
timestamp 1604681595
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_262
timestamp 1604681595
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_22
timestamp 1604681595
transform 1 0 3128 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1604681595
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10304 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9936 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_98
timestamp 1604681595
transform 1 0 10120 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_123
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16836 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17848 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_168
timestamp 1604681595
transform 1 0 16560 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_180
timestamp 1604681595
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_184
timestamp 1604681595
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 18952 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_188
timestamp 1604681595
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_192
timestamp 1604681595
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1604681595
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_210
timestamp 1604681595
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 21160 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_225
timestamp 1604681595
transform 1 0 21804 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1604681595
transform 1 0 21436 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 21620 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 22172 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_248
timestamp 1604681595
transform 1 0 23920 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24656 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24472 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_252
timestamp 1604681595
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_265
timestamp 1604681595
transform 1 0 25484 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_273
timestamp 1604681595
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9476 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_96
timestamp 1604681595
transform 1 0 9936 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_97
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10304 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_123
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_119
timestamp 1604681595
transform 1 0 12052 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13708 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12788 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_129
timestamp 1604681595
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_133
timestamp 1604681595
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_147
timestamp 1604681595
transform 1 0 14628 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_163
timestamp 1604681595
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_164
timestamp 1604681595
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1604681595
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_156
timestamp 1604681595
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16836 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_168
timestamp 1604681595
transform 1 0 16560 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1604681595
transform 1 0 18952 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1604681595
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_195
timestamp 1604681595
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_190
timestamp 1604681595
transform 1 0 18584 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19136 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 18768 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_204
timestamp 1604681595
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19320 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19412 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_208
timestamp 1604681595
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_218
timestamp 1604681595
transform 1 0 21160 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_212
timestamp 1604681595
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604681595
transform 1 0 20976 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_223
timestamp 1604681595
transform 1 0 21620 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_223
timestamp 1604681595
transform 1 0 21620 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_219
timestamp 1604681595
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21804 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21988 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 22080 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 24104 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_247
timestamp 1604681595
transform 1 0 23828 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24564 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 25944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_264
timestamp 1604681595
transform 1 0 25392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_268
timestamp 1604681595
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_252
timestamp 1604681595
transform 1 0 24288 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_264
timestamp 1604681595
transform 1 0 25392 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 26312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_272
timestamp 1604681595
transform 1 0 26128 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_276
timestamp 1604681595
transform 1 0 26496 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_272
timestamp 1604681595
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_86
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_94
timestamp 1604681595
transform 1 0 9752 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1604681595
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 12512 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12052 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1604681595
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_116
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1604681595
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13524 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 13340 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12972 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_127
timestamp 1604681595
transform 1 0 12788 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_131
timestamp 1604681595
transform 1 0 13156 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_154
timestamp 1604681595
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1604681595
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1604681595
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18216 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18952 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18768 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_188
timestamp 1604681595
transform 1 0 18400 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 21804 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_213
timestamp 1604681595
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1604681595
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1604681595
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 24104 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_234
timestamp 1604681595
transform 1 0 22632 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_249
timestamp 1604681595
transform 1 0 24012 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_101
timestamp 1604681595
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12052 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_111
timestamp 1604681595
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_115
timestamp 1604681595
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_128
timestamp 1604681595
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1604681595
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_163
timestamp 1604681595
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 17756 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 17572 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17020 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_167
timestamp 1604681595
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_171
timestamp 1604681595
transform 1 0 16836 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_175
timestamp 1604681595
transform 1 0 17204 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_200
timestamp 1604681595
transform 1 0 19504 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21896 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1604681595
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_224
timestamp 1604681595
transform 1 0 21712 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_228
timestamp 1604681595
transform 1 0 22080 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22448 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23828 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22264 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23184 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_238
timestamp 1604681595
transform 1 0 23000 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_242
timestamp 1604681595
transform 1 0 23368 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 25392 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 24840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_256
timestamp 1604681595
transform 1 0 24656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_260
timestamp 1604681595
transform 1 0 25024 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_267
timestamp 1604681595
transform 1 0 25668 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604681595
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_98
timestamp 1604681595
transform 1 0 10120 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 11316 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_105
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13892 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_126
timestamp 1604681595
transform 1 0 12696 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_136
timestamp 1604681595
transform 1 0 13616 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15456 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_148
timestamp 1604681595
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_152
timestamp 1604681595
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19872 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_193
timestamp 1604681595
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_197
timestamp 1604681595
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_201
timestamp 1604681595
transform 1 0 19596 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21436 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_213
timestamp 1604681595
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_217
timestamp 1604681595
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_234
timestamp 1604681595
transform 1 0 22632 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_230
timestamp 1604681595
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23828 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 24012 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_23_268
timestamp 1604681595
transform 1 0 25760 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_276
timestamp 1604681595
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10580 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_101
timestamp 1604681595
transform 1 0 10396 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12512 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_122
timestamp 1604681595
transform 1 0 12328 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13064 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_126
timestamp 1604681595
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_139
timestamp 1604681595
transform 1 0 13892 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1604681595
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16100 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 15640 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_147
timestamp 1604681595
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_160
timestamp 1604681595
transform 1 0 15824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 17664 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 17204 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_172
timestamp 1604681595
transform 1 0 16928 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_177
timestamp 1604681595
transform 1 0 17388 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1604681595
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_193
timestamp 1604681595
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21436 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_219
timestamp 1604681595
transform 1 0 21252 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23920 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23644 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_240
timestamp 1604681595
transform 1 0 23184 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_244
timestamp 1604681595
transform 1 0 23552 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_247
timestamp 1604681595
transform 1 0 23828 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 24932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_257
timestamp 1604681595
transform 1 0 24748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_261
timestamp 1604681595
transform 1 0 25116 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_273
timestamp 1604681595
transform 1 0 26220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1604681595
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 14168 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_132
timestamp 1604681595
transform 1 0 13248 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_138
timestamp 1604681595
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_161
timestamp 1604681595
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_165
timestamp 1604681595
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1604681595
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19688 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1604681595
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_197
timestamp 1604681595
transform 1 0 19228 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 22080 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1604681595
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_225
timestamp 1604681595
transform 1 0 21804 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22264 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_254
timestamp 1604681595
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_258
timestamp 1604681595
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_268
timestamp 1604681595
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_272
timestamp 1604681595
transform 1 0 26128 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_276
timestamp 1604681595
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1604681595
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1604681595
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_94
timestamp 1604681595
transform 1 0 9752 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_103
timestamp 1604681595
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_103
timestamp 1604681595
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_107
timestamp 1604681595
transform 1 0 10948 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_107
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1604681595
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12052 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11132 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_128
timestamp 1604681595
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_132
timestamp 1604681595
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp 1604681595
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1604681595
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_150
timestamp 1604681595
transform 1 0 14904 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_154
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_161
timestamp 1604681595
transform 1 0 15916 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_157
timestamp 1604681595
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15456 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16008 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15640 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1604681595
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_171
timestamp 1604681595
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_171
timestamp 1604681595
transform 1 0 16836 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_167
timestamp 1604681595
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17020 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 17204 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1604681595
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_184
timestamp 1604681595
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18216 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_195
timestamp 1604681595
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_188
timestamp 1604681595
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18768 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_203
timestamp 1604681595
transform 1 0 19780 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_199
timestamp 1604681595
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_205
timestamp 1604681595
transform 1 0 19964 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_201
timestamp 1604681595
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19780 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 22172 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1604681595
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_224
timestamp 1604681595
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_228
timestamp 1604681595
transform 1 0 22080 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_227
timestamp 1604681595
transform 1 0 21988 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_238
timestamp 1604681595
transform 1 0 23000 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_231
timestamp 1604681595
transform 1 0 22356 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_232
timestamp 1604681595
transform 1 0 22448 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22264 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 22540 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 22724 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 22724 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_258
timestamp 1604681595
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1604681595
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_254
timestamp 1604681595
transform 1 0 24472 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_266
timestamp 1604681595
transform 1 0 25576 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 25024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 25208 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_268
timestamp 1604681595
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_274
timestamp 1604681595
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_272
timestamp 1604681595
transform 1 0 26128 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_276
timestamp 1604681595
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10396 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 9292 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_88
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1604681595
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_97
timestamp 1604681595
transform 1 0 10028 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12052 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11500 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_110
timestamp 1604681595
transform 1 0 11224 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_115
timestamp 1604681595
transform 1 0 11684 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_128
timestamp 1604681595
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_132
timestamp 1604681595
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15732 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15456 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1604681595
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_158
timestamp 1604681595
transform 1 0 15640 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18216 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 17664 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_182
timestamp 1604681595
transform 1 0 17848 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20148 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_205
timestamp 1604681595
transform 1 0 19964 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20516 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_209
timestamp 1604681595
transform 1 0 20332 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1604681595
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23460 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23276 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22908 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_234
timestamp 1604681595
transform 1 0 22632 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 25024 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 24472 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24840 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_252
timestamp 1604681595
transform 1 0 24288 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_256
timestamp 1604681595
transform 1 0 24656 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_264
timestamp 1604681595
transform 1 0 25392 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_272
timestamp 1604681595
transform 1 0 26128 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 9292 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10304 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_92
timestamp 1604681595
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_96
timestamp 1604681595
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_109
timestamp 1604681595
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1604681595
transform 1 0 11500 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13800 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_129
timestamp 1604681595
transform 1 0 12972 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_134
timestamp 1604681595
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15364 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_147
timestamp 1604681595
transform 1 0 14628 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_151
timestamp 1604681595
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_164
timestamp 1604681595
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1604681595
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_168
timestamp 1604681595
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 16928 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1604681595
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18308 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_206
timestamp 1604681595
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 21160 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 20608 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 21712 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22080 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 20976 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1604681595
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_214
timestamp 1604681595
transform 1 0 20792 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1604681595
transform 1 0 21528 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_226
timestamp 1604681595
transform 1 0 21896 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22264 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_236
timestamp 1604681595
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604681595
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1604681595
transform 1 0 25392 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_268
timestamp 1604681595
transform 1 0 25760 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_276
timestamp 1604681595
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_73
timestamp 1604681595
transform 1 0 7820 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 9292 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1604681595
transform 1 0 8924 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12144 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11960 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_112
timestamp 1604681595
transform 1 0 11408 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 14168 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13708 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_135
timestamp 1604681595
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_139
timestamp 1604681595
transform 1 0 13892 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_145
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_149
timestamp 1604681595
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_163
timestamp 1604681595
transform 1 0 16100 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 17204 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 16928 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_168
timestamp 1604681595
transform 1 0 16560 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_184
timestamp 1604681595
transform 1 0 18032 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18860 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_189
timestamp 1604681595
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 21436 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 21068 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_210
timestamp 1604681595
transform 1 0 20424 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_219
timestamp 1604681595
transform 1 0 21252 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_225
timestamp 1604681595
transform 1 0 21804 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 22540 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23460 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_237
timestamp 1604681595
transform 1 0 22908 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_241
timestamp 1604681595
transform 1 0 23276 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 25208 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24656 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_254
timestamp 1604681595
transform 1 0 24472 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_258
timestamp 1604681595
transform 1 0 24840 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_266
timestamp 1604681595
transform 1 0 25576 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_274
timestamp 1604681595
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_68
timestamp 1604681595
transform 1 0 7360 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_90
timestamp 1604681595
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_94
timestamp 1604681595
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11868 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_107
timestamp 1604681595
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_111
timestamp 1604681595
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_115
timestamp 1604681595
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1604681595
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13340 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_129
timestamp 1604681595
transform 1 0 12972 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_152
timestamp 1604681595
transform 1 0 15088 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_156
timestamp 1604681595
transform 1 0 15456 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_162
timestamp 1604681595
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1604681595
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1604681595
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 19780 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_193
timestamp 1604681595
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1604681595
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_201
timestamp 1604681595
transform 1 0 19596 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_206
timestamp 1604681595
transform 1 0 20056 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20792 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 21804 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22172 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_210
timestamp 1604681595
transform 1 0 20424 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_223
timestamp 1604681595
transform 1 0 21620 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_227
timestamp 1604681595
transform 1 0 21988 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_231
timestamp 1604681595
transform 1 0 22356 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1604681595
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1604681595
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_264
timestamp 1604681595
transform 1 0 25392 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_276
timestamp 1604681595
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10580 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_97
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_101
timestamp 1604681595
transform 1 0 10396 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_122
timestamp 1604681595
transform 1 0 12328 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13340 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_128
timestamp 1604681595
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_132
timestamp 1604681595
transform 1 0 13248 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_142
timestamp 1604681595
transform 1 0 14168 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_146
timestamp 1604681595
transform 1 0 14536 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1604681595
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 17756 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17204 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17572 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1604681595
transform 1 0 17020 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_177
timestamp 1604681595
transform 1 0 17388 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19320 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 18768 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19136 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_190
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1604681595
transform 1 0 18952 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_204
timestamp 1604681595
transform 1 0 19872 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23368 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23184 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22816 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_234
timestamp 1604681595
transform 1 0 22632 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_238
timestamp 1604681595
transform 1 0 23000 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25300 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_261
timestamp 1604681595
transform 1 0 25116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_265
timestamp 1604681595
transform 1 0 25484 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_273
timestamp 1604681595
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_72
timestamp 1604681595
transform 1 0 7728 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_70
timestamp 1604681595
transform 1 0 7544 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_82
timestamp 1604681595
transform 1 0 8648 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_79
timestamp 1604681595
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_75
timestamp 1604681595
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_33_83
timestamp 1604681595
transform 1 0 8740 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_89
timestamp 1604681595
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_102
timestamp 1604681595
transform 1 0 10488 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_102
timestamp 1604681595
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_106
timestamp 1604681595
transform 1 0 10856 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_106
timestamp 1604681595
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11224 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_125
timestamp 1604681595
transform 1 0 12604 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_122
timestamp 1604681595
transform 1 0 12328 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_116
timestamp 1604681595
transform 1 0 11776 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13064 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12880 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_142
timestamp 1604681595
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_139
timestamp 1604681595
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_143
timestamp 1604681595
transform 1 0 14260 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_150
timestamp 1604681595
transform 1 0 14904 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_146
timestamp 1604681595
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15456 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 14628 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_158
timestamp 1604681595
transform 1 0 15640 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15916 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16100 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14904 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_33_173
timestamp 1604681595
transform 1 0 17020 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1604681595
transform 1 0 16652 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16836 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_186
timestamp 1604681595
transform 1 0 18216 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_182
timestamp 1604681595
transform 1 0 17848 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1604681595
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 18032 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 18400 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_207
timestamp 1604681595
transform 1 0 20148 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_203
timestamp 1604681595
transform 1 0 19780 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_199
timestamp 1604681595
transform 1 0 19412 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_207
timestamp 1604681595
transform 1 0 20148 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_203
timestamp 1604681595
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19596 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19964 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_210
timestamp 1604681595
transform 1 0 20424 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_211
timestamp 1604681595
transform 1 0 20516 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20700 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_34_224
timestamp 1604681595
transform 1 0 21712 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_228
timestamp 1604681595
transform 1 0 22080 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_224
timestamp 1604681595
transform 1 0 21712 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21896 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_236
timestamp 1604681595
transform 1 0 22816 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1604681595
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 22448 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_240
timestamp 1604681595
transform 1 0 23184 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604681595
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23368 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23552 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_34_253
timestamp 1604681595
transform 1 0 24380 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_258
timestamp 1604681595
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_254
timestamp 1604681595
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_265
timestamp 1604681595
transform 1 0 25484 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 25116 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_268
timestamp 1604681595
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 25944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_272
timestamp 1604681595
transform 1 0 26128 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_276
timestamp 1604681595
transform 1 0 26496 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_273
timestamp 1604681595
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604681595
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8188 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_74
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10488 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_96
timestamp 1604681595
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_100
timestamp 1604681595
transform 1 0 10304 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_113
timestamp 1604681595
transform 1 0 11500 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 1604681595
transform 1 0 12052 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13248 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13064 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12696 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14260 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_128
timestamp 1604681595
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_141
timestamp 1604681595
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_145
timestamp 1604681595
transform 1 0 14444 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_158
timestamp 1604681595
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_162
timestamp 1604681595
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1604681595
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1604681595
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19964 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19596 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_193
timestamp 1604681595
transform 1 0 18860 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_199
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_203
timestamp 1604681595
transform 1 0 19780 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_207
timestamp 1604681595
transform 1 0 20148 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20516 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20332 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23920 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_230
timestamp 1604681595
transform 1 0 22264 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_234
timestamp 1604681595
transform 1 0 22632 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 25024 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_254
timestamp 1604681595
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_258
timestamp 1604681595
transform 1 0 24840 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_268
timestamp 1604681595
transform 1 0 25760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_272
timestamp 1604681595
transform 1 0 26128 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_276
timestamp 1604681595
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604681595
transform 1 0 8556 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8188 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_68
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_76
timestamp 1604681595
transform 1 0 8096 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_79
timestamp 1604681595
transform 1 0 8372 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_84
timestamp 1604681595
transform 1 0 8832 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604681595
transform 1 0 12236 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_112
timestamp 1604681595
transform 1 0 11408 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_120
timestamp 1604681595
transform 1 0 12144 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_124
timestamp 1604681595
transform 1 0 12512 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13248 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12880 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_130
timestamp 1604681595
transform 1 0 13064 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_141
timestamp 1604681595
transform 1 0 14076 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14812 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16008 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16376 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_147
timestamp 1604681595
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_151
timestamp 1604681595
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_160
timestamp 1604681595
transform 1 0 15824 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_164
timestamp 1604681595
transform 1 0 16192 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 18032 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_168
timestamp 1604681595
transform 1 0 16560 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1604681595
transform 1 0 17664 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_186
timestamp 1604681595
transform 1 0 18216 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20240 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19044 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_194
timestamp 1604681595
transform 1 0 18952 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_206
timestamp 1604681595
transform 1 0 20056 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_210
timestamp 1604681595
transform 1 0 20424 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23736 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_234
timestamp 1604681595
transform 1 0 22632 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 25024 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_252
timestamp 1604681595
transform 1 0 24288 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_264
timestamp 1604681595
transform 1 0 25392 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_272
timestamp 1604681595
transform 1 0 26128 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1604681595
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1604681595
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1604681595
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604681595
transform 1 0 9752 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_97
timestamp 1604681595
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_101
timestamp 1604681595
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_114
timestamp 1604681595
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1604681595
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_142
timestamp 1604681595
transform 1 0 14168 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 14904 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_146
timestamp 1604681595
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16836 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1604681595
transform 1 0 16652 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_173
timestamp 1604681595
transform 1 0 17020 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_179
timestamp 1604681595
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_187
timestamp 1604681595
transform 1 0 18308 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19044 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18492 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_191
timestamp 1604681595
transform 1 0 18676 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21528 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20976 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21344 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_214
timestamp 1604681595
transform 1 0 20792 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_218
timestamp 1604681595
transform 1 0 21160 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 22540 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22908 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_231
timestamp 1604681595
transform 1 0 22356 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_235
timestamp 1604681595
transform 1 0 22724 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_239
timestamp 1604681595
transform 1 0 23092 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 24932 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 25484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 25852 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_251
timestamp 1604681595
transform 1 0 24196 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_255
timestamp 1604681595
transform 1 0 24564 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_263
timestamp 1604681595
transform 1 0 25300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_267
timestamp 1604681595
transform 1 0 25668 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_271
timestamp 1604681595
transform 1 0 26036 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10396 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10212 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12328 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_120
timestamp 1604681595
transform 1 0 12144 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_124
timestamp 1604681595
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1604681595
transform 1 0 14076 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_137
timestamp 1604681595
transform 1 0 13708 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_143
timestamp 1604681595
transform 1 0 14260 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15456 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1604681595
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_154
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 17940 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17572 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_175
timestamp 1604681595
transform 1 0 17204 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_181
timestamp 1604681595
transform 1 0 17756 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 18952 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_192
timestamp 1604681595
transform 1 0 18768 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_196
timestamp 1604681595
transform 1 0 19136 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_206
timestamp 1604681595
transform 1 0 20056 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21896 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_224
timestamp 1604681595
transform 1 0 21712 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_228
timestamp 1604681595
transform 1 0 22080 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22448 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23736 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22264 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_238
timestamp 1604681595
transform 1 0 23000 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 25024 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_252
timestamp 1604681595
transform 1 0 24288 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_264
timestamp 1604681595
transform 1 0 25392 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_272
timestamp 1604681595
transform 1 0 26128 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1604681595
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604681595
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1604681595
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604681595
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604681595
transform 1 0 12604 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_110
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_117
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_133
timestamp 1604681595
transform 1 0 13340 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_129
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_133
timestamp 1604681595
transform 1 0 13340 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_129
timestamp 1604681595
transform 1 0 12972 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1604681595
transform 1 0 13156 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604681595
transform 1 0 13064 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_145
timestamp 1604681595
transform 1 0 14444 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_137
timestamp 1604681595
transform 1 0 13708 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13892 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604681595
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14076 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16008 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16376 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_160
timestamp 1604681595
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_164
timestamp 1604681595
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_163
timestamp 1604681595
transform 1 0 16100 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_176
timestamp 1604681595
transform 1 0 17296 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_170
timestamp 1604681595
transform 1 0 16744 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_167
timestamp 1604681595
transform 1 0 16468 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_174
timestamp 1604681595
transform 1 0 17112 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16560 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17388 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16560 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_181
timestamp 1604681595
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_178
timestamp 1604681595
transform 1 0 17480 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17572 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604681595
transform 1 0 19136 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1604681595
transform 1 0 19964 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_203
timestamp 1604681595
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_207
timestamp 1604681595
transform 1 0 20148 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_188
timestamp 1604681595
transform 1 0 18400 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1604681595
transform 1 0 18768 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_200
timestamp 1604681595
transform 1 0 19504 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_212
timestamp 1604681595
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_215
timestamp 1604681595
transform 1 0 20884 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604681595
transform 1 0 21068 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 20516 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_229
timestamp 1604681595
transform 1 0 22172 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_223
timestamp 1604681595
transform 1 0 21620 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_219
timestamp 1604681595
transform 1 0 21252 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604681595
transform 1 0 21436 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_219
timestamp 1604681595
transform 1 0 21252 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_235
timestamp 1604681595
transform 1 0 22724 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1604681595
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604681595
transform 1 0 22264 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604681595
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 22356 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 23460 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_247
timestamp 1604681595
transform 1 0 23828 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_249
timestamp 1604681595
transform 1 0 24012 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604681595
transform 1 0 23828 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_259
timestamp 1604681595
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_263
timestamp 1604681595
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_259
timestamp 1604681595
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_275
timestamp 1604681595
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1604681595
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604681595
transform 1 0 14168 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_135
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_141
timestamp 1604681595
transform 1 0 14076 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604681595
transform 1 0 15272 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1604681595
transform 1 0 15824 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1604681595
transform 1 0 14720 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1604681595
transform 1 0 16376 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_146
timestamp 1604681595
transform 1 0 14536 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_150
timestamp 1604681595
transform 1 0 14904 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_158
timestamp 1604681595
transform 1 0 15640 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_162
timestamp 1604681595
transform 1 0 16008 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 16836 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1604681595
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_168
timestamp 1604681595
transform 1 0 16560 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_175
timestamp 1604681595
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_179
timestamp 1604681595
transform 1 0 17572 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_192
timestamp 1604681595
transform 1 0 18768 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_188
timestamp 1604681595
transform 1 0 18400 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_195
timestamp 1604681595
transform 1 0 19044 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_200
timestamp 1604681595
transform 1 0 19504 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_204
timestamp 1604681595
transform 1 0 19872 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 19964 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_207
timestamp 1604681595
transform 1 0 20148 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604681595
transform 1 0 21896 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604681595
transform 1 0 20792 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_212
timestamp 1604681595
transform 1 0 20608 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_216
timestamp 1604681595
transform 1 0 20976 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_224
timestamp 1604681595
transform 1 0 21712 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_228
timestamp 1604681595
transform 1 0 22080 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604681595
transform 1 0 22264 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_236
timestamp 1604681595
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_240
timestamp 1604681595
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 24564 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604681595
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_259
timestamp 1604681595
transform 1 0 24932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_263
timestamp 1604681595
transform 1 0 25300 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_275
timestamp 1604681595
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_56
timestamp 1604681595
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604681595
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604681595
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604681595
transform 1 0 16376 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_164
timestamp 1604681595
transform 1 0 16192 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_170
timestamp 1604681595
transform 1 0 16744 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_182
timestamp 1604681595
transform 1 0 17848 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 18860 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 19964 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_197
timestamp 1604681595
transform 1 0 19228 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_201
timestamp 1604681595
transform 1 0 19596 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 21436 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_209
timestamp 1604681595
transform 1 0 20332 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_225
timestamp 1604681595
transform 1 0 21804 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 22632 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_233
timestamp 1604681595
transform 1 0 22540 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_238
timestamp 1604681595
transform 1 0 23000 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_246
timestamp 1604681595
transform 1 0 23736 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 24564 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_259
timestamp 1604681595
transform 1 0 24932 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_271
timestamp 1604681595
transform 1 0 26036 0 -1 25568
box -38 -48 590 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal3 s 0 13880 480 14000 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 23264 480 23384 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 27520 4904 28000 5024 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 27520 10752 28000 10872 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 27520 11296 28000 11416 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 27520 5448 28000 5568 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 27520 6672 28000 6792 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 27520 7216 28000 7336 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 27520 7760 28000 7880 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 27520 8984 28000 9104 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 27520 9528 28000 9648 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 27520 10072 28000 10192 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 27520 22992 28000 23112 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 27520 23536 28000 23656 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 27520 24080 28000 24200 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 27520 24760 28000 24880 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 27520 25848 28000 25968 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 27520 26528 28000 26648 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 27520 27072 28000 27192 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 27520 27616 28000 27736 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 27520 17144 28000 17264 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 27520 17688 28000 17808 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 27520 18368 28000 18488 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 27520 18912 28000 19032 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 27520 19456 28000 19576 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 27520 20680 28000 20800 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 27520 21224 28000 21344 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 27520 21768 28000 21888 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1582 0 1638 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3698 0 3754 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 22742 0 22798 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 24122 0 24178 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 25502 0 25558 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 26146 0 26202 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 26882 0 26938 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 27526 0 27582 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 15290 0 15346 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 20074 0 20130 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal2 s 938 27520 994 28000 6 chany_top_in[0]
port 83 nsew default input
rlabel metal2 s 7746 27520 7802 28000 6 chany_top_in[10]
port 84 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[11]
port 85 nsew default input
rlabel metal2 s 9126 27520 9182 28000 6 chany_top_in[12]
port 86 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[13]
port 87 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[14]
port 88 nsew default input
rlabel metal2 s 11150 27520 11206 28000 6 chany_top_in[15]
port 89 nsew default input
rlabel metal2 s 11886 27520 11942 28000 6 chany_top_in[16]
port 90 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[17]
port 91 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 chany_top_in[18]
port 92 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[19]
port 93 nsew default input
rlabel metal2 s 1582 27520 1638 28000 6 chany_top_in[1]
port 94 nsew default input
rlabel metal2 s 2318 27520 2374 28000 6 chany_top_in[2]
port 95 nsew default input
rlabel metal2 s 2962 27520 3018 28000 6 chany_top_in[3]
port 96 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 chany_top_in[4]
port 97 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 chany_top_in[5]
port 98 nsew default input
rlabel metal2 s 4986 27520 5042 28000 6 chany_top_in[6]
port 99 nsew default input
rlabel metal2 s 5722 27520 5778 28000 6 chany_top_in[7]
port 100 nsew default input
rlabel metal2 s 6366 27520 6422 28000 6 chany_top_in[8]
port 101 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[9]
port 102 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_out[0]
port 103 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[10]
port 104 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[11]
port 105 nsew default tristate
rlabel metal2 s 22742 27520 22798 28000 6 chany_top_out[12]
port 106 nsew default tristate
rlabel metal2 s 23478 27520 23534 28000 6 chany_top_out[13]
port 107 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[14]
port 108 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 109 nsew default tristate
rlabel metal2 s 25502 27520 25558 28000 6 chany_top_out[16]
port 110 nsew default tristate
rlabel metal2 s 26146 27520 26202 28000 6 chany_top_out[17]
port 111 nsew default tristate
rlabel metal2 s 26882 27520 26938 28000 6 chany_top_out[18]
port 112 nsew default tristate
rlabel metal2 s 27526 27520 27582 28000 6 chany_top_out[19]
port 113 nsew default tristate
rlabel metal2 s 15290 27520 15346 28000 6 chany_top_out[1]
port 114 nsew default tristate
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_out[2]
port 115 nsew default tristate
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[3]
port 116 nsew default tristate
rlabel metal2 s 17314 27520 17370 28000 6 chany_top_out[4]
port 117 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[5]
port 118 nsew default tristate
rlabel metal2 s 18694 27520 18750 28000 6 chany_top_out[6]
port 119 nsew default tristate
rlabel metal2 s 19338 27520 19394 28000 6 chany_top_out[7]
port 120 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[8]
port 121 nsew default tristate
rlabel metal2 s 20718 27520 20774 28000 6 chany_top_out[9]
port 122 nsew default tristate
rlabel metal3 s 0 4632 480 4752 6 prog_clk
port 123 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_34_
port 124 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_bottom_grid_pin_35_
port 125 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_36_
port 126 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 right_bottom_grid_pin_37_
port 127 nsew default input
rlabel metal3 s 27520 2592 28000 2712 6 right_bottom_grid_pin_38_
port 128 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 right_bottom_grid_pin_39_
port 129 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 right_bottom_grid_pin_40_
port 130 nsew default input
rlabel metal3 s 27520 4360 28000 4480 6 right_bottom_grid_pin_41_
port 131 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 133 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
