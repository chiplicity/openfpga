//
//
//
//
//
//
//
//
`timescale 1ns / 1ps

module top_top_formal_verification (
input [0:0] a_fm,
input [0:0] b_fm,
output [0:0] out:c_fm);

//
wire [0:0] prog_clk;
wire [0:0] Test_en;
wire [0:0] clk;
wire [0:7] gfpga_pad_GPIO_Y;
wire [0:7] gfpga_pad_GPIO_A;
wire [0:7] gfpga_pad_GPIO_IE;
wire [0:7] gfpga_pad_GPIO_OE;
wire [0:0] ccff_head;
wire [0:0] ccff_tail;

//
	fpga_top U0_formal_verification (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.clk(clk[0]),
		.gfpga_pad_GPIO_A(gfpga_pad_GPIO_A[0:7]),
		.gfpga_pad_GPIO_IE(gfpga_pad_GPIO_IE[0:7]),
		.gfpga_pad_GPIO_OE(gfpga_pad_GPIO_OE[0:7]),
		.gfpga_pad_GPIO_Y(gfpga_pad_GPIO_Y[0:7]),
		.ccff_head(ccff_head[0]),
		.ccff_tail(ccff_tail[0]));

//
	assign prog_clk[0] = 1'b0;
	assign Test_en[0] = 1'b0;
//

//
//
	assign gfpga_pad_GPIO_Y[4] = a_fm[0];
//
	assign gfpga_pad_GPIO_Y[6] = b_fm[0];
//
	assign out:c_fm[0] = gfpga_pad_GPIO_Y[5];

//
	assign gfpga_pad_GPIO_Y[0] = 1'b0;
	assign gfpga_pad_GPIO_Y[1] = 1'b0;
	assign gfpga_pad_GPIO_Y[2] = 1'b0;
	assign gfpga_pad_GPIO_Y[3] = 1'b0;
	assign gfpga_pad_GPIO_Y[7] = 1'b0;

//
`ifdef ICARUS_SIMULATOR
//
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = 17'b00000000110000001;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = 2'b01;
	assign U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16] = {17{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0] = 1'b0;
	assign U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0] = 1'b1;
	assign U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:2] = 3'b010;
	assign U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:2] = {3{1'b1}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:2] = 3'b110;
	assign U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__0_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:2] = 3'b010;
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:3] = 4'b0010;
	assign U0_formal_verification.sb_1__0_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_4.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_5.mem_out[0:4] = {5{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_1__1_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_1__2_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__0_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__1_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.sb_2__2_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_12.mem_out[0:3] = {4{1'b1}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_13.mem_out[0:3] = {4{1'b1}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_bottom_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__1_.mem_bottom_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_bottom_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b1}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__1_.mem_bottom_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_1__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	assign U0_formal_verification.cby_2__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
initial begin
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = 17'b11111111001111110;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16] = {17{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_14.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_3.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_5.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_10.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__0_.mem_right_track_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_3.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_5.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_3.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_5.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_7.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_3.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_5.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_7.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_11.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_13.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_15.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_12.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_13.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_bottom_ipin_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__1_.mem_bottom_ipin_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_15.mem_outb[0:3] = {4{1'b1}};
end
//
`else
//
initial begin
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], 17'b00000000110000001);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], 17'b11111111001111110);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], 2'b01);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], 2'b10);
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0:16], {17{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.ltile_clb_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0:16], {17{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.ltile_clb_frac_logic_0.mem_frac_logic_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_fabric_out_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.ltile_clb_md_fle_mp_fabric_0.mem_ff_0_D_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_1__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_top_2__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_right_3__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_out[0], 1'b1);
	$deposit(U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_sky130_fd_sc_hd__dfxbp_1_mem.mem_outb[0], 1'b0);
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_4.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_top_track_24.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:2], 3'b010);
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_0.mem_outb[0:2], 3'b101);
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_2.mem_outb[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:2], 3'b110);
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_4.mem_outb[0:2], 3'b001);
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_6.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_10.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_12.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_16.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_18.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_20.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_22.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_24.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__0_.mem_right_track_26.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_8.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_16.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_24.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_top_track_32.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_6.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_8.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_10.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_12.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_14.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_16.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_18.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_20.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_22.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_24.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_right_track_26.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:2], 3'b010);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_outb[0:2], 3'b101);
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_0.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_4.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_right_track_24.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_6.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_8.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_10.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_10.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_12.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_16.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_18.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_20.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_22.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_24.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_28.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_28.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_30.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_30.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_32.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_32.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_34.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_34.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_36.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_36.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_38.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_top_track_38.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:3], 4'b0010);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_0.mem_outb[0:3], 4'b1101);
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_4.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_16.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_24.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_right_track_32.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_5.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_17.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_25.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__0_.mem_left_track_33.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_4.mem_outb[0:4], {5{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_16.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_24.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_top_track_32.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_4.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_4.mem_outb[0:4], {5{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_16.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_24.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_24.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_right_track_32.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_5.mem_outb[0:4], {5{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_5.mem_out[0:4], {5{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_5.mem_outb[0:4], {5{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_17.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_25.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_25.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__1_.mem_left_track_33.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_8.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_16.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_24.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_32.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_right_track_32.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_19.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_21.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_23.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_27.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_29.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_29.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_31.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_31.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_35.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_35.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_37.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_37.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_39.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_bottom_track_39.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_9.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_17.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_25.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_1__2_.mem_left_track_33.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_0.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_2.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_4.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_6.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_8.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_10.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_12.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_14.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_16.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_18.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_18.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_20.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_20.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_22.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_22.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_24.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_24.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_26.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_26.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_28.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_28.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_30.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_30.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_32.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_32.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_34.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_34.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_36.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_36.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_38.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_top_track_38.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_7.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_19.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_21.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_23.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_25.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__0_.mem_left_track_27.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_4.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_16.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_24.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_24.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_32.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_top_track_32.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_5.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_7.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_9.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_11.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_11.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_13.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_13.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_15.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_15.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_19.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_21.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_23.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__1_.mem_left_track_25.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_out[0:2], {3{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_outb[0:2], {3{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_15.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_15.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_19.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_19.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_21.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_21.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_23.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_23.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_27.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_27.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_29.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_29.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_31.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_31.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_35.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_35.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_37.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_37.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_39.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_bottom_track_39.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_1.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_5.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_5.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_9.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_25.mem_out[0:1], {2{1'b0}});
	$deposit(U0_formal_verification.sb_2__2_.mem_left_track_25.mem_outb[0:1], {2{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_4.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_5.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_6.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_7.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_10.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_11.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_12.mem_out[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_12.mem_outb[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_13.mem_out[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_13.mem_outb[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_14.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_bottom_ipin_15.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_6.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_7.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_10.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_11.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_12.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_13.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_14.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__1_.mem_bottom_ipin_15.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_4.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_5.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_6.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_7.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_10.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_11.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_12.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_13.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_14.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_bottom_ipin_15.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_outb[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_4.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_5.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_6.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_7.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_10.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_11.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_12.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_13.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_14.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__1_.mem_bottom_ipin_15.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cbx_2__2_.mem_bottom_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_left_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_6.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_7.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_10.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_11.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_12.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_13.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_14.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__1_.mem_right_ipin_15.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_left_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_10.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_11.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_12.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_13.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_14.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_1__2_.mem_right_ipin_15.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_4.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_5.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_6.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_7.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_10.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_11.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_12.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_13.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_14.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__1_.mem_right_ipin_15.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_6.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_6.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_7.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_7.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_8.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_8.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_9.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_9.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_10.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_10.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_11.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_11.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_12.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_12.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_13.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_13.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_14.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_14.mem_outb[0:3], {4{1'b1}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_15.mem_out[0:3], {4{1'b0}});
	$deposit(U0_formal_verification.cby_2__2_.mem_right_ipin_15.mem_outb[0:3], {4{1'b1}});
end
//
`endif
//
endmodule
//

