magic
tech sky130A
magscale 1 2
timestamp 1605004234
<< locali >>
rect 6929 22491 6963 22593
rect 12449 17051 12483 17221
<< viali >>
rect 5273 25449 5307 25483
rect 8217 25449 8251 25483
rect 12633 25381 12667 25415
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 5181 25313 5215 25347
rect 6929 25313 6963 25347
rect 8033 25313 8067 25347
rect 8585 25313 8619 25347
rect 9781 25313 9815 25347
rect 5365 25245 5399 25279
rect 10885 25245 10919 25279
rect 1593 25177 1627 25211
rect 7113 25177 7147 25211
rect 9965 25177 9999 25211
rect 2697 25109 2731 25143
rect 3433 25109 3467 25143
rect 4813 25109 4847 25143
rect 5825 25109 5859 25143
rect 10793 25109 10827 25143
rect 4905 24905 4939 24939
rect 2697 24837 2731 24871
rect 8125 24837 8159 24871
rect 3893 24769 3927 24803
rect 3985 24769 4019 24803
rect 5733 24769 5767 24803
rect 6285 24769 6319 24803
rect 8861 24769 8895 24803
rect 10241 24769 10275 24803
rect 11345 24769 11379 24803
rect 11897 24769 11931 24803
rect 12265 24769 12299 24803
rect 12909 24769 12943 24803
rect 13093 24769 13127 24803
rect 1409 24701 1443 24735
rect 2329 24701 2363 24735
rect 3341 24701 3375 24735
rect 3801 24701 3835 24735
rect 5549 24701 5583 24735
rect 6837 24701 6871 24735
rect 7389 24701 7423 24735
rect 7941 24701 7975 24735
rect 8493 24701 8527 24735
rect 9045 24701 9079 24735
rect 12817 24701 12851 24735
rect 5641 24633 5675 24667
rect 6561 24633 6595 24667
rect 10609 24633 10643 24667
rect 11161 24633 11195 24667
rect 1593 24565 1627 24599
rect 2053 24565 2087 24599
rect 3433 24565 3467 24599
rect 4537 24565 4571 24599
rect 5181 24565 5215 24599
rect 7021 24565 7055 24599
rect 7849 24565 7883 24599
rect 9229 24565 9263 24599
rect 9781 24565 9815 24599
rect 10701 24565 10735 24599
rect 11069 24565 11103 24599
rect 12449 24565 12483 24599
rect 3525 24361 3559 24395
rect 7665 24361 7699 24395
rect 8125 24361 8159 24395
rect 10057 24361 10091 24395
rect 13093 24361 13127 24395
rect 14197 24361 14231 24395
rect 16773 24361 16807 24395
rect 17877 24361 17911 24395
rect 19073 24361 19107 24395
rect 21097 24361 21131 24395
rect 1869 24293 1903 24327
rect 1593 24225 1627 24259
rect 2881 24225 2915 24259
rect 4077 24225 4111 24259
rect 5181 24225 5215 24259
rect 5448 24225 5482 24259
rect 8033 24225 8067 24259
rect 10416 24225 10450 24259
rect 13001 24225 13035 24259
rect 16589 24225 16623 24259
rect 17693 24225 17727 24259
rect 18889 24225 18923 24259
rect 20913 24225 20947 24259
rect 8217 24157 8251 24191
rect 10149 24157 10183 24191
rect 13277 24157 13311 24191
rect 7573 24089 7607 24123
rect 12633 24089 12667 24123
rect 3065 24021 3099 24055
rect 4261 24021 4295 24055
rect 4905 24021 4939 24055
rect 6561 24021 6595 24055
rect 7113 24021 7147 24055
rect 11529 24021 11563 24055
rect 12449 24021 12483 24055
rect 13737 24021 13771 24055
rect 1593 23817 1627 23851
rect 2605 23817 2639 23851
rect 7297 23817 7331 23851
rect 7665 23817 7699 23851
rect 11897 23817 11931 23851
rect 15577 23817 15611 23851
rect 16681 23817 16715 23851
rect 18245 23817 18279 23851
rect 19349 23817 19383 23851
rect 20453 23817 20487 23851
rect 21557 23817 21591 23851
rect 9781 23749 9815 23783
rect 12725 23749 12759 23783
rect 2053 23681 2087 23715
rect 3709 23681 3743 23715
rect 10701 23681 10735 23715
rect 10793 23681 10827 23715
rect 12265 23681 12299 23715
rect 18981 23681 19015 23715
rect 1777 23613 1811 23647
rect 3801 23613 3835 23647
rect 4068 23613 4102 23647
rect 7757 23613 7791 23647
rect 10149 23613 10183 23647
rect 10609 23613 10643 23647
rect 12909 23613 12943 23647
rect 13176 23613 13210 23647
rect 15393 23613 15427 23647
rect 15945 23613 15979 23647
rect 16497 23613 16531 23647
rect 17049 23613 17083 23647
rect 18061 23613 18095 23647
rect 19165 23613 19199 23647
rect 19717 23613 19751 23647
rect 20269 23613 20303 23647
rect 20821 23613 20855 23647
rect 21373 23613 21407 23647
rect 21925 23613 21959 23647
rect 3249 23545 3283 23579
rect 5825 23545 5859 23579
rect 8024 23545 8058 23579
rect 16405 23545 16439 23579
rect 2881 23477 2915 23511
rect 5181 23477 5215 23511
rect 6101 23477 6135 23511
rect 6561 23477 6595 23511
rect 9137 23477 9171 23511
rect 10241 23477 10275 23511
rect 11345 23477 11379 23511
rect 14289 23477 14323 23511
rect 17693 23477 17727 23511
rect 18613 23477 18647 23511
rect 21189 23477 21223 23511
rect 7021 23273 7055 23307
rect 8493 23273 8527 23307
rect 14105 23273 14139 23307
rect 16681 23273 16715 23307
rect 19625 23273 19659 23307
rect 1869 23205 1903 23239
rect 4322 23205 4356 23239
rect 10324 23205 10358 23239
rect 12992 23205 13026 23239
rect 1593 23137 1627 23171
rect 2881 23137 2915 23171
rect 3801 23137 3835 23171
rect 4077 23137 4111 23171
rect 7113 23137 7147 23171
rect 7380 23137 7414 23171
rect 9965 23137 9999 23171
rect 10057 23137 10091 23171
rect 15568 23137 15602 23171
rect 19441 23137 19475 23171
rect 12725 23069 12759 23103
rect 15301 23069 15335 23103
rect 2421 22933 2455 22967
rect 3065 22933 3099 22967
rect 3433 22933 3467 22967
rect 5457 22933 5491 22967
rect 11437 22933 11471 22967
rect 12633 22933 12667 22967
rect 2789 22729 2823 22763
rect 4169 22729 4203 22763
rect 5181 22729 5215 22763
rect 9597 22729 9631 22763
rect 13001 22729 13035 22763
rect 2329 22661 2363 22695
rect 1777 22593 1811 22627
rect 3249 22593 3283 22627
rect 3341 22593 3375 22627
rect 5825 22593 5859 22627
rect 6929 22593 6963 22627
rect 7205 22593 7239 22627
rect 9229 22593 9263 22627
rect 10701 22593 10735 22627
rect 12449 22593 12483 22627
rect 1501 22525 1535 22559
rect 5089 22525 5123 22559
rect 5549 22525 5583 22559
rect 6653 22525 6687 22559
rect 7461 22525 7495 22559
rect 9965 22525 9999 22559
rect 10517 22525 10551 22559
rect 11161 22525 11195 22559
rect 12265 22525 12299 22559
rect 13737 22525 13771 22559
rect 16037 22525 16071 22559
rect 2697 22457 2731 22491
rect 3157 22457 3191 22491
rect 4721 22457 4755 22491
rect 5641 22457 5675 22491
rect 6929 22457 6963 22491
rect 10425 22457 10459 22491
rect 13982 22457 14016 22491
rect 6193 22389 6227 22423
rect 7113 22389 7147 22423
rect 8585 22389 8619 22423
rect 10057 22389 10091 22423
rect 13553 22389 13587 22423
rect 15117 22389 15151 22423
rect 15669 22389 15703 22423
rect 19441 22389 19475 22423
rect 2605 22185 2639 22219
rect 4077 22185 4111 22219
rect 10057 22185 10091 22219
rect 15301 22185 15335 22219
rect 16313 22185 16347 22219
rect 3801 22117 3835 22151
rect 8217 22117 8251 22151
rect 10508 22117 10542 22151
rect 1501 22049 1535 22083
rect 1777 22049 1811 22083
rect 2789 22049 2823 22083
rect 4445 22049 4479 22083
rect 4537 22049 4571 22083
rect 5273 22049 5307 22083
rect 6653 22049 6687 22083
rect 8309 22049 8343 22083
rect 10241 22049 10275 22083
rect 13185 22049 13219 22083
rect 13921 22049 13955 22083
rect 14289 22049 14323 22083
rect 4721 21981 4755 22015
rect 6745 21981 6779 22015
rect 6837 21981 6871 22015
rect 8401 21981 8435 22015
rect 8861 21981 8895 22015
rect 12725 21981 12759 22015
rect 13277 21981 13311 22015
rect 13461 21981 13495 22015
rect 2329 21913 2363 21947
rect 2973 21913 3007 21947
rect 7849 21913 7883 21947
rect 3433 21845 3467 21879
rect 5549 21845 5583 21879
rect 6009 21845 6043 21879
rect 6285 21845 6319 21879
rect 7573 21845 7607 21879
rect 11621 21845 11655 21879
rect 12817 21845 12851 21879
rect 2789 21641 2823 21675
rect 4261 21641 4295 21675
rect 4813 21641 4847 21675
rect 5273 21641 5307 21675
rect 8585 21641 8619 21675
rect 9505 21641 9539 21675
rect 10609 21641 10643 21675
rect 11897 21641 11931 21675
rect 13185 21641 13219 21675
rect 7481 21573 7515 21607
rect 8861 21573 8895 21607
rect 10885 21573 10919 21607
rect 12265 21573 12299 21607
rect 1685 21505 1719 21539
rect 2421 21505 2455 21539
rect 7389 21505 7423 21539
rect 7941 21505 7975 21539
rect 8125 21505 8159 21539
rect 9965 21505 9999 21539
rect 10149 21505 10183 21539
rect 11253 21505 11287 21539
rect 12725 21505 12759 21539
rect 13737 21505 13771 21539
rect 1501 21437 1535 21471
rect 2881 21437 2915 21471
rect 3148 21437 3182 21471
rect 5365 21437 5399 21471
rect 7849 21437 7883 21471
rect 11069 21437 11103 21471
rect 6009 21369 6043 21403
rect 9413 21369 9447 21403
rect 9873 21369 9907 21403
rect 13645 21369 13679 21403
rect 13982 21369 14016 21403
rect 5549 21301 5583 21335
rect 6285 21301 6319 21335
rect 15117 21301 15151 21335
rect 2421 21097 2455 21131
rect 3525 21097 3559 21131
rect 6377 21097 6411 21131
rect 8125 21097 8159 21131
rect 12909 21097 12943 21131
rect 13369 21097 13403 21131
rect 14289 21097 14323 21131
rect 15301 21097 15335 21131
rect 1869 21029 1903 21063
rect 5089 21029 5123 21063
rect 9965 21029 9999 21063
rect 10302 21029 10336 21063
rect 1593 20961 1627 20995
rect 2881 20961 2915 20995
rect 4997 20961 5031 20995
rect 6653 20961 6687 20995
rect 7012 20961 7046 20995
rect 12725 20961 12759 20995
rect 13277 20961 13311 20995
rect 5181 20893 5215 20927
rect 6009 20893 6043 20927
rect 6745 20893 6779 20927
rect 9505 20893 9539 20927
rect 10057 20893 10091 20927
rect 13461 20893 13495 20927
rect 2789 20825 2823 20859
rect 3801 20825 3835 20859
rect 4353 20825 4387 20859
rect 6469 20825 6503 20859
rect 12541 20825 12575 20859
rect 3065 20757 3099 20791
rect 4629 20757 4663 20791
rect 8769 20757 8803 20791
rect 11437 20757 11471 20791
rect 14013 20757 14047 20791
rect 3617 20553 3651 20587
rect 5089 20553 5123 20587
rect 6009 20553 6043 20587
rect 6653 20553 6687 20587
rect 8217 20553 8251 20587
rect 9045 20553 9079 20587
rect 10609 20553 10643 20587
rect 11897 20553 11931 20587
rect 13277 20553 13311 20587
rect 15209 20553 15243 20587
rect 5733 20485 5767 20519
rect 2329 20417 2363 20451
rect 10241 20417 10275 20451
rect 11069 20417 11103 20451
rect 13829 20417 13863 20451
rect 1501 20349 1535 20383
rect 1777 20349 1811 20383
rect 3709 20349 3743 20383
rect 6837 20349 6871 20383
rect 9505 20349 9539 20383
rect 10057 20349 10091 20383
rect 12265 20349 12299 20383
rect 12449 20349 12483 20383
rect 3976 20281 4010 20315
rect 7104 20281 7138 20315
rect 9965 20281 9999 20315
rect 12725 20281 12759 20315
rect 14096 20281 14130 20315
rect 2697 20213 2731 20247
rect 3065 20213 3099 20247
rect 9597 20213 9631 20247
rect 11345 20213 11379 20247
rect 13553 20213 13587 20247
rect 16313 20213 16347 20247
rect 6929 20009 6963 20043
rect 8493 20009 8527 20043
rect 13001 20009 13035 20043
rect 13185 20009 13219 20043
rect 15761 20009 15795 20043
rect 1777 19941 1811 19975
rect 4629 19941 4663 19975
rect 4988 19941 5022 19975
rect 9045 19941 9079 19975
rect 9965 19941 9999 19975
rect 10302 19941 10336 19975
rect 13645 19941 13679 19975
rect 14197 19941 14231 19975
rect 15669 19941 15703 19975
rect 1501 19873 1535 19907
rect 2789 19873 2823 19907
rect 4721 19873 4755 19907
rect 7573 19873 7607 19907
rect 8401 19873 8435 19907
rect 9505 19873 9539 19907
rect 10057 19873 10091 19907
rect 13553 19873 13587 19907
rect 2329 19805 2363 19839
rect 7849 19805 7883 19839
rect 8677 19805 8711 19839
rect 13829 19805 13863 19839
rect 15853 19805 15887 19839
rect 8033 19737 8067 19771
rect 12633 19737 12667 19771
rect 2605 19669 2639 19703
rect 2973 19669 3007 19703
rect 3433 19669 3467 19703
rect 3801 19669 3835 19703
rect 6101 19669 6135 19703
rect 7297 19669 7331 19703
rect 7389 19669 7423 19703
rect 11437 19669 11471 19703
rect 15301 19669 15335 19703
rect 4077 19465 4111 19499
rect 5181 19465 5215 19499
rect 5457 19465 5491 19499
rect 9321 19465 9355 19499
rect 10057 19465 10091 19499
rect 10793 19465 10827 19499
rect 12817 19465 12851 19499
rect 13185 19465 13219 19499
rect 14657 19465 14691 19499
rect 15393 19465 15427 19499
rect 16313 19465 16347 19499
rect 2605 19329 2639 19363
rect 3985 19329 4019 19363
rect 4721 19329 4755 19363
rect 7941 19329 7975 19363
rect 3249 19261 3283 19295
rect 4537 19261 4571 19295
rect 5641 19261 5675 19295
rect 7481 19261 7515 19295
rect 8208 19261 8242 19295
rect 10977 19261 11011 19295
rect 11069 19261 11103 19295
rect 11897 19261 11931 19295
rect 13277 19261 13311 19295
rect 15761 19261 15795 19295
rect 16681 19261 16715 19295
rect 1961 19193 1995 19227
rect 2421 19193 2455 19227
rect 6285 19193 6319 19227
rect 11345 19193 11379 19227
rect 12265 19193 12299 19227
rect 13522 19193 13556 19227
rect 2053 19125 2087 19159
rect 2513 19125 2547 19159
rect 3617 19125 3651 19159
rect 4445 19125 4479 19159
rect 5825 19125 5859 19159
rect 6653 19125 6687 19159
rect 6837 19125 6871 19159
rect 7849 19125 7883 19159
rect 10609 19125 10643 19159
rect 15945 19125 15979 19159
rect 1409 18921 1443 18955
rect 4445 18921 4479 18955
rect 5549 18921 5583 18955
rect 6101 18921 6135 18955
rect 8769 18921 8803 18955
rect 13921 18921 13955 18955
rect 16037 18921 16071 18955
rect 5089 18853 5123 18887
rect 6193 18853 6227 18887
rect 8401 18853 8435 18887
rect 12786 18853 12820 18887
rect 15577 18853 15611 18887
rect 2789 18785 2823 18819
rect 3433 18785 3467 18819
rect 4537 18785 4571 18819
rect 7665 18785 7699 18819
rect 7757 18785 7791 18819
rect 9689 18785 9723 18819
rect 11345 18785 11379 18819
rect 15301 18785 15335 18819
rect 2881 18717 2915 18751
rect 2973 18717 3007 18751
rect 4629 18717 4663 18751
rect 6377 18717 6411 18751
rect 7849 18717 7883 18751
rect 9873 18717 9907 18751
rect 11437 18717 11471 18751
rect 11621 18717 11655 18751
rect 12541 18717 12575 18751
rect 2421 18649 2455 18683
rect 3801 18649 3835 18683
rect 4077 18649 4111 18683
rect 5733 18649 5767 18683
rect 7297 18649 7331 18683
rect 10517 18649 10551 18683
rect 10977 18649 11011 18683
rect 2145 18581 2179 18615
rect 6929 18581 6963 18615
rect 9321 18581 9355 18615
rect 10885 18581 10919 18615
rect 12081 18581 12115 18615
rect 12449 18581 12483 18615
rect 6193 18377 6227 18411
rect 10701 18377 10735 18411
rect 10793 18377 10827 18411
rect 11897 18377 11931 18411
rect 15301 18377 15335 18411
rect 16129 18377 16163 18411
rect 5641 18309 5675 18343
rect 10333 18309 10367 18343
rect 1685 18241 1719 18275
rect 7481 18241 7515 18275
rect 8217 18241 8251 18275
rect 9689 18241 9723 18275
rect 9873 18241 9907 18275
rect 11437 18241 11471 18275
rect 15669 18241 15703 18275
rect 1777 18173 1811 18207
rect 2044 18173 2078 18207
rect 4261 18173 4295 18207
rect 7297 18173 7331 18207
rect 9137 18173 9171 18207
rect 11161 18173 11195 18207
rect 12449 18173 12483 18207
rect 15393 18173 15427 18207
rect 3801 18105 3835 18139
rect 4169 18105 4203 18139
rect 4528 18105 4562 18139
rect 6561 18105 6595 18139
rect 7205 18105 7239 18139
rect 8769 18105 8803 18139
rect 9597 18105 9631 18139
rect 12265 18105 12299 18139
rect 12694 18105 12728 18139
rect 3157 18037 3191 18071
rect 6837 18037 6871 18071
rect 7941 18037 7975 18071
rect 9229 18037 9263 18071
rect 11253 18037 11287 18071
rect 13829 18037 13863 18071
rect 14381 18037 14415 18071
rect 3801 17833 3835 17867
rect 4077 17833 4111 17867
rect 5089 17833 5123 17867
rect 5641 17833 5675 17867
rect 11621 17833 11655 17867
rect 13553 17833 13587 17867
rect 14381 17833 14415 17867
rect 4445 17765 4479 17799
rect 1501 17697 1535 17731
rect 1768 17697 1802 17731
rect 5825 17697 5859 17731
rect 6276 17697 6310 17731
rect 9505 17697 9539 17731
rect 9956 17697 9990 17731
rect 12440 17697 12474 17731
rect 4537 17629 4571 17663
rect 4721 17629 4755 17663
rect 5549 17629 5583 17663
rect 6009 17629 6043 17663
rect 7941 17629 7975 17663
rect 8585 17629 8619 17663
rect 9689 17629 9723 17663
rect 12173 17629 12207 17663
rect 2881 17561 2915 17595
rect 3433 17561 3467 17595
rect 11069 17561 11103 17595
rect 7389 17493 7423 17527
rect 8309 17493 8343 17527
rect 9045 17493 9079 17527
rect 11989 17493 12023 17527
rect 2881 17289 2915 17323
rect 4169 17289 4203 17323
rect 4445 17289 4479 17323
rect 5181 17289 5215 17323
rect 6285 17289 6319 17323
rect 9413 17289 9447 17323
rect 11069 17289 11103 17323
rect 13553 17289 13587 17323
rect 11897 17221 11931 17255
rect 12449 17221 12483 17255
rect 2053 17153 2087 17187
rect 2421 17153 2455 17187
rect 3525 17153 3559 17187
rect 5641 17153 5675 17187
rect 5825 17153 5859 17187
rect 6561 17153 6595 17187
rect 6837 17153 6871 17187
rect 9321 17153 9355 17187
rect 9873 17153 9907 17187
rect 10057 17153 10091 17187
rect 11345 17153 11379 17187
rect 12265 17153 12299 17187
rect 1409 17085 1443 17119
rect 5549 17085 5583 17119
rect 8769 17085 8803 17119
rect 13001 17153 13035 17187
rect 13185 17153 13219 17187
rect 14381 17153 14415 17187
rect 2789 17017 2823 17051
rect 7104 17017 7138 17051
rect 12449 17017 12483 17051
rect 14626 17017 14660 17051
rect 1593 16949 1627 16983
rect 3249 16949 3283 16983
rect 3341 16949 3375 16983
rect 4905 16949 4939 16983
rect 8217 16949 8251 16983
rect 9781 16949 9815 16983
rect 10517 16949 10551 16983
rect 12541 16949 12575 16983
rect 12909 16949 12943 16983
rect 14197 16949 14231 16983
rect 15761 16949 15795 16983
rect 1869 16745 1903 16779
rect 3341 16745 3375 16779
rect 4077 16745 4111 16779
rect 4629 16745 4663 16779
rect 5089 16745 5123 16779
rect 6101 16745 6135 16779
rect 6653 16745 6687 16779
rect 7021 16745 7055 16779
rect 8033 16745 8067 16779
rect 9413 16745 9447 16779
rect 10149 16745 10183 16779
rect 12081 16745 12115 16779
rect 14105 16745 14139 16779
rect 2237 16677 2271 16711
rect 3617 16677 3651 16711
rect 7113 16677 7147 16711
rect 10609 16677 10643 16711
rect 13185 16677 13219 16711
rect 14013 16677 14047 16711
rect 2329 16609 2363 16643
rect 2881 16609 2915 16643
rect 5457 16609 5491 16643
rect 6561 16609 6595 16643
rect 8309 16609 8343 16643
rect 9873 16609 9907 16643
rect 10517 16609 10551 16643
rect 11161 16609 11195 16643
rect 11621 16609 11655 16643
rect 11897 16609 11931 16643
rect 12449 16609 12483 16643
rect 2513 16541 2547 16575
rect 5549 16541 5583 16575
rect 5641 16541 5675 16575
rect 7297 16541 7331 16575
rect 8493 16541 8527 16575
rect 10701 16541 10735 16575
rect 12541 16541 12575 16575
rect 12633 16541 12667 16575
rect 14197 16541 14231 16575
rect 13645 16473 13679 16507
rect 1685 16405 1719 16439
rect 4997 16405 5031 16439
rect 7757 16405 7791 16439
rect 9137 16405 9171 16439
rect 11713 16405 11747 16439
rect 2973 16201 3007 16235
rect 6285 16201 6319 16235
rect 7849 16201 7883 16235
rect 10609 16201 10643 16235
rect 13001 16201 13035 16235
rect 15301 16201 15335 16235
rect 13737 16133 13771 16167
rect 2053 16065 2087 16099
rect 5549 16065 5583 16099
rect 7389 16065 7423 16099
rect 9413 16065 9447 16099
rect 11253 16065 11287 16099
rect 13369 16065 13403 16099
rect 16681 16065 16715 16099
rect 1961 15997 1995 16031
rect 3065 15997 3099 16031
rect 3321 15997 3355 16031
rect 7205 15997 7239 16031
rect 8769 15997 8803 16031
rect 10977 15997 11011 16031
rect 11069 15997 11103 16031
rect 13921 15997 13955 16031
rect 16405 15997 16439 16031
rect 17141 15997 17175 16031
rect 7297 15929 7331 15963
rect 9321 15929 9355 15963
rect 14188 15929 14222 15963
rect 1501 15861 1535 15895
rect 1869 15861 1903 15895
rect 2605 15861 2639 15895
rect 4445 15861 4479 15895
rect 5089 15861 5123 15895
rect 6561 15861 6595 15895
rect 6837 15861 6871 15895
rect 8309 15861 8343 15895
rect 8861 15861 8895 15895
rect 9229 15861 9263 15895
rect 10149 15861 10183 15895
rect 12173 15861 12207 15895
rect 2053 15657 2087 15691
rect 3157 15657 3191 15691
rect 3525 15657 3559 15691
rect 4261 15657 4295 15691
rect 5181 15657 5215 15691
rect 6653 15657 6687 15691
rect 7297 15657 7331 15691
rect 8585 15657 8619 15691
rect 8953 15657 8987 15691
rect 10149 15657 10183 15691
rect 10793 15657 10827 15691
rect 11345 15657 11379 15691
rect 12725 15657 12759 15691
rect 13369 15657 13403 15691
rect 14657 15657 14691 15691
rect 3801 15589 3835 15623
rect 12449 15589 12483 15623
rect 15577 15589 15611 15623
rect 2421 15521 2455 15555
rect 4077 15521 4111 15555
rect 5540 15521 5574 15555
rect 7757 15521 7791 15555
rect 10057 15521 10091 15555
rect 11713 15521 11747 15555
rect 13277 15521 13311 15555
rect 15301 15521 15335 15555
rect 2513 15453 2547 15487
rect 2697 15453 2731 15487
rect 4721 15453 4755 15487
rect 5273 15453 5307 15487
rect 7941 15453 7975 15487
rect 10241 15453 10275 15487
rect 11805 15453 11839 15487
rect 11897 15453 11931 15487
rect 13461 15453 13495 15487
rect 14013 15385 14047 15419
rect 1961 15317 1995 15351
rect 7665 15317 7699 15351
rect 9229 15317 9263 15351
rect 9689 15317 9723 15351
rect 11161 15317 11195 15351
rect 12909 15317 12943 15351
rect 14289 15317 14323 15351
rect 5641 15113 5675 15147
rect 6285 15113 6319 15147
rect 7113 15113 7147 15147
rect 7573 15113 7607 15147
rect 9045 15113 9079 15147
rect 10517 15113 10551 15147
rect 11069 15113 11103 15147
rect 11529 15113 11563 15147
rect 13093 15113 13127 15147
rect 14933 15113 14967 15147
rect 15485 15113 15519 15147
rect 21833 15113 21867 15147
rect 7389 14977 7423 15011
rect 8033 14977 8067 15011
rect 8217 14977 8251 15011
rect 1501 14909 1535 14943
rect 4261 14909 4295 14943
rect 9137 14909 9171 14943
rect 13553 14909 13587 14943
rect 13820 14909 13854 14943
rect 21649 14909 21683 14943
rect 22201 14909 22235 14943
rect 1768 14841 1802 14875
rect 4169 14841 4203 14875
rect 4528 14841 4562 14875
rect 6653 14841 6687 14875
rect 8585 14841 8619 14875
rect 9404 14841 9438 14875
rect 11897 14841 11931 14875
rect 2881 14773 2915 14807
rect 3433 14773 3467 14807
rect 7941 14773 7975 14807
rect 12173 14773 12207 14807
rect 12541 14773 12575 14807
rect 13369 14773 13403 14807
rect 1409 14569 1443 14603
rect 3525 14569 3559 14603
rect 4629 14569 4663 14603
rect 8033 14569 8067 14603
rect 8493 14569 8527 14603
rect 9965 14569 9999 14603
rect 12173 14569 12207 14603
rect 12633 14569 12667 14603
rect 14105 14569 14139 14603
rect 14657 14569 14691 14603
rect 8401 14501 8435 14535
rect 10508 14501 10542 14535
rect 1777 14433 1811 14467
rect 2973 14433 3007 14467
rect 4077 14433 4111 14467
rect 5181 14433 5215 14467
rect 5448 14433 5482 14467
rect 10241 14433 10275 14467
rect 12725 14433 12759 14467
rect 12992 14433 13026 14467
rect 1869 14365 1903 14399
rect 2053 14365 2087 14399
rect 8585 14365 8619 14399
rect 2421 14297 2455 14331
rect 4261 14297 4295 14331
rect 6561 14297 6595 14331
rect 2789 14229 2823 14263
rect 3801 14229 3835 14263
rect 4997 14229 5031 14263
rect 7205 14229 7239 14263
rect 7573 14229 7607 14263
rect 9229 14229 9263 14263
rect 11621 14229 11655 14263
rect 3617 14025 3651 14059
rect 3985 14025 4019 14059
rect 6837 14025 6871 14059
rect 7941 14025 7975 14059
rect 9689 14025 9723 14059
rect 10517 14025 10551 14059
rect 11345 14025 11379 14059
rect 12173 14025 12207 14059
rect 13829 14025 13863 14059
rect 5181 13957 5215 13991
rect 11897 13957 11931 13991
rect 5089 13889 5123 13923
rect 5641 13889 5675 13923
rect 5825 13889 5859 13923
rect 7297 13889 7331 13923
rect 7389 13889 7423 13923
rect 16405 13889 16439 13923
rect 21005 13889 21039 13923
rect 1685 13821 1719 13855
rect 1952 13821 1986 13855
rect 4721 13821 4755 13855
rect 8309 13821 8343 13855
rect 8401 13821 8435 13855
rect 12449 13821 12483 13855
rect 12705 13821 12739 13855
rect 16129 13821 16163 13855
rect 16865 13821 16899 13855
rect 20729 13821 20763 13855
rect 21465 13821 21499 13855
rect 4169 13753 4203 13787
rect 5549 13753 5583 13787
rect 10885 13753 10919 13787
rect 3065 13685 3099 13719
rect 6193 13685 6227 13719
rect 6561 13685 6595 13719
rect 7205 13685 7239 13719
rect 2789 13481 2823 13515
rect 3065 13481 3099 13515
rect 3433 13481 3467 13515
rect 5733 13481 5767 13515
rect 7941 13481 7975 13515
rect 10149 13481 10183 13515
rect 12449 13481 12483 13515
rect 12909 13481 12943 13515
rect 5641 13413 5675 13447
rect 6929 13413 6963 13447
rect 7573 13413 7607 13447
rect 9505 13413 9539 13447
rect 13461 13413 13495 13447
rect 17693 13413 17727 13447
rect 2053 13345 2087 13379
rect 3617 13345 3651 13379
rect 8401 13345 8435 13379
rect 10057 13345 10091 13379
rect 12817 13345 12851 13379
rect 17417 13345 17451 13379
rect 2145 13277 2179 13311
rect 2329 13277 2363 13311
rect 4077 13277 4111 13311
rect 4813 13277 4847 13311
rect 5917 13277 5951 13311
rect 7021 13277 7055 13311
rect 8493 13277 8527 13311
rect 8677 13277 8711 13311
rect 10241 13277 10275 13311
rect 13093 13277 13127 13311
rect 5273 13209 5307 13243
rect 6469 13209 6503 13243
rect 8033 13209 8067 13243
rect 9689 13209 9723 13243
rect 11069 13209 11103 13243
rect 11897 13209 11931 13243
rect 1685 13141 1719 13175
rect 9137 13141 9171 13175
rect 10793 13141 10827 13175
rect 11437 13141 11471 13175
rect 1685 12937 1719 12971
rect 2145 12937 2179 12971
rect 4813 12937 4847 12971
rect 5917 12937 5951 12971
rect 7941 12937 7975 12971
rect 9781 12937 9815 12971
rect 11437 12937 11471 12971
rect 11897 12937 11931 12971
rect 12449 12937 12483 12971
rect 13829 12937 13863 12971
rect 15485 12937 15519 12971
rect 4721 12869 4755 12903
rect 6561 12869 6595 12903
rect 10425 12869 10459 12903
rect 13553 12869 13587 12903
rect 17785 12869 17819 12903
rect 2329 12801 2363 12835
rect 5273 12801 5307 12835
rect 5365 12801 5399 12835
rect 8401 12801 8435 12835
rect 10885 12801 10919 12835
rect 10977 12801 11011 12835
rect 12909 12801 12943 12835
rect 13001 12801 13035 12835
rect 14289 12801 14323 12835
rect 16957 12801 16991 12835
rect 18337 12801 18371 12835
rect 2585 12733 2619 12767
rect 5181 12733 5215 12767
rect 8309 12733 8343 12767
rect 12173 12733 12207 12767
rect 12817 12733 12851 12767
rect 14013 12733 14047 12767
rect 14749 12733 14783 12767
rect 15301 12733 15335 12767
rect 15853 12733 15887 12767
rect 16681 12733 16715 12767
rect 17417 12733 17451 12767
rect 18061 12733 18095 12767
rect 18797 12733 18831 12767
rect 4353 12665 4387 12699
rect 6193 12665 6227 12699
rect 7665 12665 7699 12699
rect 8668 12665 8702 12699
rect 3709 12597 3743 12631
rect 6837 12597 6871 12631
rect 8125 12597 8159 12631
rect 10793 12597 10827 12631
rect 1685 12393 1719 12427
rect 2789 12393 2823 12427
rect 7021 12393 7055 12427
rect 7481 12393 7515 12427
rect 9229 12393 9263 12427
rect 9781 12393 9815 12427
rect 10701 12393 10735 12427
rect 12725 12393 12759 12427
rect 13093 12393 13127 12427
rect 13277 12393 13311 12427
rect 6561 12325 6595 12359
rect 11038 12325 11072 12359
rect 2145 12257 2179 12291
rect 3525 12257 3559 12291
rect 4077 12257 4111 12291
rect 4344 12257 4378 12291
rect 7389 12257 7423 12291
rect 8116 12257 8150 12291
rect 13645 12257 13679 12291
rect 2237 12189 2271 12223
rect 2421 12189 2455 12223
rect 7573 12189 7607 12223
rect 7849 12189 7883 12223
rect 10793 12189 10827 12223
rect 13737 12189 13771 12223
rect 13829 12189 13863 12223
rect 1777 12121 1811 12155
rect 3157 12053 3191 12087
rect 5457 12053 5491 12087
rect 6009 12053 6043 12087
rect 6929 12053 6963 12087
rect 10241 12053 10275 12087
rect 12173 12053 12207 12087
rect 2697 11849 2731 11883
rect 3525 11849 3559 11883
rect 5365 11849 5399 11883
rect 6285 11849 6319 11883
rect 10701 11849 10735 11883
rect 11253 11849 11287 11883
rect 11897 11849 11931 11883
rect 12173 11849 12207 11883
rect 14381 11849 14415 11883
rect 8217 11781 8251 11815
rect 2237 11713 2271 11747
rect 6837 11713 6871 11747
rect 9229 11713 9263 11747
rect 14933 11713 14967 11747
rect 2053 11645 2087 11679
rect 3893 11645 3927 11679
rect 3985 11645 4019 11679
rect 4241 11645 4275 11679
rect 7093 11645 7127 11679
rect 9321 11645 9355 11679
rect 9588 11645 9622 11679
rect 12449 11645 12483 11679
rect 12705 11645 12739 11679
rect 1685 11509 1719 11543
rect 2145 11509 2179 11543
rect 3065 11509 3099 11543
rect 3709 11509 3743 11543
rect 6561 11509 6595 11543
rect 8861 11509 8895 11543
rect 13829 11509 13863 11543
rect 14749 11509 14783 11543
rect 1777 11305 1811 11339
rect 3157 11305 3191 11339
rect 4721 11305 4755 11339
rect 6377 11305 6411 11339
rect 7113 11305 7147 11339
rect 8493 11305 8527 11339
rect 8953 11305 8987 11339
rect 11253 11305 11287 11339
rect 11621 11305 11655 11339
rect 11989 11305 12023 11339
rect 12541 11305 12575 11339
rect 14105 11305 14139 11339
rect 3525 11237 3559 11271
rect 5264 11237 5298 11271
rect 12992 11237 13026 11271
rect 2145 11169 2179 11203
rect 4353 11169 4387 11203
rect 4997 11169 5031 11203
rect 7849 11169 7883 11203
rect 9229 11169 9263 11203
rect 10609 11169 10643 11203
rect 12725 11169 12759 11203
rect 18521 11169 18555 11203
rect 18797 11169 18831 11203
rect 2237 11101 2271 11135
rect 2421 11101 2455 11135
rect 7941 11101 7975 11135
rect 8125 11101 8159 11135
rect 10701 11101 10735 11135
rect 10793 11101 10827 11135
rect 2789 11033 2823 11067
rect 7481 11033 7515 11067
rect 9045 11033 9079 11067
rect 10241 11033 10275 11067
rect 1685 10965 1719 10999
rect 10149 10965 10183 10999
rect 3249 10761 3283 10795
rect 4169 10761 4203 10795
rect 5457 10761 5491 10795
rect 5733 10761 5767 10795
rect 6101 10761 6135 10795
rect 9045 10761 9079 10795
rect 9689 10761 9723 10795
rect 10149 10761 10183 10795
rect 12449 10761 12483 10795
rect 13553 10761 13587 10795
rect 18521 10761 18555 10795
rect 3893 10625 3927 10659
rect 4997 10625 5031 10659
rect 7665 10625 7699 10659
rect 10609 10625 10643 10659
rect 10793 10625 10827 10659
rect 13001 10625 13035 10659
rect 20453 10625 20487 10659
rect 1869 10557 1903 10591
rect 4721 10557 4755 10591
rect 20177 10557 20211 10591
rect 20913 10557 20947 10591
rect 2136 10489 2170 10523
rect 4813 10489 4847 10523
rect 6653 10489 6687 10523
rect 7573 10489 7607 10523
rect 7932 10489 7966 10523
rect 10517 10489 10551 10523
rect 12173 10489 12207 10523
rect 12817 10489 12851 10523
rect 1777 10421 1811 10455
rect 4353 10421 4387 10455
rect 7205 10421 7239 10455
rect 9965 10421 9999 10455
rect 11161 10421 11195 10455
rect 11529 10421 11563 10455
rect 12909 10421 12943 10455
rect 1869 10217 1903 10251
rect 2237 10217 2271 10251
rect 2605 10217 2639 10251
rect 5457 10217 5491 10251
rect 5641 10217 5675 10251
rect 6009 10217 6043 10251
rect 7297 10217 7331 10251
rect 7757 10217 7791 10251
rect 9045 10217 9079 10251
rect 10057 10217 10091 10251
rect 12541 10217 12575 10251
rect 12817 10217 12851 10251
rect 13185 10217 13219 10251
rect 6101 10149 6135 10183
rect 10416 10149 10450 10183
rect 2697 10081 2731 10115
rect 4445 10081 4479 10115
rect 7665 10081 7699 10115
rect 18889 10081 18923 10115
rect 19165 10081 19199 10115
rect 2789 10013 2823 10047
rect 3249 10013 3283 10047
rect 4537 10013 4571 10047
rect 4721 10013 4755 10047
rect 6285 10013 6319 10047
rect 7205 10013 7239 10047
rect 7849 10013 7883 10047
rect 8309 10013 8343 10047
rect 10149 10013 10183 10047
rect 4077 9945 4111 9979
rect 5089 9945 5123 9979
rect 3893 9877 3927 9911
rect 6837 9877 6871 9911
rect 8677 9877 8711 9911
rect 9413 9877 9447 9911
rect 11529 9877 11563 9911
rect 6009 9673 6043 9707
rect 10241 9673 10275 9707
rect 18889 9673 18923 9707
rect 3985 9605 4019 9639
rect 6653 9605 6687 9639
rect 9689 9605 9723 9639
rect 10425 9537 10459 9571
rect 19625 9537 19659 9571
rect 1593 9469 1627 9503
rect 4077 9469 4111 9503
rect 7665 9469 7699 9503
rect 7932 9469 7966 9503
rect 19349 9469 19383 9503
rect 20085 9469 20119 9503
rect 1860 9401 1894 9435
rect 3525 9401 3559 9435
rect 4344 9401 4378 9435
rect 7389 9401 7423 9435
rect 2973 9333 3007 9367
rect 5457 9333 5491 9367
rect 9045 9333 9079 9367
rect 10885 9333 10919 9367
rect 2697 9129 2731 9163
rect 2973 9129 3007 9163
rect 3433 9129 3467 9163
rect 6377 9129 6411 9163
rect 8309 9129 8343 9163
rect 11897 9129 11931 9163
rect 1961 9061 1995 9095
rect 4353 9061 4387 9095
rect 4712 9061 4746 9095
rect 3617 8993 3651 9027
rect 4445 8993 4479 9027
rect 7196 8993 7230 9027
rect 10517 8993 10551 9027
rect 10773 8993 10807 9027
rect 2053 8925 2087 8959
rect 2237 8925 2271 8959
rect 6929 8925 6963 8959
rect 1593 8789 1627 8823
rect 5825 8789 5859 8823
rect 6745 8789 6779 8823
rect 1593 8585 1627 8619
rect 2697 8585 2731 8619
rect 2973 8585 3007 8619
rect 3157 8585 3191 8619
rect 4537 8585 4571 8619
rect 4905 8585 4939 8619
rect 5089 8585 5123 8619
rect 8309 8585 8343 8619
rect 10609 8585 10643 8619
rect 6837 8517 6871 8551
rect 8401 8517 8435 8551
rect 10885 8517 10919 8551
rect 2053 8449 2087 8483
rect 2145 8449 2179 8483
rect 3617 8449 3651 8483
rect 3801 8449 3835 8483
rect 5641 8449 5675 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 8861 8449 8895 8483
rect 8953 8449 8987 8483
rect 3525 8381 3559 8415
rect 5457 8381 5491 8415
rect 6285 8381 6319 8415
rect 5549 8313 5583 8347
rect 6653 8313 6687 8347
rect 7205 8313 7239 8347
rect 8769 8313 8803 8347
rect 1961 8245 1995 8279
rect 7941 8245 7975 8279
rect 1593 8041 1627 8075
rect 2421 8041 2455 8075
rect 2789 8041 2823 8075
rect 3157 8041 3191 8075
rect 3617 8041 3651 8075
rect 4169 8041 4203 8075
rect 4629 8041 4663 8075
rect 5089 8041 5123 8075
rect 5549 8041 5583 8075
rect 7021 8041 7055 8075
rect 7573 8041 7607 8075
rect 8125 8041 8159 8075
rect 8677 8041 8711 8075
rect 2053 7973 2087 8007
rect 5886 7973 5920 8007
rect 5641 7837 5675 7871
rect 2053 7497 2087 7531
rect 2421 7497 2455 7531
rect 3525 7497 3559 7531
rect 4537 7497 4571 7531
rect 6009 7497 6043 7531
rect 7297 7497 7331 7531
rect 8125 7497 8159 7531
rect 8585 7497 8619 7531
rect 22477 7497 22511 7531
rect 5733 7361 5767 7395
rect 6837 7361 6871 7395
rect 8309 7293 8343 7327
rect 22293 7293 22327 7327
rect 22845 7293 22879 7327
rect 1685 7157 1719 7191
rect 22753 6817 22787 6851
rect 22937 6681 22971 6715
rect 22753 6409 22787 6443
rect 23857 6409 23891 6443
rect 23673 6205 23707 6239
rect 24225 6205 24259 6239
rect 24225 5865 24259 5899
rect 24041 5729 24075 5763
rect 24041 5321 24075 5355
rect 24777 5321 24811 5355
rect 24593 5117 24627 5151
rect 25145 5117 25179 5151
rect 24777 4777 24811 4811
rect 24593 4641 24627 4675
rect 24593 4165 24627 4199
rect 2329 3009 2363 3043
rect 2237 2873 2271 2907
rect 2596 2873 2630 2907
rect 3709 2805 3743 2839
rect 2329 2601 2363 2635
<< metal1 >>
rect 3418 27344 3424 27396
rect 3476 27384 3482 27396
rect 7190 27384 7196 27396
rect 3476 27356 7196 27384
rect 3476 27344 3482 27356
rect 7190 27344 7196 27356
rect 7248 27344 7254 27396
rect 3510 26324 3516 26376
rect 3568 26364 3574 26376
rect 9214 26364 9220 26376
rect 3568 26336 9220 26364
rect 3568 26324 3574 26336
rect 9214 26324 9220 26336
rect 9272 26324 9278 26376
rect 3418 26256 3424 26308
rect 3476 26296 3482 26308
rect 8110 26296 8116 26308
rect 3476 26268 8116 26296
rect 3476 26256 3482 26268
rect 8110 26256 8116 26268
rect 8168 26256 8174 26308
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 4890 25440 4896 25492
rect 4948 25480 4954 25492
rect 5261 25483 5319 25489
rect 5261 25480 5273 25483
rect 4948 25452 5273 25480
rect 4948 25440 4954 25452
rect 5261 25449 5273 25452
rect 5307 25480 5319 25483
rect 7650 25480 7656 25492
rect 5307 25452 7656 25480
rect 5307 25449 5319 25452
rect 5261 25443 5319 25449
rect 7650 25440 7656 25452
rect 7708 25440 7714 25492
rect 8110 25440 8116 25492
rect 8168 25480 8174 25492
rect 8205 25483 8263 25489
rect 8205 25480 8217 25483
rect 8168 25452 8217 25480
rect 8168 25440 8174 25452
rect 8205 25449 8217 25452
rect 8251 25449 8263 25483
rect 8205 25443 8263 25449
rect 1946 25372 1952 25424
rect 2004 25412 2010 25424
rect 2004 25384 5488 25412
rect 2004 25372 2010 25384
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 2038 25344 2044 25356
rect 1443 25316 2044 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 2038 25304 2044 25316
rect 2096 25304 2102 25356
rect 2314 25304 2320 25356
rect 2372 25344 2378 25356
rect 2501 25347 2559 25353
rect 2501 25344 2513 25347
rect 2372 25316 2513 25344
rect 2372 25304 2378 25316
rect 2501 25313 2513 25316
rect 2547 25313 2559 25347
rect 2501 25307 2559 25313
rect 4614 25304 4620 25356
rect 4672 25344 4678 25356
rect 5166 25344 5172 25356
rect 4672 25316 5172 25344
rect 4672 25304 4678 25316
rect 5166 25304 5172 25316
rect 5224 25304 5230 25356
rect 5074 25236 5080 25288
rect 5132 25276 5138 25288
rect 5353 25279 5411 25285
rect 5353 25276 5365 25279
rect 5132 25248 5365 25276
rect 5132 25236 5138 25248
rect 5353 25245 5365 25248
rect 5399 25245 5411 25279
rect 5460 25276 5488 25384
rect 6270 25372 6276 25424
rect 6328 25412 6334 25424
rect 12621 25415 12679 25421
rect 12621 25412 12633 25415
rect 6328 25384 12633 25412
rect 6328 25372 6334 25384
rect 12621 25381 12633 25384
rect 12667 25381 12679 25415
rect 12621 25375 12679 25381
rect 6917 25347 6975 25353
rect 6917 25313 6929 25347
rect 6963 25344 6975 25347
rect 7098 25344 7104 25356
rect 6963 25316 7104 25344
rect 6963 25313 6975 25316
rect 6917 25307 6975 25313
rect 7098 25304 7104 25316
rect 7156 25304 7162 25356
rect 8021 25347 8079 25353
rect 8021 25313 8033 25347
rect 8067 25344 8079 25347
rect 8573 25347 8631 25353
rect 8573 25344 8585 25347
rect 8067 25316 8585 25344
rect 8067 25313 8079 25316
rect 8021 25307 8079 25313
rect 8573 25313 8585 25316
rect 8619 25313 8631 25347
rect 9766 25344 9772 25356
rect 9727 25316 9772 25344
rect 8573 25307 8631 25313
rect 8036 25276 8064 25307
rect 9766 25304 9772 25316
rect 9824 25304 9830 25356
rect 10870 25276 10876 25288
rect 5460 25248 8064 25276
rect 10831 25248 10876 25276
rect 5353 25239 5411 25245
rect 10870 25236 10876 25248
rect 10928 25236 10934 25288
rect 1581 25211 1639 25217
rect 1581 25177 1593 25211
rect 1627 25208 1639 25211
rect 2774 25208 2780 25220
rect 1627 25180 2780 25208
rect 1627 25177 1639 25180
rect 1581 25171 1639 25177
rect 2774 25168 2780 25180
rect 2832 25168 2838 25220
rect 3510 25168 3516 25220
rect 3568 25208 3574 25220
rect 7101 25211 7159 25217
rect 7101 25208 7113 25211
rect 3568 25180 7113 25208
rect 3568 25168 3574 25180
rect 7101 25177 7113 25180
rect 7147 25177 7159 25211
rect 7101 25171 7159 25177
rect 7190 25168 7196 25220
rect 7248 25208 7254 25220
rect 9953 25211 10011 25217
rect 9953 25208 9965 25211
rect 7248 25180 9965 25208
rect 7248 25168 7254 25180
rect 9953 25177 9965 25180
rect 9999 25177 10011 25211
rect 9953 25171 10011 25177
rect 2685 25143 2743 25149
rect 2685 25109 2697 25143
rect 2731 25140 2743 25143
rect 2866 25140 2872 25152
rect 2731 25112 2872 25140
rect 2731 25109 2743 25112
rect 2685 25103 2743 25109
rect 2866 25100 2872 25112
rect 2924 25100 2930 25152
rect 3421 25143 3479 25149
rect 3421 25109 3433 25143
rect 3467 25140 3479 25143
rect 3878 25140 3884 25152
rect 3467 25112 3884 25140
rect 3467 25109 3479 25112
rect 3421 25103 3479 25109
rect 3878 25100 3884 25112
rect 3936 25140 3942 25152
rect 4801 25143 4859 25149
rect 4801 25140 4813 25143
rect 3936 25112 4813 25140
rect 3936 25100 3942 25112
rect 4801 25109 4813 25112
rect 4847 25109 4859 25143
rect 4801 25103 4859 25109
rect 5534 25100 5540 25152
rect 5592 25140 5598 25152
rect 5813 25143 5871 25149
rect 5813 25140 5825 25143
rect 5592 25112 5825 25140
rect 5592 25100 5598 25112
rect 5813 25109 5825 25112
rect 5859 25109 5871 25143
rect 5813 25103 5871 25109
rect 10781 25143 10839 25149
rect 10781 25109 10793 25143
rect 10827 25140 10839 25143
rect 11606 25140 11612 25152
rect 10827 25112 11612 25140
rect 10827 25109 10839 25112
rect 10781 25103 10839 25109
rect 11606 25100 11612 25112
rect 11664 25100 11670 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 4890 24936 4896 24948
rect 4851 24908 4896 24936
rect 4890 24896 4896 24908
rect 4948 24896 4954 24948
rect 5166 24896 5172 24948
rect 5224 24936 5230 24948
rect 11606 24936 11612 24948
rect 5224 24908 11612 24936
rect 5224 24896 5230 24908
rect 11606 24896 11612 24908
rect 11664 24896 11670 24948
rect 2314 24828 2320 24880
rect 2372 24868 2378 24880
rect 2685 24871 2743 24877
rect 2685 24868 2697 24871
rect 2372 24840 2697 24868
rect 2372 24828 2378 24840
rect 2685 24837 2697 24840
rect 2731 24837 2743 24871
rect 2685 24831 2743 24837
rect 3234 24828 3240 24880
rect 3292 24868 3298 24880
rect 8113 24871 8171 24877
rect 8113 24868 8125 24871
rect 3292 24840 8125 24868
rect 3292 24828 3298 24840
rect 8113 24837 8125 24840
rect 8159 24837 8171 24871
rect 12986 24868 12992 24880
rect 8113 24831 8171 24837
rect 12176 24840 12992 24868
rect 3878 24800 3884 24812
rect 3839 24772 3884 24800
rect 3878 24760 3884 24772
rect 3936 24760 3942 24812
rect 3970 24760 3976 24812
rect 4028 24800 4034 24812
rect 4028 24772 4073 24800
rect 4028 24760 4034 24772
rect 5442 24760 5448 24812
rect 5500 24800 5506 24812
rect 5721 24803 5779 24809
rect 5721 24800 5733 24803
rect 5500 24772 5733 24800
rect 5500 24760 5506 24772
rect 5721 24769 5733 24772
rect 5767 24769 5779 24803
rect 6270 24800 6276 24812
rect 6231 24772 6276 24800
rect 5721 24763 5779 24769
rect 6270 24760 6276 24772
rect 6328 24760 6334 24812
rect 8846 24800 8852 24812
rect 8807 24772 8852 24800
rect 8846 24760 8852 24772
rect 8904 24800 8910 24812
rect 10229 24803 10287 24809
rect 8904 24772 9076 24800
rect 8904 24760 8910 24772
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 1670 24732 1676 24744
rect 1443 24704 1676 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 1670 24692 1676 24704
rect 1728 24732 1734 24744
rect 2317 24735 2375 24741
rect 2317 24732 2329 24735
rect 1728 24704 2329 24732
rect 1728 24692 1734 24704
rect 2317 24701 2329 24704
rect 2363 24701 2375 24735
rect 2317 24695 2375 24701
rect 3329 24735 3387 24741
rect 3329 24701 3341 24735
rect 3375 24732 3387 24735
rect 3786 24732 3792 24744
rect 3375 24704 3792 24732
rect 3375 24701 3387 24704
rect 3329 24695 3387 24701
rect 3786 24692 3792 24704
rect 3844 24692 3850 24744
rect 5537 24735 5595 24741
rect 5537 24701 5549 24735
rect 5583 24732 5595 24735
rect 6288 24732 6316 24760
rect 6822 24732 6828 24744
rect 5583 24704 6316 24732
rect 6783 24704 6828 24732
rect 5583 24701 5595 24704
rect 5537 24695 5595 24701
rect 6822 24692 6828 24704
rect 6880 24732 6886 24744
rect 7377 24735 7435 24741
rect 7377 24732 7389 24735
rect 6880 24704 7389 24732
rect 6880 24692 6886 24704
rect 7377 24701 7389 24704
rect 7423 24701 7435 24735
rect 7926 24732 7932 24744
rect 7887 24704 7932 24732
rect 7377 24695 7435 24701
rect 7926 24692 7932 24704
rect 7984 24732 7990 24744
rect 9048 24741 9076 24772
rect 10229 24769 10241 24803
rect 10275 24800 10287 24803
rect 11330 24800 11336 24812
rect 10275 24772 11336 24800
rect 10275 24769 10287 24772
rect 10229 24763 10287 24769
rect 11330 24760 11336 24772
rect 11388 24760 11394 24812
rect 11885 24803 11943 24809
rect 11885 24769 11897 24803
rect 11931 24800 11943 24803
rect 12176 24800 12204 24840
rect 12986 24828 12992 24840
rect 13044 24868 13050 24880
rect 13044 24840 13124 24868
rect 13044 24828 13050 24840
rect 11931 24772 12204 24800
rect 12253 24803 12311 24809
rect 11931 24769 11943 24772
rect 11885 24763 11943 24769
rect 12253 24769 12265 24803
rect 12299 24800 12311 24803
rect 12894 24800 12900 24812
rect 12299 24772 12900 24800
rect 12299 24769 12311 24772
rect 12253 24763 12311 24769
rect 12894 24760 12900 24772
rect 12952 24760 12958 24812
rect 13096 24809 13124 24840
rect 13081 24803 13139 24809
rect 13081 24769 13093 24803
rect 13127 24769 13139 24803
rect 13081 24763 13139 24769
rect 8481 24735 8539 24741
rect 8481 24732 8493 24735
rect 7984 24704 8493 24732
rect 7984 24692 7990 24704
rect 8481 24701 8493 24704
rect 8527 24701 8539 24735
rect 8481 24695 8539 24701
rect 9033 24735 9091 24741
rect 9033 24701 9045 24735
rect 9079 24701 9091 24735
rect 9033 24695 9091 24701
rect 12434 24692 12440 24744
rect 12492 24732 12498 24744
rect 12805 24735 12863 24741
rect 12805 24732 12817 24735
rect 12492 24704 12817 24732
rect 12492 24692 12498 24704
rect 12805 24701 12817 24704
rect 12851 24701 12863 24735
rect 12805 24695 12863 24701
rect 5629 24667 5687 24673
rect 5629 24633 5641 24667
rect 5675 24664 5687 24667
rect 6546 24664 6552 24676
rect 5675 24636 6552 24664
rect 5675 24633 5687 24636
rect 5629 24627 5687 24633
rect 6546 24624 6552 24636
rect 6604 24624 6610 24676
rect 10597 24667 10655 24673
rect 10597 24633 10609 24667
rect 10643 24664 10655 24667
rect 11149 24667 11207 24673
rect 11149 24664 11161 24667
rect 10643 24636 11161 24664
rect 10643 24633 10655 24636
rect 10597 24627 10655 24633
rect 11149 24633 11161 24636
rect 11195 24664 11207 24667
rect 12250 24664 12256 24676
rect 11195 24636 12256 24664
rect 11195 24633 11207 24636
rect 11149 24627 11207 24633
rect 12250 24624 12256 24636
rect 12308 24624 12314 24676
rect 1394 24556 1400 24608
rect 1452 24596 1458 24608
rect 1581 24599 1639 24605
rect 1581 24596 1593 24599
rect 1452 24568 1593 24596
rect 1452 24556 1458 24568
rect 1581 24565 1593 24568
rect 1627 24565 1639 24599
rect 2038 24596 2044 24608
rect 1999 24568 2044 24596
rect 1581 24559 1639 24565
rect 2038 24556 2044 24568
rect 2096 24556 2102 24608
rect 3418 24596 3424 24608
rect 3379 24568 3424 24596
rect 3418 24556 3424 24568
rect 3476 24556 3482 24608
rect 4525 24599 4583 24605
rect 4525 24565 4537 24599
rect 4571 24596 4583 24599
rect 4614 24596 4620 24608
rect 4571 24568 4620 24596
rect 4571 24565 4583 24568
rect 4525 24559 4583 24565
rect 4614 24556 4620 24568
rect 4672 24556 4678 24608
rect 5166 24596 5172 24608
rect 5127 24568 5172 24596
rect 5166 24556 5172 24568
rect 5224 24556 5230 24608
rect 7006 24596 7012 24608
rect 6967 24568 7012 24596
rect 7006 24556 7012 24568
rect 7064 24556 7070 24608
rect 7837 24599 7895 24605
rect 7837 24565 7849 24599
rect 7883 24596 7895 24599
rect 8202 24596 8208 24608
rect 7883 24568 8208 24596
rect 7883 24565 7895 24568
rect 7837 24559 7895 24565
rect 8202 24556 8208 24568
rect 8260 24556 8266 24608
rect 9214 24596 9220 24608
rect 9175 24568 9220 24596
rect 9214 24556 9220 24568
rect 9272 24556 9278 24608
rect 9766 24596 9772 24608
rect 9727 24568 9772 24596
rect 9766 24556 9772 24568
rect 9824 24556 9830 24608
rect 10686 24596 10692 24608
rect 10647 24568 10692 24596
rect 10686 24556 10692 24568
rect 10744 24556 10750 24608
rect 11057 24599 11115 24605
rect 11057 24565 11069 24599
rect 11103 24596 11115 24599
rect 11606 24596 11612 24608
rect 11103 24568 11612 24596
rect 11103 24565 11115 24568
rect 11057 24559 11115 24565
rect 11606 24556 11612 24568
rect 11664 24556 11670 24608
rect 12437 24599 12495 24605
rect 12437 24565 12449 24599
rect 12483 24596 12495 24599
rect 12802 24596 12808 24608
rect 12483 24568 12808 24596
rect 12483 24565 12495 24568
rect 12437 24559 12495 24565
rect 12802 24556 12808 24568
rect 12860 24556 12866 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 3513 24395 3571 24401
rect 3513 24361 3525 24395
rect 3559 24392 3571 24395
rect 3970 24392 3976 24404
rect 3559 24364 3976 24392
rect 3559 24361 3571 24364
rect 3513 24355 3571 24361
rect 3970 24352 3976 24364
rect 4028 24352 4034 24404
rect 6546 24352 6552 24404
rect 6604 24392 6610 24404
rect 7653 24395 7711 24401
rect 7653 24392 7665 24395
rect 6604 24364 7665 24392
rect 6604 24352 6610 24364
rect 7653 24361 7665 24364
rect 7699 24361 7711 24395
rect 8110 24392 8116 24404
rect 8071 24364 8116 24392
rect 7653 24355 7711 24361
rect 8110 24352 8116 24364
rect 8168 24352 8174 24404
rect 10045 24395 10103 24401
rect 10045 24361 10057 24395
rect 10091 24392 10103 24395
rect 10686 24392 10692 24404
rect 10091 24364 10692 24392
rect 10091 24361 10103 24364
rect 10045 24355 10103 24361
rect 10686 24352 10692 24364
rect 10744 24352 10750 24404
rect 12802 24352 12808 24404
rect 12860 24392 12866 24404
rect 13081 24395 13139 24401
rect 13081 24392 13093 24395
rect 12860 24364 13093 24392
rect 12860 24352 12866 24364
rect 13081 24361 13093 24364
rect 13127 24361 13139 24395
rect 14182 24392 14188 24404
rect 14143 24364 14188 24392
rect 13081 24355 13139 24361
rect 14182 24352 14188 24364
rect 14240 24352 14246 24404
rect 16758 24392 16764 24404
rect 16719 24364 16764 24392
rect 16758 24352 16764 24364
rect 16816 24352 16822 24404
rect 17862 24392 17868 24404
rect 17823 24364 17868 24392
rect 17862 24352 17868 24364
rect 17920 24352 17926 24404
rect 19058 24392 19064 24404
rect 19019 24364 19064 24392
rect 19058 24352 19064 24364
rect 19116 24352 19122 24404
rect 21085 24395 21143 24401
rect 21085 24361 21097 24395
rect 21131 24392 21143 24395
rect 22462 24392 22468 24404
rect 21131 24364 22468 24392
rect 21131 24361 21143 24364
rect 21085 24355 21143 24361
rect 22462 24352 22468 24364
rect 22520 24352 22526 24404
rect 1854 24324 1860 24336
rect 1815 24296 1860 24324
rect 1854 24284 1860 24296
rect 1912 24284 1918 24336
rect 3786 24284 3792 24336
rect 3844 24324 3850 24336
rect 5994 24324 6000 24336
rect 3844 24296 6000 24324
rect 3844 24284 3850 24296
rect 1578 24256 1584 24268
rect 1539 24228 1584 24256
rect 1578 24216 1584 24228
rect 1636 24216 1642 24268
rect 2869 24259 2927 24265
rect 2869 24225 2881 24259
rect 2915 24256 2927 24259
rect 2958 24256 2964 24268
rect 2915 24228 2964 24256
rect 2915 24225 2927 24228
rect 2869 24219 2927 24225
rect 2958 24216 2964 24228
rect 3016 24216 3022 24268
rect 3878 24216 3884 24268
rect 3936 24256 3942 24268
rect 5184 24265 5212 24296
rect 5994 24284 6000 24296
rect 6052 24284 6058 24336
rect 5442 24265 5448 24268
rect 4065 24259 4123 24265
rect 4065 24256 4077 24259
rect 3936 24228 4077 24256
rect 3936 24216 3942 24228
rect 4065 24225 4077 24228
rect 4111 24225 4123 24259
rect 4065 24219 4123 24225
rect 5169 24259 5227 24265
rect 5169 24225 5181 24259
rect 5215 24225 5227 24259
rect 5436 24256 5448 24265
rect 5403 24228 5448 24256
rect 5169 24219 5227 24225
rect 5436 24219 5448 24228
rect 5442 24216 5448 24219
rect 5500 24216 5506 24268
rect 7282 24216 7288 24268
rect 7340 24256 7346 24268
rect 8018 24256 8024 24268
rect 7340 24228 8024 24256
rect 7340 24216 7346 24228
rect 8018 24216 8024 24228
rect 8076 24216 8082 24268
rect 10404 24259 10462 24265
rect 10404 24225 10416 24259
rect 10450 24256 10462 24259
rect 11330 24256 11336 24268
rect 10450 24228 11336 24256
rect 10450 24225 10462 24228
rect 10404 24219 10462 24225
rect 11330 24216 11336 24228
rect 11388 24216 11394 24268
rect 12710 24216 12716 24268
rect 12768 24256 12774 24268
rect 12989 24259 13047 24265
rect 12989 24256 13001 24259
rect 12768 24228 13001 24256
rect 12768 24216 12774 24228
rect 12989 24225 13001 24228
rect 13035 24225 13047 24259
rect 12989 24219 13047 24225
rect 16577 24259 16635 24265
rect 16577 24225 16589 24259
rect 16623 24256 16635 24259
rect 16758 24256 16764 24268
rect 16623 24228 16764 24256
rect 16623 24225 16635 24228
rect 16577 24219 16635 24225
rect 16758 24216 16764 24228
rect 16816 24216 16822 24268
rect 17678 24256 17684 24268
rect 17639 24228 17684 24256
rect 17678 24216 17684 24228
rect 17736 24216 17742 24268
rect 18874 24256 18880 24268
rect 18835 24228 18880 24256
rect 18874 24216 18880 24228
rect 18932 24216 18938 24268
rect 20898 24256 20904 24268
rect 20859 24228 20904 24256
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 8202 24148 8208 24200
rect 8260 24188 8266 24200
rect 10134 24188 10140 24200
rect 8260 24160 8305 24188
rect 10095 24160 10140 24188
rect 8260 24148 8266 24160
rect 10134 24148 10140 24160
rect 10192 24148 10198 24200
rect 13265 24191 13323 24197
rect 13265 24157 13277 24191
rect 13311 24188 13323 24191
rect 13311 24160 13768 24188
rect 13311 24157 13323 24160
rect 13265 24151 13323 24157
rect 7561 24123 7619 24129
rect 7561 24089 7573 24123
rect 7607 24120 7619 24123
rect 8220 24120 8248 24148
rect 7607 24092 8248 24120
rect 7607 24089 7619 24092
rect 7561 24083 7619 24089
rect 12342 24080 12348 24132
rect 12400 24120 12406 24132
rect 12621 24123 12679 24129
rect 12621 24120 12633 24123
rect 12400 24092 12633 24120
rect 12400 24080 12406 24092
rect 12621 24089 12633 24092
rect 12667 24089 12679 24123
rect 12621 24083 12679 24089
rect 13740 24064 13768 24160
rect 3050 24052 3056 24064
rect 3011 24024 3056 24052
rect 3050 24012 3056 24024
rect 3108 24012 3114 24064
rect 4246 24052 4252 24064
rect 4207 24024 4252 24052
rect 4246 24012 4252 24024
rect 4304 24012 4310 24064
rect 4893 24055 4951 24061
rect 4893 24021 4905 24055
rect 4939 24052 4951 24055
rect 5074 24052 5080 24064
rect 4939 24024 5080 24052
rect 4939 24021 4951 24024
rect 4893 24015 4951 24021
rect 5074 24012 5080 24024
rect 5132 24052 5138 24064
rect 6549 24055 6607 24061
rect 6549 24052 6561 24055
rect 5132 24024 6561 24052
rect 5132 24012 5138 24024
rect 6549 24021 6561 24024
rect 6595 24021 6607 24055
rect 7098 24052 7104 24064
rect 7059 24024 7104 24052
rect 6549 24015 6607 24021
rect 7098 24012 7104 24024
rect 7156 24012 7162 24064
rect 11514 24052 11520 24064
rect 11475 24024 11520 24052
rect 11514 24012 11520 24024
rect 11572 24012 11578 24064
rect 12434 24012 12440 24064
rect 12492 24052 12498 24064
rect 13722 24052 13728 24064
rect 12492 24024 12537 24052
rect 13683 24024 13728 24052
rect 12492 24012 12498 24024
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 2593 23851 2651 23857
rect 2593 23817 2605 23851
rect 2639 23848 2651 23851
rect 3418 23848 3424 23860
rect 2639 23820 3424 23848
rect 2639 23817 2651 23820
rect 2593 23811 2651 23817
rect 2038 23712 2044 23724
rect 1999 23684 2044 23712
rect 2038 23672 2044 23684
rect 2096 23672 2102 23724
rect 1765 23647 1823 23653
rect 1765 23613 1777 23647
rect 1811 23644 1823 23647
rect 2608 23644 2636 23811
rect 3418 23808 3424 23820
rect 3476 23808 3482 23860
rect 7282 23848 7288 23860
rect 7243 23820 7288 23848
rect 7282 23808 7288 23820
rect 7340 23808 7346 23860
rect 7653 23851 7711 23857
rect 7653 23817 7665 23851
rect 7699 23848 7711 23851
rect 8110 23848 8116 23860
rect 7699 23820 8116 23848
rect 7699 23817 7711 23820
rect 7653 23811 7711 23817
rect 8110 23808 8116 23820
rect 8168 23808 8174 23860
rect 11885 23851 11943 23857
rect 11885 23817 11897 23851
rect 11931 23848 11943 23851
rect 12802 23848 12808 23860
rect 11931 23820 12808 23848
rect 11931 23817 11943 23820
rect 11885 23811 11943 23817
rect 12802 23808 12808 23820
rect 12860 23808 12866 23860
rect 15565 23851 15623 23857
rect 15565 23817 15577 23851
rect 15611 23848 15623 23851
rect 16482 23848 16488 23860
rect 15611 23820 16488 23848
rect 15611 23817 15623 23820
rect 15565 23811 15623 23817
rect 16482 23808 16488 23820
rect 16540 23808 16546 23860
rect 16669 23851 16727 23857
rect 16669 23817 16681 23851
rect 16715 23848 16727 23851
rect 17862 23848 17868 23860
rect 16715 23820 17868 23848
rect 16715 23817 16727 23820
rect 16669 23811 16727 23817
rect 17862 23808 17868 23820
rect 17920 23808 17926 23860
rect 18233 23851 18291 23857
rect 18233 23817 18245 23851
rect 18279 23848 18291 23851
rect 19242 23848 19248 23860
rect 18279 23820 19248 23848
rect 18279 23817 18291 23820
rect 18233 23811 18291 23817
rect 19242 23808 19248 23820
rect 19300 23808 19306 23860
rect 19337 23851 19395 23857
rect 19337 23817 19349 23851
rect 19383 23848 19395 23851
rect 20254 23848 20260 23860
rect 19383 23820 20260 23848
rect 19383 23817 19395 23820
rect 19337 23811 19395 23817
rect 20254 23808 20260 23820
rect 20312 23808 20318 23860
rect 20438 23848 20444 23860
rect 20399 23820 20444 23848
rect 20438 23808 20444 23820
rect 20496 23808 20502 23860
rect 21542 23848 21548 23860
rect 21503 23820 21548 23848
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 9769 23783 9827 23789
rect 9769 23749 9781 23783
rect 9815 23780 9827 23783
rect 12710 23780 12716 23792
rect 9815 23752 10824 23780
rect 12671 23752 12716 23780
rect 9815 23749 9827 23752
rect 9769 23743 9827 23749
rect 10796 23724 10824 23752
rect 12710 23740 12716 23752
rect 12768 23740 12774 23792
rect 3697 23715 3755 23721
rect 3697 23681 3709 23715
rect 3743 23712 3755 23715
rect 10686 23712 10692 23724
rect 3743 23684 3924 23712
rect 10647 23684 10692 23712
rect 3743 23681 3755 23684
rect 3697 23675 3755 23681
rect 3786 23644 3792 23656
rect 1811 23616 2636 23644
rect 3747 23616 3792 23644
rect 1811 23613 1823 23616
rect 1765 23607 1823 23613
rect 3786 23604 3792 23616
rect 3844 23604 3850 23656
rect 3896 23644 3924 23684
rect 10686 23672 10692 23684
rect 10744 23672 10750 23724
rect 10778 23672 10784 23724
rect 10836 23712 10842 23724
rect 11514 23712 11520 23724
rect 10836 23684 11520 23712
rect 10836 23672 10842 23684
rect 11514 23672 11520 23684
rect 11572 23672 11578 23724
rect 12253 23715 12311 23721
rect 12253 23681 12265 23715
rect 12299 23712 12311 23715
rect 12299 23684 13032 23712
rect 12299 23681 12311 23684
rect 12253 23675 12311 23681
rect 4056 23647 4114 23653
rect 4056 23644 4068 23647
rect 3896 23616 4068 23644
rect 4056 23613 4068 23616
rect 4102 23644 4114 23647
rect 5074 23644 5080 23656
rect 4102 23616 5080 23644
rect 4102 23613 4114 23616
rect 4056 23607 4114 23613
rect 5074 23604 5080 23616
rect 5132 23604 5138 23656
rect 7006 23604 7012 23656
rect 7064 23644 7070 23656
rect 7745 23647 7803 23653
rect 7745 23644 7757 23647
rect 7064 23616 7757 23644
rect 7064 23604 7070 23616
rect 7745 23613 7757 23616
rect 7791 23613 7803 23647
rect 7745 23607 7803 23613
rect 10137 23647 10195 23653
rect 10137 23613 10149 23647
rect 10183 23644 10195 23647
rect 10597 23647 10655 23653
rect 10597 23644 10609 23647
rect 10183 23616 10609 23644
rect 10183 23613 10195 23616
rect 10137 23607 10195 23613
rect 10597 23613 10609 23616
rect 10643 23644 10655 23647
rect 10870 23644 10876 23656
rect 10643 23616 10876 23644
rect 10643 23613 10655 23616
rect 10597 23607 10655 23613
rect 10870 23604 10876 23616
rect 10928 23604 10934 23656
rect 12618 23604 12624 23656
rect 12676 23644 12682 23656
rect 12897 23647 12955 23653
rect 12897 23644 12909 23647
rect 12676 23616 12909 23644
rect 12676 23604 12682 23616
rect 12897 23613 12909 23616
rect 12943 23613 12955 23647
rect 13004 23644 13032 23684
rect 18322 23672 18328 23724
rect 18380 23712 18386 23724
rect 18874 23712 18880 23724
rect 18380 23684 18880 23712
rect 18380 23672 18386 23684
rect 18874 23672 18880 23684
rect 18932 23712 18938 23724
rect 18969 23715 19027 23721
rect 18969 23712 18981 23715
rect 18932 23684 18981 23712
rect 18932 23672 18938 23684
rect 18969 23681 18981 23684
rect 19015 23681 19027 23715
rect 18969 23675 19027 23681
rect 13164 23647 13222 23653
rect 13164 23644 13176 23647
rect 13004 23616 13176 23644
rect 12897 23607 12955 23613
rect 13164 23613 13176 23616
rect 13210 23644 13222 23647
rect 13722 23644 13728 23656
rect 13210 23616 13728 23644
rect 13210 23613 13222 23616
rect 13164 23607 13222 23613
rect 13722 23604 13728 23616
rect 13780 23604 13786 23656
rect 15381 23647 15439 23653
rect 15381 23613 15393 23647
rect 15427 23644 15439 23647
rect 15470 23644 15476 23656
rect 15427 23616 15476 23644
rect 15427 23613 15439 23616
rect 15381 23607 15439 23613
rect 15470 23604 15476 23616
rect 15528 23644 15534 23656
rect 15933 23647 15991 23653
rect 15933 23644 15945 23647
rect 15528 23616 15945 23644
rect 15528 23604 15534 23616
rect 15933 23613 15945 23616
rect 15979 23613 15991 23647
rect 15933 23607 15991 23613
rect 16114 23604 16120 23656
rect 16172 23644 16178 23656
rect 16485 23647 16543 23653
rect 16485 23644 16497 23647
rect 16172 23616 16497 23644
rect 16172 23604 16178 23616
rect 16485 23613 16497 23616
rect 16531 23644 16543 23647
rect 17037 23647 17095 23653
rect 17037 23644 17049 23647
rect 16531 23616 17049 23644
rect 16531 23613 16543 23616
rect 16485 23607 16543 23613
rect 17037 23613 17049 23616
rect 17083 23613 17095 23647
rect 17037 23607 17095 23613
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23644 18107 23647
rect 19150 23644 19156 23656
rect 18095 23616 18644 23644
rect 19111 23616 19156 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 2498 23536 2504 23588
rect 2556 23576 2562 23588
rect 3237 23579 3295 23585
rect 3237 23576 3249 23579
rect 2556 23548 3249 23576
rect 2556 23536 2562 23548
rect 3237 23545 3249 23548
rect 3283 23576 3295 23579
rect 3878 23576 3884 23588
rect 3283 23548 3884 23576
rect 3283 23545 3295 23548
rect 3237 23539 3295 23545
rect 3878 23536 3884 23548
rect 3936 23536 3942 23588
rect 4798 23536 4804 23588
rect 4856 23576 4862 23588
rect 5350 23576 5356 23588
rect 4856 23548 5356 23576
rect 4856 23536 4862 23548
rect 5350 23536 5356 23548
rect 5408 23536 5414 23588
rect 5442 23536 5448 23588
rect 5500 23576 5506 23588
rect 5813 23579 5871 23585
rect 5813 23576 5825 23579
rect 5500 23548 5825 23576
rect 5500 23536 5506 23548
rect 5813 23545 5825 23548
rect 5859 23576 5871 23579
rect 8012 23579 8070 23585
rect 5859 23548 7788 23576
rect 5859 23545 5871 23548
rect 5813 23539 5871 23545
rect 2222 23468 2228 23520
rect 2280 23508 2286 23520
rect 2869 23511 2927 23517
rect 2869 23508 2881 23511
rect 2280 23480 2881 23508
rect 2280 23468 2286 23480
rect 2869 23477 2881 23480
rect 2915 23508 2927 23511
rect 2958 23508 2964 23520
rect 2915 23480 2964 23508
rect 2915 23477 2927 23480
rect 2869 23471 2927 23477
rect 2958 23468 2964 23480
rect 3016 23468 3022 23520
rect 4154 23468 4160 23520
rect 4212 23508 4218 23520
rect 5169 23511 5227 23517
rect 5169 23508 5181 23511
rect 4212 23480 5181 23508
rect 4212 23468 4218 23480
rect 5169 23477 5181 23480
rect 5215 23477 5227 23511
rect 5169 23471 5227 23477
rect 5994 23468 6000 23520
rect 6052 23508 6058 23520
rect 6089 23511 6147 23517
rect 6089 23508 6101 23511
rect 6052 23480 6101 23508
rect 6052 23468 6058 23480
rect 6089 23477 6101 23480
rect 6135 23508 6147 23511
rect 6549 23511 6607 23517
rect 6549 23508 6561 23511
rect 6135 23480 6561 23508
rect 6135 23477 6147 23480
rect 6089 23471 6147 23477
rect 6549 23477 6561 23480
rect 6595 23477 6607 23511
rect 7760 23508 7788 23548
rect 8012 23545 8024 23579
rect 8058 23576 8070 23579
rect 8202 23576 8208 23588
rect 8058 23548 8208 23576
rect 8058 23545 8070 23548
rect 8012 23539 8070 23545
rect 8202 23536 8208 23548
rect 8260 23536 8266 23588
rect 16393 23579 16451 23585
rect 16393 23545 16405 23579
rect 16439 23576 16451 23579
rect 16758 23576 16764 23588
rect 16439 23548 16764 23576
rect 16439 23545 16451 23548
rect 16393 23539 16451 23545
rect 16758 23536 16764 23548
rect 16816 23536 16822 23588
rect 18616 23520 18644 23616
rect 19150 23604 19156 23616
rect 19208 23644 19214 23656
rect 19705 23647 19763 23653
rect 19705 23644 19717 23647
rect 19208 23616 19717 23644
rect 19208 23604 19214 23616
rect 19705 23613 19717 23616
rect 19751 23613 19763 23647
rect 20254 23644 20260 23656
rect 20215 23616 20260 23644
rect 19705 23607 19763 23613
rect 20254 23604 20260 23616
rect 20312 23644 20318 23656
rect 20809 23647 20867 23653
rect 20809 23644 20821 23647
rect 20312 23616 20821 23644
rect 20312 23604 20318 23616
rect 20809 23613 20821 23616
rect 20855 23613 20867 23647
rect 21358 23644 21364 23656
rect 21319 23616 21364 23644
rect 20809 23607 20867 23613
rect 21358 23604 21364 23616
rect 21416 23644 21422 23656
rect 21913 23647 21971 23653
rect 21913 23644 21925 23647
rect 21416 23616 21925 23644
rect 21416 23604 21422 23616
rect 21913 23613 21925 23616
rect 21959 23613 21971 23647
rect 21913 23607 21971 23613
rect 23474 23536 23480 23588
rect 23532 23576 23538 23588
rect 24762 23576 24768 23588
rect 23532 23548 24768 23576
rect 23532 23536 23538 23548
rect 24762 23536 24768 23548
rect 24820 23536 24826 23588
rect 9125 23511 9183 23517
rect 9125 23508 9137 23511
rect 7760 23480 9137 23508
rect 6549 23471 6607 23477
rect 9125 23477 9137 23480
rect 9171 23477 9183 23511
rect 9125 23471 9183 23477
rect 9674 23468 9680 23520
rect 9732 23508 9738 23520
rect 10229 23511 10287 23517
rect 10229 23508 10241 23511
rect 9732 23480 10241 23508
rect 9732 23468 9738 23480
rect 10229 23477 10241 23480
rect 10275 23477 10287 23511
rect 11330 23508 11336 23520
rect 11243 23480 11336 23508
rect 10229 23471 10287 23477
rect 11330 23468 11336 23480
rect 11388 23508 11394 23520
rect 14277 23511 14335 23517
rect 14277 23508 14289 23511
rect 11388 23480 14289 23508
rect 11388 23468 11394 23480
rect 14277 23477 14289 23480
rect 14323 23477 14335 23511
rect 14277 23471 14335 23477
rect 16574 23468 16580 23520
rect 16632 23508 16638 23520
rect 17678 23508 17684 23520
rect 16632 23480 17684 23508
rect 16632 23468 16638 23480
rect 17678 23468 17684 23480
rect 17736 23468 17742 23520
rect 18598 23508 18604 23520
rect 18559 23480 18604 23508
rect 18598 23468 18604 23480
rect 18656 23468 18662 23520
rect 20898 23468 20904 23520
rect 20956 23508 20962 23520
rect 21177 23511 21235 23517
rect 21177 23508 21189 23511
rect 20956 23480 21189 23508
rect 20956 23468 20962 23480
rect 21177 23477 21189 23480
rect 21223 23477 21235 23511
rect 21177 23471 21235 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 7006 23304 7012 23316
rect 6967 23276 7012 23304
rect 7006 23264 7012 23276
rect 7064 23264 7070 23316
rect 8202 23264 8208 23316
rect 8260 23304 8266 23316
rect 8481 23307 8539 23313
rect 8481 23304 8493 23307
rect 8260 23276 8493 23304
rect 8260 23264 8266 23276
rect 8481 23273 8493 23276
rect 8527 23273 8539 23307
rect 8481 23267 8539 23273
rect 13814 23264 13820 23316
rect 13872 23304 13878 23316
rect 14093 23307 14151 23313
rect 14093 23304 14105 23307
rect 13872 23276 14105 23304
rect 13872 23264 13878 23276
rect 14093 23273 14105 23276
rect 14139 23273 14151 23307
rect 16666 23304 16672 23316
rect 16627 23276 16672 23304
rect 14093 23267 14151 23273
rect 16666 23264 16672 23276
rect 16724 23264 16730 23316
rect 19613 23307 19671 23313
rect 19613 23273 19625 23307
rect 19659 23304 19671 23307
rect 19978 23304 19984 23316
rect 19659 23276 19984 23304
rect 19659 23273 19671 23276
rect 19613 23267 19671 23273
rect 19978 23264 19984 23276
rect 20036 23264 20042 23316
rect 1854 23236 1860 23248
rect 1815 23208 1860 23236
rect 1854 23196 1860 23208
rect 1912 23196 1918 23248
rect 4154 23196 4160 23248
rect 4212 23236 4218 23248
rect 4310 23239 4368 23245
rect 4310 23236 4322 23239
rect 4212 23208 4322 23236
rect 4212 23196 4218 23208
rect 4310 23205 4322 23208
rect 4356 23205 4368 23239
rect 4310 23199 4368 23205
rect 1578 23168 1584 23180
rect 1539 23140 1584 23168
rect 1578 23128 1584 23140
rect 1636 23128 1642 23180
rect 2869 23171 2927 23177
rect 2869 23137 2881 23171
rect 2915 23168 2927 23171
rect 3418 23168 3424 23180
rect 2915 23140 3424 23168
rect 2915 23137 2927 23140
rect 2869 23131 2927 23137
rect 3418 23128 3424 23140
rect 3476 23128 3482 23180
rect 3786 23168 3792 23180
rect 3747 23140 3792 23168
rect 3786 23128 3792 23140
rect 3844 23168 3850 23180
rect 4065 23171 4123 23177
rect 4065 23168 4077 23171
rect 3844 23140 4077 23168
rect 3844 23128 3850 23140
rect 4065 23137 4077 23140
rect 4111 23137 4123 23171
rect 7024 23168 7052 23264
rect 9582 23196 9588 23248
rect 9640 23236 9646 23248
rect 10312 23239 10370 23245
rect 10312 23236 10324 23239
rect 9640 23208 10324 23236
rect 9640 23196 9646 23208
rect 10312 23205 10324 23208
rect 10358 23236 10370 23239
rect 10778 23236 10784 23248
rect 10358 23208 10784 23236
rect 10358 23205 10370 23208
rect 10312 23199 10370 23205
rect 10778 23196 10784 23208
rect 10836 23196 10842 23248
rect 12986 23245 12992 23248
rect 12980 23236 12992 23245
rect 12947 23208 12992 23236
rect 12980 23199 12992 23208
rect 12986 23196 12992 23199
rect 13044 23196 13050 23248
rect 7374 23177 7380 23180
rect 7101 23171 7159 23177
rect 7101 23168 7113 23171
rect 7024 23140 7113 23168
rect 4065 23131 4123 23137
rect 7101 23137 7113 23140
rect 7147 23137 7159 23171
rect 7368 23168 7380 23177
rect 7335 23140 7380 23168
rect 7101 23131 7159 23137
rect 7368 23131 7380 23140
rect 7374 23128 7380 23131
rect 7432 23128 7438 23180
rect 9953 23171 10011 23177
rect 9953 23137 9965 23171
rect 9999 23168 10011 23171
rect 10045 23171 10103 23177
rect 10045 23168 10057 23171
rect 9999 23140 10057 23168
rect 9999 23137 10011 23140
rect 9953 23131 10011 23137
rect 10045 23137 10057 23140
rect 10091 23168 10103 23171
rect 10134 23168 10140 23180
rect 10091 23140 10140 23168
rect 10091 23137 10103 23140
rect 10045 23131 10103 23137
rect 10134 23128 10140 23140
rect 10192 23128 10198 23180
rect 15562 23177 15568 23180
rect 15556 23168 15568 23177
rect 15523 23140 15568 23168
rect 15556 23131 15568 23140
rect 15562 23128 15568 23131
rect 15620 23128 15626 23180
rect 19426 23168 19432 23180
rect 19387 23140 19432 23168
rect 19426 23128 19432 23140
rect 19484 23128 19490 23180
rect 12713 23103 12771 23109
rect 12713 23100 12725 23103
rect 12636 23072 12725 23100
rect 12636 22976 12664 23072
rect 12713 23069 12725 23072
rect 12759 23069 12771 23103
rect 15286 23100 15292 23112
rect 15247 23072 15292 23100
rect 12713 23063 12771 23069
rect 15286 23060 15292 23072
rect 15344 23060 15350 23112
rect 2406 22964 2412 22976
rect 2367 22936 2412 22964
rect 2406 22924 2412 22936
rect 2464 22924 2470 22976
rect 2866 22924 2872 22976
rect 2924 22964 2930 22976
rect 3053 22967 3111 22973
rect 3053 22964 3065 22967
rect 2924 22936 3065 22964
rect 2924 22924 2930 22936
rect 3053 22933 3065 22936
rect 3099 22933 3111 22967
rect 3053 22927 3111 22933
rect 3234 22924 3240 22976
rect 3292 22964 3298 22976
rect 3421 22967 3479 22973
rect 3421 22964 3433 22967
rect 3292 22936 3433 22964
rect 3292 22924 3298 22936
rect 3421 22933 3433 22936
rect 3467 22933 3479 22967
rect 3421 22927 3479 22933
rect 5258 22924 5264 22976
rect 5316 22964 5322 22976
rect 5445 22967 5503 22973
rect 5445 22964 5457 22967
rect 5316 22936 5457 22964
rect 5316 22924 5322 22936
rect 5445 22933 5457 22936
rect 5491 22933 5503 22967
rect 5445 22927 5503 22933
rect 10686 22924 10692 22976
rect 10744 22964 10750 22976
rect 11425 22967 11483 22973
rect 11425 22964 11437 22967
rect 10744 22936 11437 22964
rect 10744 22924 10750 22936
rect 11425 22933 11437 22936
rect 11471 22933 11483 22967
rect 12618 22964 12624 22976
rect 12579 22936 12624 22964
rect 11425 22927 11483 22933
rect 12618 22924 12624 22936
rect 12676 22924 12682 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1578 22720 1584 22772
rect 1636 22760 1642 22772
rect 2590 22760 2596 22772
rect 1636 22732 2596 22760
rect 1636 22720 1642 22732
rect 2590 22720 2596 22732
rect 2648 22760 2654 22772
rect 2777 22763 2835 22769
rect 2777 22760 2789 22763
rect 2648 22732 2789 22760
rect 2648 22720 2654 22732
rect 2777 22729 2789 22732
rect 2823 22729 2835 22763
rect 4154 22760 4160 22772
rect 4115 22732 4160 22760
rect 2777 22723 2835 22729
rect 4154 22720 4160 22732
rect 4212 22720 4218 22772
rect 5166 22760 5172 22772
rect 5127 22732 5172 22760
rect 5166 22720 5172 22732
rect 5224 22720 5230 22772
rect 9582 22760 9588 22772
rect 9543 22732 9588 22760
rect 9582 22720 9588 22732
rect 9640 22720 9646 22772
rect 12986 22760 12992 22772
rect 12947 22732 12992 22760
rect 12986 22720 12992 22732
rect 13044 22720 13050 22772
rect 2317 22695 2375 22701
rect 2317 22661 2329 22695
rect 2363 22692 2375 22695
rect 2363 22664 3372 22692
rect 2363 22661 2375 22664
rect 2317 22655 2375 22661
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 2498 22624 2504 22636
rect 1811 22596 2504 22624
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 2498 22584 2504 22596
rect 2556 22584 2562 22636
rect 3234 22624 3240 22636
rect 3195 22596 3240 22624
rect 3234 22584 3240 22596
rect 3292 22584 3298 22636
rect 3344 22633 3372 22664
rect 3329 22627 3387 22633
rect 3329 22593 3341 22627
rect 3375 22624 3387 22627
rect 4062 22624 4068 22636
rect 3375 22596 4068 22624
rect 3375 22593 3387 22596
rect 3329 22587 3387 22593
rect 4062 22584 4068 22596
rect 4120 22584 4126 22636
rect 5442 22584 5448 22636
rect 5500 22624 5506 22636
rect 5813 22627 5871 22633
rect 5813 22624 5825 22627
rect 5500 22596 5825 22624
rect 5500 22584 5506 22596
rect 5813 22593 5825 22596
rect 5859 22624 5871 22627
rect 6917 22627 6975 22633
rect 6917 22624 6929 22627
rect 5859 22596 6929 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 6917 22593 6929 22596
rect 6963 22593 6975 22627
rect 6917 22587 6975 22593
rect 7006 22584 7012 22636
rect 7064 22624 7070 22636
rect 7193 22627 7251 22633
rect 7193 22624 7205 22627
rect 7064 22596 7205 22624
rect 7064 22584 7070 22596
rect 7193 22593 7205 22596
rect 7239 22593 7251 22627
rect 7193 22587 7251 22593
rect 9217 22627 9275 22633
rect 9217 22593 9229 22627
rect 9263 22624 9275 22627
rect 10686 22624 10692 22636
rect 9263 22596 10692 22624
rect 9263 22593 9275 22596
rect 9217 22587 9275 22593
rect 10686 22584 10692 22596
rect 10744 22584 10750 22636
rect 12437 22627 12495 22633
rect 12437 22593 12449 22627
rect 12483 22624 12495 22627
rect 12710 22624 12716 22636
rect 12483 22596 12716 22624
rect 12483 22593 12495 22596
rect 12437 22587 12495 22593
rect 12710 22584 12716 22596
rect 12768 22584 12774 22636
rect 1489 22559 1547 22565
rect 1489 22525 1501 22559
rect 1535 22556 1547 22559
rect 2406 22556 2412 22568
rect 1535 22528 2412 22556
rect 1535 22525 1547 22528
rect 1489 22519 1547 22525
rect 2406 22516 2412 22528
rect 2464 22516 2470 22568
rect 5077 22559 5135 22565
rect 5077 22525 5089 22559
rect 5123 22556 5135 22559
rect 5534 22556 5540 22568
rect 5123 22528 5540 22556
rect 5123 22525 5135 22528
rect 5077 22519 5135 22525
rect 5534 22516 5540 22528
rect 5592 22516 5598 22568
rect 6641 22559 6699 22565
rect 6641 22525 6653 22559
rect 6687 22556 6699 22559
rect 7449 22559 7507 22565
rect 7449 22556 7461 22559
rect 6687 22528 7461 22556
rect 6687 22525 6699 22528
rect 6641 22519 6699 22525
rect 7449 22525 7461 22528
rect 7495 22556 7507 22559
rect 8018 22556 8024 22568
rect 7495 22528 8024 22556
rect 7495 22525 7507 22528
rect 7449 22519 7507 22525
rect 8018 22516 8024 22528
rect 8076 22516 8082 22568
rect 9953 22559 10011 22565
rect 9953 22525 9965 22559
rect 9999 22556 10011 22559
rect 10505 22559 10563 22565
rect 10505 22556 10517 22559
rect 9999 22528 10517 22556
rect 9999 22525 10011 22528
rect 9953 22519 10011 22525
rect 10505 22525 10517 22528
rect 10551 22556 10563 22559
rect 10870 22556 10876 22568
rect 10551 22528 10876 22556
rect 10551 22525 10563 22528
rect 10505 22519 10563 22525
rect 10870 22516 10876 22528
rect 10928 22516 10934 22568
rect 10962 22516 10968 22568
rect 11020 22556 11026 22568
rect 11149 22559 11207 22565
rect 11149 22556 11161 22559
rect 11020 22528 11161 22556
rect 11020 22516 11026 22528
rect 11149 22525 11161 22528
rect 11195 22556 11207 22559
rect 12253 22559 12311 22565
rect 12253 22556 12265 22559
rect 11195 22528 12265 22556
rect 11195 22525 11207 22528
rect 11149 22519 11207 22525
rect 12253 22525 12265 22528
rect 12299 22556 12311 22559
rect 12618 22556 12624 22568
rect 12299 22528 12624 22556
rect 12299 22525 12311 22528
rect 12253 22519 12311 22525
rect 12618 22516 12624 22528
rect 12676 22556 12682 22568
rect 13630 22556 13636 22568
rect 12676 22528 13636 22556
rect 12676 22516 12682 22528
rect 13630 22516 13636 22528
rect 13688 22556 13694 22568
rect 13725 22559 13783 22565
rect 13725 22556 13737 22559
rect 13688 22528 13737 22556
rect 13688 22516 13694 22528
rect 13725 22525 13737 22528
rect 13771 22525 13783 22559
rect 13725 22519 13783 22525
rect 15286 22516 15292 22568
rect 15344 22556 15350 22568
rect 16025 22559 16083 22565
rect 16025 22556 16037 22559
rect 15344 22528 16037 22556
rect 15344 22516 15350 22528
rect 16025 22525 16037 22528
rect 16071 22525 16083 22559
rect 16025 22519 16083 22525
rect 2685 22491 2743 22497
rect 2685 22457 2697 22491
rect 2731 22488 2743 22491
rect 3142 22488 3148 22500
rect 2731 22460 3148 22488
rect 2731 22457 2743 22460
rect 2685 22451 2743 22457
rect 3142 22448 3148 22460
rect 3200 22448 3206 22500
rect 4709 22491 4767 22497
rect 4709 22457 4721 22491
rect 4755 22488 4767 22491
rect 5629 22491 5687 22497
rect 5629 22488 5641 22491
rect 4755 22460 5641 22488
rect 4755 22457 4767 22460
rect 4709 22451 4767 22457
rect 5629 22457 5641 22460
rect 5675 22488 5687 22491
rect 6822 22488 6828 22500
rect 5675 22460 6828 22488
rect 5675 22457 5687 22460
rect 5629 22451 5687 22457
rect 6822 22448 6828 22460
rect 6880 22448 6886 22500
rect 6917 22491 6975 22497
rect 6917 22457 6929 22491
rect 6963 22488 6975 22491
rect 6963 22460 7144 22488
rect 6963 22457 6975 22460
rect 6917 22451 6975 22457
rect 5994 22380 6000 22432
rect 6052 22420 6058 22432
rect 6181 22423 6239 22429
rect 6181 22420 6193 22423
rect 6052 22392 6193 22420
rect 6052 22380 6058 22392
rect 6181 22389 6193 22392
rect 6227 22420 6239 22423
rect 7006 22420 7012 22432
rect 6227 22392 7012 22420
rect 6227 22389 6239 22392
rect 6181 22383 6239 22389
rect 7006 22380 7012 22392
rect 7064 22380 7070 22432
rect 7116 22429 7144 22460
rect 9858 22448 9864 22500
rect 9916 22488 9922 22500
rect 10413 22491 10471 22497
rect 10413 22488 10425 22491
rect 9916 22460 10425 22488
rect 9916 22448 9922 22460
rect 10413 22457 10425 22460
rect 10459 22457 10471 22491
rect 13970 22491 14028 22497
rect 13970 22488 13982 22491
rect 10413 22451 10471 22457
rect 13556 22460 13982 22488
rect 13556 22432 13584 22460
rect 13970 22457 13982 22460
rect 14016 22457 14028 22491
rect 13970 22451 14028 22457
rect 7101 22423 7159 22429
rect 7101 22389 7113 22423
rect 7147 22420 7159 22423
rect 7374 22420 7380 22432
rect 7147 22392 7380 22420
rect 7147 22389 7159 22392
rect 7101 22383 7159 22389
rect 7374 22380 7380 22392
rect 7432 22420 7438 22432
rect 8573 22423 8631 22429
rect 8573 22420 8585 22423
rect 7432 22392 8585 22420
rect 7432 22380 7438 22392
rect 8573 22389 8585 22392
rect 8619 22389 8631 22423
rect 8573 22383 8631 22389
rect 9950 22380 9956 22432
rect 10008 22420 10014 22432
rect 10045 22423 10103 22429
rect 10045 22420 10057 22423
rect 10008 22392 10057 22420
rect 10008 22380 10014 22392
rect 10045 22389 10057 22392
rect 10091 22389 10103 22423
rect 13538 22420 13544 22432
rect 13499 22392 13544 22420
rect 10045 22383 10103 22389
rect 13538 22380 13544 22392
rect 13596 22380 13602 22432
rect 13814 22380 13820 22432
rect 13872 22420 13878 22432
rect 15105 22423 15163 22429
rect 15105 22420 15117 22423
rect 13872 22392 15117 22420
rect 13872 22380 13878 22392
rect 15105 22389 15117 22392
rect 15151 22420 15163 22423
rect 15562 22420 15568 22432
rect 15151 22392 15568 22420
rect 15151 22389 15163 22392
rect 15105 22383 15163 22389
rect 15562 22380 15568 22392
rect 15620 22420 15626 22432
rect 15657 22423 15715 22429
rect 15657 22420 15669 22423
rect 15620 22392 15669 22420
rect 15620 22380 15626 22392
rect 15657 22389 15669 22392
rect 15703 22389 15715 22423
rect 19426 22420 19432 22432
rect 19387 22392 19432 22420
rect 15657 22383 15715 22389
rect 19426 22380 19432 22392
rect 19484 22380 19490 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 2590 22216 2596 22228
rect 2551 22188 2596 22216
rect 2590 22176 2596 22188
rect 2648 22176 2654 22228
rect 3234 22176 3240 22228
rect 3292 22216 3298 22228
rect 4065 22219 4123 22225
rect 4065 22216 4077 22219
rect 3292 22188 4077 22216
rect 3292 22176 3298 22188
rect 4065 22185 4077 22188
rect 4111 22185 4123 22219
rect 4065 22179 4123 22185
rect 9858 22176 9864 22228
rect 9916 22216 9922 22228
rect 10045 22219 10103 22225
rect 10045 22216 10057 22219
rect 9916 22188 10057 22216
rect 9916 22176 9922 22188
rect 10045 22185 10057 22188
rect 10091 22185 10103 22219
rect 10045 22179 10103 22185
rect 15289 22219 15347 22225
rect 15289 22185 15301 22219
rect 15335 22216 15347 22219
rect 15378 22216 15384 22228
rect 15335 22188 15384 22216
rect 15335 22185 15347 22188
rect 15289 22179 15347 22185
rect 15378 22176 15384 22188
rect 15436 22176 15442 22228
rect 16298 22216 16304 22228
rect 16259 22188 16304 22216
rect 16298 22176 16304 22188
rect 16356 22176 16362 22228
rect 3786 22148 3792 22160
rect 3747 22120 3792 22148
rect 3786 22108 3792 22120
rect 3844 22108 3850 22160
rect 8202 22148 8208 22160
rect 8163 22120 8208 22148
rect 8202 22108 8208 22120
rect 8260 22108 8266 22160
rect 10496 22151 10554 22157
rect 10496 22117 10508 22151
rect 10542 22148 10554 22151
rect 10686 22148 10692 22160
rect 10542 22120 10692 22148
rect 10542 22117 10554 22120
rect 10496 22111 10554 22117
rect 10686 22108 10692 22120
rect 10744 22108 10750 22160
rect 13630 22108 13636 22160
rect 13688 22108 13694 22160
rect 15194 22148 15200 22160
rect 15120 22120 15200 22148
rect 1489 22083 1547 22089
rect 1489 22049 1501 22083
rect 1535 22049 1547 22083
rect 1489 22043 1547 22049
rect 1765 22083 1823 22089
rect 1765 22049 1777 22083
rect 1811 22080 1823 22083
rect 2314 22080 2320 22092
rect 1811 22052 2320 22080
rect 1811 22049 1823 22052
rect 1765 22043 1823 22049
rect 1504 22012 1532 22043
rect 2314 22040 2320 22052
rect 2372 22040 2378 22092
rect 2774 22080 2780 22092
rect 2735 22052 2780 22080
rect 2774 22040 2780 22052
rect 2832 22040 2838 22092
rect 4430 22080 4436 22092
rect 4391 22052 4436 22080
rect 4430 22040 4436 22052
rect 4488 22040 4494 22092
rect 4522 22040 4528 22092
rect 4580 22080 4586 22092
rect 5261 22083 5319 22089
rect 4580 22052 4625 22080
rect 4580 22040 4586 22052
rect 5261 22049 5273 22083
rect 5307 22080 5319 22083
rect 5442 22080 5448 22092
rect 5307 22052 5448 22080
rect 5307 22049 5319 22052
rect 5261 22043 5319 22049
rect 5442 22040 5448 22052
rect 5500 22040 5506 22092
rect 6178 22040 6184 22092
rect 6236 22080 6242 22092
rect 6641 22083 6699 22089
rect 6641 22080 6653 22083
rect 6236 22052 6653 22080
rect 6236 22040 6242 22052
rect 6641 22049 6653 22052
rect 6687 22049 6699 22083
rect 6641 22043 6699 22049
rect 8297 22083 8355 22089
rect 8297 22049 8309 22083
rect 8343 22080 8355 22083
rect 8754 22080 8760 22092
rect 8343 22052 8760 22080
rect 8343 22049 8355 22052
rect 8297 22043 8355 22049
rect 8754 22040 8760 22052
rect 8812 22040 8818 22092
rect 10134 22040 10140 22092
rect 10192 22080 10198 22092
rect 10229 22083 10287 22089
rect 10229 22080 10241 22083
rect 10192 22052 10241 22080
rect 10192 22040 10198 22052
rect 10229 22049 10241 22052
rect 10275 22080 10287 22083
rect 10962 22080 10968 22092
rect 10275 22052 10968 22080
rect 10275 22049 10287 22052
rect 10229 22043 10287 22049
rect 10962 22040 10968 22052
rect 11020 22040 11026 22092
rect 13170 22080 13176 22092
rect 13131 22052 13176 22080
rect 13170 22040 13176 22052
rect 13228 22040 13234 22092
rect 13648 22080 13676 22108
rect 13909 22083 13967 22089
rect 13909 22080 13921 22083
rect 13648 22052 13921 22080
rect 13909 22049 13921 22052
rect 13955 22080 13967 22083
rect 14277 22083 14335 22089
rect 14277 22080 14289 22083
rect 13955 22052 14289 22080
rect 13955 22049 13967 22052
rect 13909 22043 13967 22049
rect 14277 22049 14289 22052
rect 14323 22080 14335 22083
rect 15120 22080 15148 22120
rect 15194 22108 15200 22120
rect 15252 22108 15258 22160
rect 14323 22052 15148 22080
rect 14323 22049 14335 22052
rect 14277 22043 14335 22049
rect 2406 22012 2412 22024
rect 1504 21984 2412 22012
rect 2406 21972 2412 21984
rect 2464 21972 2470 22024
rect 4709 22015 4767 22021
rect 4709 21981 4721 22015
rect 4755 22012 4767 22015
rect 5166 22012 5172 22024
rect 4755 21984 5172 22012
rect 4755 21981 4767 21984
rect 4709 21975 4767 21981
rect 5166 21972 5172 21984
rect 5224 21972 5230 22024
rect 6730 22012 6736 22024
rect 6691 21984 6736 22012
rect 6730 21972 6736 21984
rect 6788 21972 6794 22024
rect 6825 22015 6883 22021
rect 6825 21981 6837 22015
rect 6871 22012 6883 22015
rect 7006 22012 7012 22024
rect 6871 21984 7012 22012
rect 6871 21981 6883 21984
rect 6825 21975 6883 21981
rect 7006 21972 7012 21984
rect 7064 21972 7070 22024
rect 8018 21972 8024 22024
rect 8076 22012 8082 22024
rect 8389 22015 8447 22021
rect 8389 22012 8401 22015
rect 8076 21984 8401 22012
rect 8076 21972 8082 21984
rect 8389 21981 8401 21984
rect 8435 22012 8447 22015
rect 8849 22015 8907 22021
rect 8849 22012 8861 22015
rect 8435 21984 8861 22012
rect 8435 21981 8447 21984
rect 8389 21975 8447 21981
rect 8849 21981 8861 21984
rect 8895 21981 8907 22015
rect 8849 21975 8907 21981
rect 12713 22015 12771 22021
rect 12713 21981 12725 22015
rect 12759 22012 12771 22015
rect 12894 22012 12900 22024
rect 12759 21984 12900 22012
rect 12759 21981 12771 21984
rect 12713 21975 12771 21981
rect 12894 21972 12900 21984
rect 12952 22012 12958 22024
rect 13265 22015 13323 22021
rect 13265 22012 13277 22015
rect 12952 21984 13277 22012
rect 12952 21972 12958 21984
rect 13265 21981 13277 21984
rect 13311 21981 13323 22015
rect 13265 21975 13323 21981
rect 13449 22015 13507 22021
rect 13449 21981 13461 22015
rect 13495 22012 13507 22015
rect 13722 22012 13728 22024
rect 13495 21984 13728 22012
rect 13495 21981 13507 21984
rect 13449 21975 13507 21981
rect 2314 21944 2320 21956
rect 2275 21916 2320 21944
rect 2314 21904 2320 21916
rect 2372 21904 2378 21956
rect 2958 21944 2964 21956
rect 2919 21916 2964 21944
rect 2958 21904 2964 21916
rect 3016 21904 3022 21956
rect 6914 21904 6920 21956
rect 6972 21944 6978 21956
rect 7837 21947 7895 21953
rect 7837 21944 7849 21947
rect 6972 21916 7849 21944
rect 6972 21904 6978 21916
rect 7837 21913 7849 21916
rect 7883 21913 7895 21947
rect 7837 21907 7895 21913
rect 12250 21904 12256 21956
rect 12308 21944 12314 21956
rect 13464 21944 13492 21975
rect 13722 21972 13728 21984
rect 13780 21972 13786 22024
rect 12308 21916 13492 21944
rect 12308 21904 12314 21916
rect 3418 21876 3424 21888
rect 3379 21848 3424 21876
rect 3418 21836 3424 21848
rect 3476 21836 3482 21888
rect 5166 21836 5172 21888
rect 5224 21876 5230 21888
rect 5537 21879 5595 21885
rect 5537 21876 5549 21879
rect 5224 21848 5549 21876
rect 5224 21836 5230 21848
rect 5537 21845 5549 21848
rect 5583 21845 5595 21879
rect 5994 21876 6000 21888
rect 5955 21848 6000 21876
rect 5537 21839 5595 21845
rect 5994 21836 6000 21848
rect 6052 21836 6058 21888
rect 6270 21876 6276 21888
rect 6231 21848 6276 21876
rect 6270 21836 6276 21848
rect 6328 21836 6334 21888
rect 7558 21876 7564 21888
rect 7519 21848 7564 21876
rect 7558 21836 7564 21848
rect 7616 21836 7622 21888
rect 10134 21836 10140 21888
rect 10192 21876 10198 21888
rect 11609 21879 11667 21885
rect 11609 21876 11621 21879
rect 10192 21848 11621 21876
rect 10192 21836 10198 21848
rect 11609 21845 11621 21848
rect 11655 21845 11667 21879
rect 12802 21876 12808 21888
rect 12763 21848 12808 21876
rect 11609 21839 11667 21845
rect 12802 21836 12808 21848
rect 12860 21836 12866 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2774 21672 2780 21684
rect 2687 21644 2780 21672
rect 2774 21632 2780 21644
rect 2832 21672 2838 21684
rect 3510 21672 3516 21684
rect 2832 21644 3516 21672
rect 2832 21632 2838 21644
rect 3510 21632 3516 21644
rect 3568 21632 3574 21684
rect 4154 21632 4160 21684
rect 4212 21672 4218 21684
rect 4249 21675 4307 21681
rect 4249 21672 4261 21675
rect 4212 21644 4261 21672
rect 4212 21632 4218 21644
rect 4249 21641 4261 21644
rect 4295 21641 4307 21675
rect 4249 21635 4307 21641
rect 4522 21632 4528 21684
rect 4580 21672 4586 21684
rect 4801 21675 4859 21681
rect 4801 21672 4813 21675
rect 4580 21644 4813 21672
rect 4580 21632 4586 21644
rect 4801 21641 4813 21644
rect 4847 21641 4859 21675
rect 5258 21672 5264 21684
rect 5219 21644 5264 21672
rect 4801 21635 4859 21641
rect 5258 21632 5264 21644
rect 5316 21632 5322 21684
rect 8573 21675 8631 21681
rect 8573 21641 8585 21675
rect 8619 21672 8631 21675
rect 8754 21672 8760 21684
rect 8619 21644 8760 21672
rect 8619 21641 8631 21644
rect 8573 21635 8631 21641
rect 8754 21632 8760 21644
rect 8812 21632 8818 21684
rect 9490 21672 9496 21684
rect 9451 21644 9496 21672
rect 9490 21632 9496 21644
rect 9548 21632 9554 21684
rect 10597 21675 10655 21681
rect 10597 21641 10609 21675
rect 10643 21672 10655 21675
rect 10686 21672 10692 21684
rect 10643 21644 10692 21672
rect 10643 21641 10655 21644
rect 10597 21635 10655 21641
rect 10686 21632 10692 21644
rect 10744 21632 10750 21684
rect 11885 21675 11943 21681
rect 11885 21641 11897 21675
rect 11931 21672 11943 21675
rect 12342 21672 12348 21684
rect 11931 21644 12348 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 6730 21564 6736 21616
rect 6788 21604 6794 21616
rect 7469 21607 7527 21613
rect 7469 21604 7481 21607
rect 6788 21576 7481 21604
rect 6788 21564 6794 21576
rect 7469 21573 7481 21576
rect 7515 21573 7527 21607
rect 7469 21567 7527 21573
rect 8294 21564 8300 21616
rect 8352 21604 8358 21616
rect 8846 21604 8852 21616
rect 8352 21576 8852 21604
rect 8352 21564 8358 21576
rect 8846 21564 8852 21576
rect 8904 21564 8910 21616
rect 10873 21607 10931 21613
rect 10873 21604 10885 21607
rect 9968 21576 10885 21604
rect 9968 21548 9996 21576
rect 10873 21573 10885 21576
rect 10919 21573 10931 21607
rect 10873 21567 10931 21573
rect 1670 21536 1676 21548
rect 1631 21508 1676 21536
rect 1670 21496 1676 21508
rect 1728 21496 1734 21548
rect 2409 21539 2467 21545
rect 2409 21505 2421 21539
rect 2455 21536 2467 21539
rect 7377 21539 7435 21545
rect 2455 21508 3004 21536
rect 2455 21505 2467 21508
rect 2409 21499 2467 21505
rect 1489 21471 1547 21477
rect 1489 21437 1501 21471
rect 1535 21468 1547 21471
rect 2314 21468 2320 21480
rect 1535 21440 2320 21468
rect 1535 21437 1547 21440
rect 1489 21431 1547 21437
rect 2314 21428 2320 21440
rect 2372 21428 2378 21480
rect 2869 21471 2927 21477
rect 2869 21437 2881 21471
rect 2915 21437 2927 21471
rect 2976 21468 3004 21508
rect 7377 21505 7389 21539
rect 7423 21536 7435 21539
rect 7926 21536 7932 21548
rect 7423 21508 7932 21536
rect 7423 21505 7435 21508
rect 7377 21499 7435 21505
rect 7926 21496 7932 21508
rect 7984 21496 7990 21548
rect 8113 21539 8171 21545
rect 8113 21505 8125 21539
rect 8159 21536 8171 21539
rect 8202 21536 8208 21548
rect 8159 21508 8208 21536
rect 8159 21505 8171 21508
rect 8113 21499 8171 21505
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 9950 21536 9956 21548
rect 9911 21508 9956 21536
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 10134 21536 10140 21548
rect 10095 21508 10140 21536
rect 10134 21496 10140 21508
rect 10192 21496 10198 21548
rect 11238 21536 11244 21548
rect 11199 21508 11244 21536
rect 11238 21496 11244 21508
rect 11296 21496 11302 21548
rect 3136 21471 3194 21477
rect 3136 21468 3148 21471
rect 2976 21440 3148 21468
rect 2869 21431 2927 21437
rect 3136 21437 3148 21440
rect 3182 21468 3194 21471
rect 5258 21468 5264 21480
rect 3182 21440 5264 21468
rect 3182 21437 3194 21440
rect 3136 21431 3194 21437
rect 2884 21400 2912 21431
rect 5258 21428 5264 21440
rect 5316 21428 5322 21480
rect 5353 21471 5411 21477
rect 5353 21437 5365 21471
rect 5399 21437 5411 21471
rect 5353 21431 5411 21437
rect 3786 21400 3792 21412
rect 2884 21372 3792 21400
rect 3786 21360 3792 21372
rect 3844 21360 3850 21412
rect 5166 21360 5172 21412
rect 5224 21400 5230 21412
rect 5368 21400 5396 21431
rect 7558 21428 7564 21480
rect 7616 21468 7622 21480
rect 7837 21471 7895 21477
rect 7837 21468 7849 21471
rect 7616 21440 7849 21468
rect 7616 21428 7622 21440
rect 7837 21437 7849 21440
rect 7883 21437 7895 21471
rect 7837 21431 7895 21437
rect 11057 21471 11115 21477
rect 11057 21437 11069 21471
rect 11103 21468 11115 21471
rect 11900 21468 11928 21635
rect 12342 21632 12348 21644
rect 12400 21632 12406 21684
rect 13170 21672 13176 21684
rect 13131 21644 13176 21672
rect 13170 21632 13176 21644
rect 13228 21632 13234 21684
rect 12250 21604 12256 21616
rect 12211 21576 12256 21604
rect 12250 21564 12256 21576
rect 12308 21564 12314 21616
rect 12713 21539 12771 21545
rect 12713 21505 12725 21539
rect 12759 21536 12771 21539
rect 13188 21536 13216 21632
rect 12759 21508 13216 21536
rect 12759 21505 12771 21508
rect 12713 21499 12771 21505
rect 13630 21496 13636 21548
rect 13688 21536 13694 21548
rect 13725 21539 13783 21545
rect 13725 21536 13737 21539
rect 13688 21508 13737 21536
rect 13688 21496 13694 21508
rect 13725 21505 13737 21508
rect 13771 21505 13783 21539
rect 13725 21499 13783 21505
rect 11103 21440 11928 21468
rect 11103 21437 11115 21440
rect 11057 21431 11115 21437
rect 5224 21372 5396 21400
rect 5997 21403 6055 21409
rect 5224 21360 5230 21372
rect 5997 21369 6009 21403
rect 6043 21400 6055 21403
rect 7006 21400 7012 21412
rect 6043 21372 7012 21400
rect 6043 21369 6055 21372
rect 5997 21363 6055 21369
rect 7006 21360 7012 21372
rect 7064 21360 7070 21412
rect 9401 21403 9459 21409
rect 9401 21369 9413 21403
rect 9447 21400 9459 21403
rect 9861 21403 9919 21409
rect 9861 21400 9873 21403
rect 9447 21372 9873 21400
rect 9447 21369 9459 21372
rect 9401 21363 9459 21369
rect 9861 21369 9873 21372
rect 9907 21400 9919 21403
rect 10686 21400 10692 21412
rect 9907 21372 10692 21400
rect 9907 21369 9919 21372
rect 9861 21363 9919 21369
rect 10686 21360 10692 21372
rect 10744 21360 10750 21412
rect 13633 21403 13691 21409
rect 13633 21369 13645 21403
rect 13679 21400 13691 21403
rect 13970 21403 14028 21409
rect 13970 21400 13982 21403
rect 13679 21372 13982 21400
rect 13679 21369 13691 21372
rect 13633 21363 13691 21369
rect 13970 21369 13982 21372
rect 14016 21400 14028 21403
rect 15194 21400 15200 21412
rect 14016 21372 15200 21400
rect 14016 21369 14028 21372
rect 13970 21363 14028 21369
rect 15194 21360 15200 21372
rect 15252 21360 15258 21412
rect 23566 21360 23572 21412
rect 23624 21400 23630 21412
rect 24210 21400 24216 21412
rect 23624 21372 24216 21400
rect 23624 21360 23630 21372
rect 24210 21360 24216 21372
rect 24268 21360 24274 21412
rect 24854 21360 24860 21412
rect 24912 21400 24918 21412
rect 25958 21400 25964 21412
rect 24912 21372 25964 21400
rect 24912 21360 24918 21372
rect 25958 21360 25964 21372
rect 26016 21360 26022 21412
rect 5534 21332 5540 21344
rect 5495 21304 5540 21332
rect 5534 21292 5540 21304
rect 5592 21292 5598 21344
rect 6178 21292 6184 21344
rect 6236 21332 6242 21344
rect 6273 21335 6331 21341
rect 6273 21332 6285 21335
rect 6236 21304 6285 21332
rect 6236 21292 6242 21304
rect 6273 21301 6285 21304
rect 6319 21301 6331 21335
rect 6273 21295 6331 21301
rect 13538 21292 13544 21344
rect 13596 21332 13602 21344
rect 15105 21335 15163 21341
rect 15105 21332 15117 21335
rect 13596 21304 15117 21332
rect 13596 21292 13602 21304
rect 15105 21301 15117 21304
rect 15151 21301 15163 21335
rect 15105 21295 15163 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 2406 21128 2412 21140
rect 2367 21100 2412 21128
rect 2406 21088 2412 21100
rect 2464 21088 2470 21140
rect 3513 21131 3571 21137
rect 3513 21097 3525 21131
rect 3559 21128 3571 21131
rect 3786 21128 3792 21140
rect 3559 21100 3792 21128
rect 3559 21097 3571 21100
rect 3513 21091 3571 21097
rect 3786 21088 3792 21100
rect 3844 21088 3850 21140
rect 6365 21131 6423 21137
rect 6365 21097 6377 21131
rect 6411 21128 6423 21131
rect 6730 21128 6736 21140
rect 6411 21100 6736 21128
rect 6411 21097 6423 21100
rect 6365 21091 6423 21097
rect 6730 21088 6736 21100
rect 6788 21088 6794 21140
rect 8018 21088 8024 21140
rect 8076 21128 8082 21140
rect 8113 21131 8171 21137
rect 8113 21128 8125 21131
rect 8076 21100 8125 21128
rect 8076 21088 8082 21100
rect 8113 21097 8125 21100
rect 8159 21097 8171 21131
rect 12894 21128 12900 21140
rect 12855 21100 12900 21128
rect 8113 21091 8171 21097
rect 12894 21088 12900 21100
rect 12952 21088 12958 21140
rect 13354 21128 13360 21140
rect 13315 21100 13360 21128
rect 13354 21088 13360 21100
rect 13412 21088 13418 21140
rect 13630 21088 13636 21140
rect 13688 21128 13694 21140
rect 13814 21128 13820 21140
rect 13688 21100 13820 21128
rect 13688 21088 13694 21100
rect 13814 21088 13820 21100
rect 13872 21128 13878 21140
rect 14277 21131 14335 21137
rect 14277 21128 14289 21131
rect 13872 21100 14289 21128
rect 13872 21088 13878 21100
rect 14277 21097 14289 21100
rect 14323 21097 14335 21131
rect 15286 21128 15292 21140
rect 15247 21100 15292 21128
rect 14277 21091 14335 21097
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 1857 21063 1915 21069
rect 1857 21029 1869 21063
rect 1903 21060 1915 21063
rect 1946 21060 1952 21072
rect 1903 21032 1952 21060
rect 1903 21029 1915 21032
rect 1857 21023 1915 21029
rect 1946 21020 1952 21032
rect 2004 21020 2010 21072
rect 5077 21063 5135 21069
rect 5077 21029 5089 21063
rect 5123 21060 5135 21063
rect 5258 21060 5264 21072
rect 5123 21032 5264 21060
rect 5123 21029 5135 21032
rect 5077 21023 5135 21029
rect 5258 21020 5264 21032
rect 5316 21020 5322 21072
rect 9953 21063 10011 21069
rect 9953 21029 9965 21063
rect 9999 21060 10011 21063
rect 10134 21060 10140 21072
rect 9999 21032 10140 21060
rect 9999 21029 10011 21032
rect 9953 21023 10011 21029
rect 10134 21020 10140 21032
rect 10192 21060 10198 21072
rect 10290 21063 10348 21069
rect 10290 21060 10302 21063
rect 10192 21032 10302 21060
rect 10192 21020 10198 21032
rect 10290 21029 10302 21032
rect 10336 21029 10348 21063
rect 10290 21023 10348 21029
rect 1581 20995 1639 21001
rect 1581 20961 1593 20995
rect 1627 20992 1639 20995
rect 2682 20992 2688 21004
rect 1627 20964 2688 20992
rect 1627 20961 1639 20964
rect 1581 20955 1639 20961
rect 2682 20952 2688 20964
rect 2740 20952 2746 21004
rect 2869 20995 2927 21001
rect 2869 20961 2881 20995
rect 2915 20992 2927 20995
rect 3050 20992 3056 21004
rect 2915 20964 3056 20992
rect 2915 20961 2927 20964
rect 2869 20955 2927 20961
rect 3050 20952 3056 20964
rect 3108 20952 3114 21004
rect 4985 20995 5043 21001
rect 4985 20961 4997 20995
rect 5031 20992 5043 20995
rect 5442 20992 5448 21004
rect 5031 20964 5448 20992
rect 5031 20961 5043 20964
rect 4985 20955 5043 20961
rect 5442 20952 5448 20964
rect 5500 20952 5506 21004
rect 6641 20995 6699 21001
rect 6641 20961 6653 20995
rect 6687 20992 6699 20995
rect 6822 20992 6828 21004
rect 6687 20964 6828 20992
rect 6687 20961 6699 20964
rect 6641 20955 6699 20961
rect 6822 20952 6828 20964
rect 6880 20952 6886 21004
rect 7006 21001 7012 21004
rect 7000 20992 7012 21001
rect 6967 20964 7012 20992
rect 7000 20955 7012 20964
rect 7006 20952 7012 20955
rect 7064 20952 7070 21004
rect 12434 20952 12440 21004
rect 12492 20992 12498 21004
rect 12713 20995 12771 21001
rect 12713 20992 12725 20995
rect 12492 20964 12725 20992
rect 12492 20952 12498 20964
rect 12713 20961 12725 20964
rect 12759 20961 12771 20995
rect 12713 20955 12771 20961
rect 13170 20952 13176 21004
rect 13228 20992 13234 21004
rect 13265 20995 13323 21001
rect 13265 20992 13277 20995
rect 13228 20964 13277 20992
rect 13228 20952 13234 20964
rect 13265 20961 13277 20964
rect 13311 20961 13323 20995
rect 13265 20955 13323 20961
rect 5166 20924 5172 20936
rect 5127 20896 5172 20924
rect 5166 20884 5172 20896
rect 5224 20884 5230 20936
rect 5994 20924 6000 20936
rect 5907 20896 6000 20924
rect 5994 20884 6000 20896
rect 6052 20924 6058 20936
rect 6730 20924 6736 20936
rect 6052 20896 6736 20924
rect 6052 20884 6058 20896
rect 2777 20859 2835 20865
rect 2777 20825 2789 20859
rect 2823 20856 2835 20859
rect 3789 20859 3847 20865
rect 3789 20856 3801 20859
rect 2823 20828 3801 20856
rect 2823 20825 2835 20828
rect 2777 20819 2835 20825
rect 3789 20825 3801 20828
rect 3835 20856 3847 20859
rect 3970 20856 3976 20868
rect 3835 20828 3976 20856
rect 3835 20825 3847 20828
rect 3789 20819 3847 20825
rect 3970 20816 3976 20828
rect 4028 20816 4034 20868
rect 4341 20859 4399 20865
rect 4341 20825 4353 20859
rect 4387 20856 4399 20859
rect 4430 20856 4436 20868
rect 4387 20828 4436 20856
rect 4387 20825 4399 20828
rect 4341 20819 4399 20825
rect 4430 20816 4436 20828
rect 4488 20856 4494 20868
rect 4890 20856 4896 20868
rect 4488 20828 4896 20856
rect 4488 20816 4494 20828
rect 4890 20816 4896 20828
rect 4948 20816 4954 20868
rect 6472 20865 6500 20896
rect 6730 20884 6736 20896
rect 6788 20884 6794 20936
rect 9493 20927 9551 20933
rect 9493 20893 9505 20927
rect 9539 20924 9551 20927
rect 10042 20924 10048 20936
rect 9539 20896 10048 20924
rect 9539 20893 9551 20896
rect 9493 20887 9551 20893
rect 10042 20884 10048 20896
rect 10100 20884 10106 20936
rect 12986 20884 12992 20936
rect 13044 20924 13050 20936
rect 13449 20927 13507 20933
rect 13449 20924 13461 20927
rect 13044 20896 13461 20924
rect 13044 20884 13050 20896
rect 13449 20893 13461 20896
rect 13495 20924 13507 20927
rect 13538 20924 13544 20936
rect 13495 20896 13544 20924
rect 13495 20893 13507 20896
rect 13449 20887 13507 20893
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 6457 20859 6515 20865
rect 6457 20825 6469 20859
rect 6503 20825 6515 20859
rect 12526 20856 12532 20868
rect 12439 20828 12532 20856
rect 6457 20819 6515 20825
rect 12526 20816 12532 20828
rect 12584 20856 12590 20868
rect 13814 20856 13820 20868
rect 12584 20828 13820 20856
rect 12584 20816 12590 20828
rect 13814 20816 13820 20828
rect 13872 20816 13878 20868
rect 3053 20791 3111 20797
rect 3053 20757 3065 20791
rect 3099 20788 3111 20791
rect 3142 20788 3148 20800
rect 3099 20760 3148 20788
rect 3099 20757 3111 20760
rect 3053 20751 3111 20757
rect 3142 20748 3148 20760
rect 3200 20748 3206 20800
rect 4522 20748 4528 20800
rect 4580 20788 4586 20800
rect 4617 20791 4675 20797
rect 4617 20788 4629 20791
rect 4580 20760 4629 20788
rect 4580 20748 4586 20760
rect 4617 20757 4629 20760
rect 4663 20757 4675 20791
rect 4617 20751 4675 20757
rect 8202 20748 8208 20800
rect 8260 20788 8266 20800
rect 8757 20791 8815 20797
rect 8757 20788 8769 20791
rect 8260 20760 8769 20788
rect 8260 20748 8266 20760
rect 8757 20757 8769 20760
rect 8803 20788 8815 20791
rect 9306 20788 9312 20800
rect 8803 20760 9312 20788
rect 8803 20757 8815 20760
rect 8757 20751 8815 20757
rect 9306 20748 9312 20760
rect 9364 20748 9370 20800
rect 11054 20748 11060 20800
rect 11112 20788 11118 20800
rect 11425 20791 11483 20797
rect 11425 20788 11437 20791
rect 11112 20760 11437 20788
rect 11112 20748 11118 20760
rect 11425 20757 11437 20760
rect 11471 20757 11483 20791
rect 11425 20751 11483 20757
rect 14001 20791 14059 20797
rect 14001 20757 14013 20791
rect 14047 20788 14059 20791
rect 14090 20788 14096 20800
rect 14047 20760 14096 20788
rect 14047 20757 14059 20760
rect 14001 20751 14059 20757
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 3605 20587 3663 20593
rect 3605 20553 3617 20587
rect 3651 20584 3663 20587
rect 4062 20584 4068 20596
rect 3651 20556 4068 20584
rect 3651 20553 3663 20556
rect 3605 20547 3663 20553
rect 4062 20544 4068 20556
rect 4120 20544 4126 20596
rect 5077 20587 5135 20593
rect 5077 20553 5089 20587
rect 5123 20584 5135 20587
rect 5166 20584 5172 20596
rect 5123 20556 5172 20584
rect 5123 20553 5135 20556
rect 5077 20547 5135 20553
rect 5166 20544 5172 20556
rect 5224 20544 5230 20596
rect 5534 20544 5540 20596
rect 5592 20584 5598 20596
rect 5994 20584 6000 20596
rect 5592 20556 6000 20584
rect 5592 20544 5598 20556
rect 5994 20544 6000 20556
rect 6052 20544 6058 20596
rect 6641 20587 6699 20593
rect 6641 20553 6653 20587
rect 6687 20584 6699 20587
rect 7006 20584 7012 20596
rect 6687 20556 7012 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 7006 20544 7012 20556
rect 7064 20584 7070 20596
rect 8205 20587 8263 20593
rect 8205 20584 8217 20587
rect 7064 20556 8217 20584
rect 7064 20544 7070 20556
rect 8205 20553 8217 20556
rect 8251 20553 8263 20587
rect 9030 20584 9036 20596
rect 8991 20556 9036 20584
rect 8205 20547 8263 20553
rect 9030 20544 9036 20556
rect 9088 20544 9094 20596
rect 10134 20544 10140 20596
rect 10192 20584 10198 20596
rect 10597 20587 10655 20593
rect 10597 20584 10609 20587
rect 10192 20556 10609 20584
rect 10192 20544 10198 20556
rect 10597 20553 10609 20556
rect 10643 20553 10655 20587
rect 11882 20584 11888 20596
rect 11795 20556 11888 20584
rect 10597 20547 10655 20553
rect 11882 20544 11888 20556
rect 11940 20584 11946 20596
rect 12342 20584 12348 20596
rect 11940 20556 12348 20584
rect 11940 20544 11946 20556
rect 12342 20544 12348 20556
rect 12400 20544 12406 20596
rect 13265 20587 13323 20593
rect 13265 20553 13277 20587
rect 13311 20584 13323 20587
rect 13354 20584 13360 20596
rect 13311 20556 13360 20584
rect 13311 20553 13323 20556
rect 13265 20547 13323 20553
rect 13354 20544 13360 20556
rect 13412 20544 13418 20596
rect 15197 20587 15255 20593
rect 15197 20553 15209 20587
rect 15243 20584 15255 20587
rect 15286 20584 15292 20596
rect 15243 20556 15292 20584
rect 15243 20553 15255 20556
rect 15197 20547 15255 20553
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 5258 20476 5264 20528
rect 5316 20516 5322 20528
rect 5721 20519 5779 20525
rect 5721 20516 5733 20519
rect 5316 20488 5733 20516
rect 5316 20476 5322 20488
rect 5721 20485 5733 20488
rect 5767 20516 5779 20519
rect 6454 20516 6460 20528
rect 5767 20488 6460 20516
rect 5767 20485 5779 20488
rect 5721 20479 5779 20485
rect 6454 20476 6460 20488
rect 6512 20476 6518 20528
rect 2314 20448 2320 20460
rect 1504 20420 2320 20448
rect 1504 20389 1532 20420
rect 2314 20408 2320 20420
rect 2372 20408 2378 20460
rect 9048 20448 9076 20544
rect 9048 20420 9444 20448
rect 1489 20383 1547 20389
rect 1489 20349 1501 20383
rect 1535 20349 1547 20383
rect 1762 20380 1768 20392
rect 1723 20352 1768 20380
rect 1489 20343 1547 20349
rect 1762 20340 1768 20352
rect 1820 20340 1826 20392
rect 3697 20383 3755 20389
rect 3697 20349 3709 20383
rect 3743 20380 3755 20383
rect 3786 20380 3792 20392
rect 3743 20352 3792 20380
rect 3743 20349 3755 20352
rect 3697 20343 3755 20349
rect 3786 20340 3792 20352
rect 3844 20340 3850 20392
rect 6730 20340 6736 20392
rect 6788 20380 6794 20392
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 6788 20352 6837 20380
rect 6788 20340 6794 20352
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 9030 20380 9036 20392
rect 6825 20343 6883 20349
rect 7024 20352 9036 20380
rect 3964 20315 4022 20321
rect 3964 20281 3976 20315
rect 4010 20312 4022 20315
rect 4062 20312 4068 20324
rect 4010 20284 4068 20312
rect 4010 20281 4022 20284
rect 3964 20275 4022 20281
rect 4062 20272 4068 20284
rect 4120 20272 4126 20324
rect 6840 20312 6868 20343
rect 7024 20312 7052 20352
rect 9030 20340 9036 20352
rect 9088 20340 9094 20392
rect 7098 20321 7104 20324
rect 6840 20284 7052 20312
rect 7092 20275 7104 20321
rect 7156 20312 7162 20324
rect 8202 20312 8208 20324
rect 7156 20284 8208 20312
rect 7098 20272 7104 20275
rect 7156 20272 7162 20284
rect 8202 20272 8208 20284
rect 8260 20272 8266 20324
rect 9416 20312 9444 20420
rect 9950 20408 9956 20460
rect 10008 20448 10014 20460
rect 10229 20451 10287 20457
rect 10229 20448 10241 20451
rect 10008 20420 10241 20448
rect 10008 20408 10014 20420
rect 10229 20417 10241 20420
rect 10275 20448 10287 20451
rect 10962 20448 10968 20460
rect 10275 20420 10968 20448
rect 10275 20417 10287 20420
rect 10229 20411 10287 20417
rect 10962 20408 10968 20420
rect 11020 20408 11026 20460
rect 11057 20451 11115 20457
rect 11057 20417 11069 20451
rect 11103 20448 11115 20451
rect 11146 20448 11152 20460
rect 11103 20420 11152 20448
rect 11103 20417 11115 20420
rect 11057 20411 11115 20417
rect 11146 20408 11152 20420
rect 11204 20448 11210 20460
rect 12342 20448 12348 20460
rect 11204 20420 12348 20448
rect 11204 20408 11210 20420
rect 12342 20408 12348 20420
rect 12400 20408 12406 20460
rect 13814 20448 13820 20460
rect 13775 20420 13820 20448
rect 13814 20408 13820 20420
rect 13872 20408 13878 20460
rect 9493 20383 9551 20389
rect 9493 20349 9505 20383
rect 9539 20380 9551 20383
rect 10045 20383 10103 20389
rect 10045 20380 10057 20383
rect 9539 20352 10057 20380
rect 9539 20349 9551 20352
rect 9493 20343 9551 20349
rect 10045 20349 10057 20352
rect 10091 20380 10103 20383
rect 10870 20380 10876 20392
rect 10091 20352 10876 20380
rect 10091 20349 10103 20352
rect 10045 20343 10103 20349
rect 10870 20340 10876 20352
rect 10928 20340 10934 20392
rect 12253 20383 12311 20389
rect 12253 20349 12265 20383
rect 12299 20380 12311 20383
rect 12437 20383 12495 20389
rect 12437 20380 12449 20383
rect 12299 20352 12449 20380
rect 12299 20349 12311 20352
rect 12253 20343 12311 20349
rect 12437 20349 12449 20352
rect 12483 20380 12495 20383
rect 12802 20380 12808 20392
rect 12483 20352 12808 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 13354 20340 13360 20392
rect 13412 20380 13418 20392
rect 13832 20380 13860 20408
rect 13412 20352 14228 20380
rect 13412 20340 13418 20352
rect 14200 20324 14228 20352
rect 9953 20315 10011 20321
rect 9953 20312 9965 20315
rect 9416 20284 9965 20312
rect 9953 20281 9965 20284
rect 9999 20312 10011 20315
rect 10686 20312 10692 20324
rect 9999 20284 10692 20312
rect 9999 20281 10011 20284
rect 9953 20275 10011 20281
rect 10686 20272 10692 20284
rect 10744 20272 10750 20324
rect 12710 20312 12716 20324
rect 12671 20284 12716 20312
rect 12710 20272 12716 20284
rect 12768 20272 12774 20324
rect 14090 20321 14096 20324
rect 14084 20312 14096 20321
rect 14051 20284 14096 20312
rect 14084 20275 14096 20284
rect 14090 20272 14096 20275
rect 14148 20272 14154 20324
rect 14182 20272 14188 20324
rect 14240 20272 14246 20324
rect 2682 20244 2688 20256
rect 2643 20216 2688 20244
rect 2682 20204 2688 20216
rect 2740 20204 2746 20256
rect 3050 20244 3056 20256
rect 2963 20216 3056 20244
rect 3050 20204 3056 20216
rect 3108 20244 3114 20256
rect 3510 20244 3516 20256
rect 3108 20216 3516 20244
rect 3108 20204 3114 20216
rect 3510 20204 3516 20216
rect 3568 20204 3574 20256
rect 9582 20244 9588 20256
rect 9543 20216 9588 20244
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 11330 20244 11336 20256
rect 11291 20216 11336 20244
rect 11330 20204 11336 20216
rect 11388 20204 11394 20256
rect 13170 20204 13176 20256
rect 13228 20244 13234 20256
rect 13541 20247 13599 20253
rect 13541 20244 13553 20247
rect 13228 20216 13553 20244
rect 13228 20204 13234 20216
rect 13541 20213 13553 20216
rect 13587 20213 13599 20247
rect 16298 20244 16304 20256
rect 16259 20216 16304 20244
rect 13541 20207 13599 20213
rect 16298 20204 16304 20216
rect 16356 20204 16362 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 6917 20043 6975 20049
rect 6917 20009 6929 20043
rect 6963 20040 6975 20043
rect 7098 20040 7104 20052
rect 6963 20012 7104 20040
rect 6963 20009 6975 20012
rect 6917 20003 6975 20009
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 8481 20043 8539 20049
rect 8481 20009 8493 20043
rect 8527 20040 8539 20043
rect 8754 20040 8760 20052
rect 8527 20012 8760 20040
rect 8527 20009 8539 20012
rect 8481 20003 8539 20009
rect 8754 20000 8760 20012
rect 8812 20040 8818 20052
rect 9582 20040 9588 20052
rect 8812 20012 9588 20040
rect 8812 20000 8818 20012
rect 9582 20000 9588 20012
rect 9640 20000 9646 20052
rect 12986 20040 12992 20052
rect 12947 20012 12992 20040
rect 12986 20000 12992 20012
rect 13044 20000 13050 20052
rect 13173 20043 13231 20049
rect 13173 20009 13185 20043
rect 13219 20040 13231 20043
rect 15749 20043 15807 20049
rect 15749 20040 15761 20043
rect 13219 20012 15761 20040
rect 13219 20009 13231 20012
rect 13173 20003 13231 20009
rect 15749 20009 15761 20012
rect 15795 20040 15807 20043
rect 16022 20040 16028 20052
rect 15795 20012 16028 20040
rect 15795 20009 15807 20012
rect 15749 20003 15807 20009
rect 16022 20000 16028 20012
rect 16080 20000 16086 20052
rect 1765 19975 1823 19981
rect 1765 19941 1777 19975
rect 1811 19972 1823 19975
rect 2222 19972 2228 19984
rect 1811 19944 2228 19972
rect 1811 19941 1823 19944
rect 1765 19935 1823 19941
rect 2222 19932 2228 19944
rect 2280 19932 2286 19984
rect 4617 19975 4675 19981
rect 4617 19941 4629 19975
rect 4663 19972 4675 19975
rect 4976 19975 5034 19981
rect 4976 19972 4988 19975
rect 4663 19944 4988 19972
rect 4663 19941 4675 19944
rect 4617 19935 4675 19941
rect 4976 19941 4988 19944
rect 5022 19972 5034 19975
rect 5166 19972 5172 19984
rect 5022 19944 5172 19972
rect 5022 19941 5034 19944
rect 4976 19935 5034 19941
rect 5166 19932 5172 19944
rect 5224 19932 5230 19984
rect 9030 19972 9036 19984
rect 8991 19944 9036 19972
rect 9030 19932 9036 19944
rect 9088 19932 9094 19984
rect 9950 19972 9956 19984
rect 9911 19944 9956 19972
rect 9950 19932 9956 19944
rect 10008 19972 10014 19984
rect 10290 19975 10348 19981
rect 10290 19972 10302 19975
rect 10008 19944 10302 19972
rect 10008 19932 10014 19944
rect 10290 19941 10302 19944
rect 10336 19941 10348 19975
rect 10290 19935 10348 19941
rect 13633 19975 13691 19981
rect 13633 19941 13645 19975
rect 13679 19972 13691 19975
rect 13722 19972 13728 19984
rect 13679 19944 13728 19972
rect 13679 19941 13691 19944
rect 13633 19935 13691 19941
rect 13722 19932 13728 19944
rect 13780 19932 13786 19984
rect 14182 19972 14188 19984
rect 14143 19944 14188 19972
rect 14182 19932 14188 19944
rect 14240 19932 14246 19984
rect 15654 19972 15660 19984
rect 15615 19944 15660 19972
rect 15654 19932 15660 19944
rect 15712 19932 15718 19984
rect 1489 19907 1547 19913
rect 1489 19873 1501 19907
rect 1535 19904 1547 19907
rect 2777 19907 2835 19913
rect 1535 19876 2360 19904
rect 1535 19873 1547 19876
rect 1489 19867 1547 19873
rect 2332 19848 2360 19876
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 3418 19904 3424 19916
rect 2823 19876 3424 19904
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 3418 19864 3424 19876
rect 3476 19864 3482 19916
rect 3970 19864 3976 19916
rect 4028 19904 4034 19916
rect 4430 19904 4436 19916
rect 4028 19876 4436 19904
rect 4028 19864 4034 19876
rect 4430 19864 4436 19876
rect 4488 19904 4494 19916
rect 4709 19907 4767 19913
rect 4709 19904 4721 19907
rect 4488 19876 4721 19904
rect 4488 19864 4494 19876
rect 4709 19873 4721 19876
rect 4755 19904 4767 19907
rect 5442 19904 5448 19916
rect 4755 19876 5448 19904
rect 4755 19873 4767 19876
rect 4709 19867 4767 19873
rect 5442 19864 5448 19876
rect 5500 19904 5506 19916
rect 5500 19876 6592 19904
rect 5500 19864 5506 19876
rect 2314 19836 2320 19848
rect 2275 19808 2320 19836
rect 2314 19796 2320 19808
rect 2372 19796 2378 19848
rect 6564 19836 6592 19876
rect 7006 19864 7012 19916
rect 7064 19904 7070 19916
rect 7561 19907 7619 19913
rect 7561 19904 7573 19907
rect 7064 19876 7573 19904
rect 7064 19864 7070 19876
rect 7561 19873 7573 19876
rect 7607 19873 7619 19907
rect 8386 19904 8392 19916
rect 8347 19876 8392 19904
rect 7561 19867 7619 19873
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 9493 19907 9551 19913
rect 9493 19873 9505 19907
rect 9539 19904 9551 19907
rect 10042 19904 10048 19916
rect 9539 19876 10048 19904
rect 9539 19873 9551 19876
rect 9493 19867 9551 19873
rect 10042 19864 10048 19876
rect 10100 19904 10106 19916
rect 11146 19904 11152 19916
rect 10100 19876 11152 19904
rect 10100 19864 10106 19876
rect 11146 19864 11152 19876
rect 11204 19864 11210 19916
rect 12802 19864 12808 19916
rect 12860 19904 12866 19916
rect 13538 19904 13544 19916
rect 12860 19876 13544 19904
rect 12860 19864 12866 19876
rect 13538 19864 13544 19876
rect 13596 19864 13602 19916
rect 7837 19839 7895 19845
rect 7837 19836 7849 19839
rect 6564 19808 7849 19836
rect 7837 19805 7849 19808
rect 7883 19836 7895 19839
rect 7926 19836 7932 19848
rect 7883 19808 7932 19836
rect 7883 19805 7895 19808
rect 7837 19799 7895 19805
rect 7926 19796 7932 19808
rect 7984 19796 7990 19848
rect 8662 19836 8668 19848
rect 8575 19808 8668 19836
rect 8662 19796 8668 19808
rect 8720 19836 8726 19848
rect 13817 19839 13875 19845
rect 8720 19808 9536 19836
rect 8720 19796 8726 19808
rect 8018 19768 8024 19780
rect 7979 19740 8024 19768
rect 8018 19728 8024 19740
rect 8076 19728 8082 19780
rect 2498 19660 2504 19712
rect 2556 19700 2562 19712
rect 2593 19703 2651 19709
rect 2593 19700 2605 19703
rect 2556 19672 2605 19700
rect 2556 19660 2562 19672
rect 2593 19669 2605 19672
rect 2639 19669 2651 19703
rect 2593 19663 2651 19669
rect 2961 19703 3019 19709
rect 2961 19669 2973 19703
rect 3007 19700 3019 19703
rect 3050 19700 3056 19712
rect 3007 19672 3056 19700
rect 3007 19669 3019 19672
rect 2961 19663 3019 19669
rect 3050 19660 3056 19672
rect 3108 19660 3114 19712
rect 3418 19700 3424 19712
rect 3379 19672 3424 19700
rect 3418 19660 3424 19672
rect 3476 19660 3482 19712
rect 3789 19703 3847 19709
rect 3789 19669 3801 19703
rect 3835 19700 3847 19703
rect 3970 19700 3976 19712
rect 3835 19672 3976 19700
rect 3835 19669 3847 19672
rect 3789 19663 3847 19669
rect 3970 19660 3976 19672
rect 4028 19660 4034 19712
rect 6089 19703 6147 19709
rect 6089 19669 6101 19703
rect 6135 19700 6147 19703
rect 6178 19700 6184 19712
rect 6135 19672 6184 19700
rect 6135 19669 6147 19672
rect 6089 19663 6147 19669
rect 6178 19660 6184 19672
rect 6236 19660 6242 19712
rect 6914 19660 6920 19712
rect 6972 19700 6978 19712
rect 7285 19703 7343 19709
rect 7285 19700 7297 19703
rect 6972 19672 7297 19700
rect 6972 19660 6978 19672
rect 7285 19669 7297 19672
rect 7331 19700 7343 19703
rect 7374 19700 7380 19712
rect 7331 19672 7380 19700
rect 7331 19669 7343 19672
rect 7285 19663 7343 19669
rect 7374 19660 7380 19672
rect 7432 19660 7438 19712
rect 9508 19700 9536 19808
rect 13817 19805 13829 19839
rect 13863 19836 13875 19839
rect 14090 19836 14096 19848
rect 13863 19808 14096 19836
rect 13863 19805 13875 19808
rect 13817 19799 13875 19805
rect 12621 19771 12679 19777
rect 12621 19737 12633 19771
rect 12667 19768 12679 19771
rect 13832 19768 13860 19799
rect 14090 19796 14096 19808
rect 14148 19836 14154 19848
rect 14642 19836 14648 19848
rect 14148 19808 14648 19836
rect 14148 19796 14154 19808
rect 14642 19796 14648 19808
rect 14700 19796 14706 19848
rect 15286 19796 15292 19848
rect 15344 19836 15350 19848
rect 15841 19839 15899 19845
rect 15841 19836 15853 19839
rect 15344 19808 15853 19836
rect 15344 19796 15350 19808
rect 15841 19805 15853 19808
rect 15887 19836 15899 19839
rect 16298 19836 16304 19848
rect 15887 19808 16304 19836
rect 15887 19805 15899 19808
rect 15841 19799 15899 19805
rect 16298 19796 16304 19808
rect 16356 19796 16362 19848
rect 12667 19740 13860 19768
rect 12667 19737 12679 19740
rect 12621 19731 12679 19737
rect 11425 19703 11483 19709
rect 11425 19700 11437 19703
rect 9508 19672 11437 19700
rect 11425 19669 11437 19672
rect 11471 19669 11483 19703
rect 15286 19700 15292 19712
rect 15247 19672 15292 19700
rect 11425 19663 11483 19669
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 4062 19496 4068 19508
rect 4023 19468 4068 19496
rect 4062 19456 4068 19468
rect 4120 19456 4126 19508
rect 5166 19496 5172 19508
rect 5127 19468 5172 19496
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 5442 19496 5448 19508
rect 5403 19468 5448 19496
rect 5442 19456 5448 19468
rect 5500 19456 5506 19508
rect 9306 19496 9312 19508
rect 9267 19468 9312 19496
rect 9306 19456 9312 19468
rect 9364 19456 9370 19508
rect 9950 19456 9956 19508
rect 10008 19496 10014 19508
rect 10045 19499 10103 19505
rect 10045 19496 10057 19499
rect 10008 19468 10057 19496
rect 10008 19456 10014 19468
rect 10045 19465 10057 19468
rect 10091 19465 10103 19499
rect 10045 19459 10103 19465
rect 10781 19499 10839 19505
rect 10781 19465 10793 19499
rect 10827 19496 10839 19499
rect 11606 19496 11612 19508
rect 10827 19468 11612 19496
rect 10827 19465 10839 19468
rect 10781 19459 10839 19465
rect 11606 19456 11612 19468
rect 11664 19496 11670 19508
rect 11882 19496 11888 19508
rect 11664 19468 11888 19496
rect 11664 19456 11670 19468
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 12802 19496 12808 19508
rect 12763 19468 12808 19496
rect 12802 19456 12808 19468
rect 12860 19456 12866 19508
rect 13173 19499 13231 19505
rect 13173 19465 13185 19499
rect 13219 19496 13231 19499
rect 13630 19496 13636 19508
rect 13219 19468 13636 19496
rect 13219 19465 13231 19468
rect 13173 19459 13231 19465
rect 13630 19456 13636 19468
rect 13688 19456 13694 19508
rect 14642 19496 14648 19508
rect 14603 19468 14648 19496
rect 14642 19456 14648 19468
rect 14700 19456 14706 19508
rect 15381 19499 15439 19505
rect 15381 19465 15393 19499
rect 15427 19496 15439 19499
rect 15654 19496 15660 19508
rect 15427 19468 15660 19496
rect 15427 19465 15439 19468
rect 15381 19459 15439 19465
rect 15654 19456 15660 19468
rect 15712 19456 15718 19508
rect 16298 19496 16304 19508
rect 16259 19468 16304 19496
rect 16298 19456 16304 19468
rect 16356 19456 16362 19508
rect 2590 19360 2596 19372
rect 2551 19332 2596 19360
rect 2590 19320 2596 19332
rect 2648 19320 2654 19372
rect 3973 19363 4031 19369
rect 3973 19329 3985 19363
rect 4019 19360 4031 19363
rect 4709 19363 4767 19369
rect 4709 19360 4721 19363
rect 4019 19332 4721 19360
rect 4019 19329 4031 19332
rect 3973 19323 4031 19329
rect 4709 19329 4721 19332
rect 4755 19360 4767 19363
rect 6086 19360 6092 19372
rect 4755 19332 6092 19360
rect 4755 19329 4767 19332
rect 4709 19323 4767 19329
rect 6086 19320 6092 19332
rect 6144 19320 6150 19372
rect 7926 19360 7932 19372
rect 7887 19332 7932 19360
rect 7926 19320 7932 19332
rect 7984 19320 7990 19372
rect 3237 19295 3295 19301
rect 3237 19261 3249 19295
rect 3283 19292 3295 19295
rect 4522 19292 4528 19304
rect 3283 19264 4528 19292
rect 3283 19261 3295 19264
rect 3237 19255 3295 19261
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 5629 19295 5687 19301
rect 5629 19261 5641 19295
rect 5675 19261 5687 19295
rect 5629 19255 5687 19261
rect 7469 19295 7527 19301
rect 7469 19261 7481 19295
rect 7515 19292 7527 19295
rect 8196 19295 8254 19301
rect 8196 19292 8208 19295
rect 7515 19264 8208 19292
rect 7515 19261 7527 19264
rect 7469 19255 7527 19261
rect 8196 19261 8208 19264
rect 8242 19292 8254 19295
rect 8662 19292 8668 19304
rect 8242 19264 8668 19292
rect 8242 19261 8254 19264
rect 8196 19255 8254 19261
rect 1394 19184 1400 19236
rect 1452 19224 1458 19236
rect 1949 19227 2007 19233
rect 1949 19224 1961 19227
rect 1452 19196 1961 19224
rect 1452 19184 1458 19196
rect 1949 19193 1961 19196
rect 1995 19224 2007 19227
rect 2409 19227 2467 19233
rect 2409 19224 2421 19227
rect 1995 19196 2421 19224
rect 1995 19193 2007 19196
rect 1949 19187 2007 19193
rect 2409 19193 2421 19196
rect 2455 19193 2467 19227
rect 2409 19187 2467 19193
rect 2958 19184 2964 19236
rect 3016 19224 3022 19236
rect 5644 19224 5672 19255
rect 8662 19252 8668 19264
rect 8720 19252 8726 19304
rect 10965 19295 11023 19301
rect 10965 19292 10977 19295
rect 10612 19264 10977 19292
rect 6270 19224 6276 19236
rect 3016 19196 5580 19224
rect 5644 19196 6276 19224
rect 3016 19184 3022 19196
rect 2038 19156 2044 19168
rect 1999 19128 2044 19156
rect 2038 19116 2044 19128
rect 2096 19116 2102 19168
rect 2498 19156 2504 19168
rect 2459 19128 2504 19156
rect 2498 19116 2504 19128
rect 2556 19116 2562 19168
rect 3605 19159 3663 19165
rect 3605 19125 3617 19159
rect 3651 19156 3663 19159
rect 3786 19156 3792 19168
rect 3651 19128 3792 19156
rect 3651 19125 3663 19128
rect 3605 19119 3663 19125
rect 3786 19116 3792 19128
rect 3844 19116 3850 19168
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4433 19159 4491 19165
rect 4433 19156 4445 19159
rect 4212 19128 4445 19156
rect 4212 19116 4218 19128
rect 4433 19125 4445 19128
rect 4479 19125 4491 19159
rect 5552 19156 5580 19196
rect 6270 19184 6276 19196
rect 6328 19184 6334 19236
rect 5813 19159 5871 19165
rect 5813 19156 5825 19159
rect 5552 19128 5825 19156
rect 4433 19119 4491 19125
rect 5813 19125 5825 19128
rect 5859 19125 5871 19159
rect 6638 19156 6644 19168
rect 6599 19128 6644 19156
rect 5813 19119 5871 19125
rect 6638 19116 6644 19128
rect 6696 19116 6702 19168
rect 6822 19156 6828 19168
rect 6783 19128 6828 19156
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 7837 19159 7895 19165
rect 7837 19125 7849 19159
rect 7883 19156 7895 19159
rect 8202 19156 8208 19168
rect 7883 19128 8208 19156
rect 7883 19125 7895 19128
rect 7837 19119 7895 19125
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 10612 19165 10640 19264
rect 10965 19261 10977 19264
rect 11011 19261 11023 19295
rect 10965 19255 11023 19261
rect 11057 19295 11115 19301
rect 11057 19261 11069 19295
rect 11103 19292 11115 19295
rect 11882 19292 11888 19304
rect 11103 19264 11888 19292
rect 11103 19261 11115 19264
rect 11057 19255 11115 19261
rect 11882 19252 11888 19264
rect 11940 19252 11946 19304
rect 13265 19295 13323 19301
rect 13265 19261 13277 19295
rect 13311 19292 13323 19295
rect 13354 19292 13360 19304
rect 13311 19264 13360 19292
rect 13311 19261 13323 19264
rect 13265 19255 13323 19261
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 15562 19252 15568 19304
rect 15620 19292 15626 19304
rect 15749 19295 15807 19301
rect 15749 19292 15761 19295
rect 15620 19264 15761 19292
rect 15620 19252 15626 19264
rect 15749 19261 15761 19264
rect 15795 19292 15807 19295
rect 16669 19295 16727 19301
rect 16669 19292 16681 19295
rect 15795 19264 16681 19292
rect 15795 19261 15807 19264
rect 15749 19255 15807 19261
rect 16669 19261 16681 19264
rect 16715 19261 16727 19295
rect 16669 19255 16727 19261
rect 11146 19184 11152 19236
rect 11204 19224 11210 19236
rect 11333 19227 11391 19233
rect 11333 19224 11345 19227
rect 11204 19196 11345 19224
rect 11204 19184 11210 19196
rect 11333 19193 11345 19196
rect 11379 19193 11391 19227
rect 11333 19187 11391 19193
rect 11974 19184 11980 19236
rect 12032 19224 12038 19236
rect 12253 19227 12311 19233
rect 12253 19224 12265 19227
rect 12032 19196 12265 19224
rect 12032 19184 12038 19196
rect 12253 19193 12265 19196
rect 12299 19224 12311 19227
rect 13510 19227 13568 19233
rect 13510 19224 13522 19227
rect 12299 19196 13522 19224
rect 12299 19193 12311 19196
rect 12253 19187 12311 19193
rect 13510 19193 13522 19196
rect 13556 19224 13568 19227
rect 13906 19224 13912 19236
rect 13556 19196 13912 19224
rect 13556 19193 13568 19196
rect 13510 19187 13568 19193
rect 13906 19184 13912 19196
rect 13964 19184 13970 19236
rect 10597 19159 10655 19165
rect 10597 19156 10609 19159
rect 10192 19128 10609 19156
rect 10192 19116 10198 19128
rect 10597 19125 10609 19128
rect 10643 19125 10655 19159
rect 15930 19156 15936 19168
rect 15891 19128 15936 19156
rect 10597 19119 10655 19125
rect 15930 19116 15936 19128
rect 15988 19116 15994 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1394 18952 1400 18964
rect 1355 18924 1400 18952
rect 1394 18912 1400 18924
rect 1452 18912 1458 18964
rect 4430 18952 4436 18964
rect 4391 18924 4436 18952
rect 4430 18912 4436 18924
rect 4488 18952 4494 18964
rect 4706 18952 4712 18964
rect 4488 18924 4712 18952
rect 4488 18912 4494 18924
rect 4706 18912 4712 18924
rect 4764 18912 4770 18964
rect 5534 18952 5540 18964
rect 5495 18924 5540 18952
rect 5534 18912 5540 18924
rect 5592 18952 5598 18964
rect 6086 18952 6092 18964
rect 5592 18924 6092 18952
rect 5592 18912 5598 18924
rect 6086 18912 6092 18924
rect 6144 18912 6150 18964
rect 8754 18952 8760 18964
rect 8715 18924 8760 18952
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 13906 18952 13912 18964
rect 13867 18924 13912 18952
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 16022 18952 16028 18964
rect 15983 18924 16028 18952
rect 16022 18912 16028 18924
rect 16080 18912 16086 18964
rect 4246 18844 4252 18896
rect 4304 18884 4310 18896
rect 5077 18887 5135 18893
rect 5077 18884 5089 18887
rect 4304 18856 5089 18884
rect 4304 18844 4310 18856
rect 5077 18853 5089 18856
rect 5123 18884 5135 18887
rect 5258 18884 5264 18896
rect 5123 18856 5264 18884
rect 5123 18853 5135 18856
rect 5077 18847 5135 18853
rect 5258 18844 5264 18856
rect 5316 18844 5322 18896
rect 5994 18844 6000 18896
rect 6052 18884 6058 18896
rect 6181 18887 6239 18893
rect 6181 18884 6193 18887
rect 6052 18856 6193 18884
rect 6052 18844 6058 18856
rect 6181 18853 6193 18856
rect 6227 18853 6239 18887
rect 6181 18847 6239 18853
rect 8389 18887 8447 18893
rect 8389 18853 8401 18887
rect 8435 18884 8447 18887
rect 8662 18884 8668 18896
rect 8435 18856 8668 18884
rect 8435 18853 8447 18856
rect 8389 18847 8447 18853
rect 8662 18844 8668 18856
rect 8720 18844 8726 18896
rect 12526 18844 12532 18896
rect 12584 18884 12590 18896
rect 12774 18887 12832 18893
rect 12774 18884 12786 18887
rect 12584 18856 12786 18884
rect 12584 18844 12590 18856
rect 12774 18853 12786 18856
rect 12820 18853 12832 18887
rect 15562 18884 15568 18896
rect 15523 18856 15568 18884
rect 12774 18847 12832 18853
rect 15562 18844 15568 18856
rect 15620 18844 15626 18896
rect 2774 18816 2780 18828
rect 2735 18788 2780 18816
rect 2774 18776 2780 18788
rect 2832 18776 2838 18828
rect 3421 18819 3479 18825
rect 3421 18816 3433 18819
rect 2884 18788 3433 18816
rect 2884 18760 2912 18788
rect 3421 18785 3433 18788
rect 3467 18785 3479 18819
rect 4525 18819 4583 18825
rect 4525 18816 4537 18819
rect 3421 18779 3479 18785
rect 3804 18788 4537 18816
rect 2866 18748 2872 18760
rect 2827 18720 2872 18748
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 2958 18708 2964 18760
rect 3016 18748 3022 18760
rect 3016 18720 3061 18748
rect 3016 18708 3022 18720
rect 3804 18689 3832 18788
rect 4525 18785 4537 18788
rect 4571 18785 4583 18819
rect 7650 18816 7656 18828
rect 7611 18788 7656 18816
rect 4525 18779 4583 18785
rect 7650 18776 7656 18788
rect 7708 18776 7714 18828
rect 7745 18819 7803 18825
rect 7745 18785 7757 18819
rect 7791 18816 7803 18819
rect 7926 18816 7932 18828
rect 7791 18788 7932 18816
rect 7791 18785 7803 18788
rect 7745 18779 7803 18785
rect 7926 18776 7932 18788
rect 7984 18776 7990 18828
rect 9677 18819 9735 18825
rect 9677 18785 9689 18819
rect 9723 18816 9735 18819
rect 11330 18816 11336 18828
rect 9723 18788 10548 18816
rect 11291 18788 11336 18816
rect 9723 18785 9735 18788
rect 9677 18779 9735 18785
rect 4614 18748 4620 18760
rect 4575 18720 4620 18748
rect 4614 18708 4620 18720
rect 4672 18708 4678 18760
rect 6362 18748 6368 18760
rect 6323 18720 6368 18748
rect 6362 18708 6368 18720
rect 6420 18708 6426 18760
rect 7837 18751 7895 18757
rect 7837 18717 7849 18751
rect 7883 18748 7895 18751
rect 8202 18748 8208 18760
rect 7883 18720 8208 18748
rect 7883 18717 7895 18720
rect 7837 18711 7895 18717
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 9858 18748 9864 18760
rect 9819 18720 9864 18748
rect 9858 18708 9864 18720
rect 9916 18708 9922 18760
rect 2409 18683 2467 18689
rect 2409 18649 2421 18683
rect 2455 18680 2467 18683
rect 3789 18683 3847 18689
rect 3789 18680 3801 18683
rect 2455 18652 3801 18680
rect 2455 18649 2467 18652
rect 2409 18643 2467 18649
rect 3789 18649 3801 18652
rect 3835 18649 3847 18683
rect 4062 18680 4068 18692
rect 4023 18652 4068 18680
rect 3789 18643 3847 18649
rect 4062 18640 4068 18652
rect 4120 18640 4126 18692
rect 5626 18640 5632 18692
rect 5684 18680 5690 18692
rect 5721 18683 5779 18689
rect 5721 18680 5733 18683
rect 5684 18652 5733 18680
rect 5684 18640 5690 18652
rect 5721 18649 5733 18652
rect 5767 18649 5779 18683
rect 7282 18680 7288 18692
rect 7243 18652 7288 18680
rect 5721 18643 5779 18649
rect 7282 18640 7288 18652
rect 7340 18640 7346 18692
rect 10520 18689 10548 18788
rect 11330 18776 11336 18788
rect 11388 18776 11394 18828
rect 15286 18816 15292 18828
rect 15247 18788 15292 18816
rect 15286 18776 15292 18788
rect 15344 18776 15350 18828
rect 11422 18748 11428 18760
rect 11383 18720 11428 18748
rect 11422 18708 11428 18720
rect 11480 18708 11486 18760
rect 11609 18751 11667 18757
rect 11609 18717 11621 18751
rect 11655 18748 11667 18751
rect 11974 18748 11980 18760
rect 11655 18720 11980 18748
rect 11655 18717 11667 18720
rect 11609 18711 11667 18717
rect 11974 18708 11980 18720
rect 12032 18708 12038 18760
rect 12529 18751 12587 18757
rect 12529 18748 12541 18751
rect 12176 18720 12541 18748
rect 10505 18683 10563 18689
rect 10505 18649 10517 18683
rect 10551 18680 10563 18683
rect 10965 18683 11023 18689
rect 10965 18680 10977 18683
rect 10551 18652 10977 18680
rect 10551 18649 10563 18652
rect 10505 18643 10563 18649
rect 10965 18649 10977 18652
rect 11011 18649 11023 18683
rect 10965 18643 11023 18649
rect 12176 18624 12204 18720
rect 12529 18717 12541 18720
rect 12575 18717 12587 18751
rect 12529 18711 12587 18717
rect 2038 18572 2044 18624
rect 2096 18612 2102 18624
rect 2133 18615 2191 18621
rect 2133 18612 2145 18615
rect 2096 18584 2145 18612
rect 2096 18572 2102 18584
rect 2133 18581 2145 18584
rect 2179 18612 2191 18615
rect 2590 18612 2596 18624
rect 2179 18584 2596 18612
rect 2179 18581 2191 18584
rect 2133 18575 2191 18581
rect 2590 18572 2596 18584
rect 2648 18612 2654 18624
rect 2958 18612 2964 18624
rect 2648 18584 2964 18612
rect 2648 18572 2654 18584
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 6917 18615 6975 18621
rect 6917 18581 6929 18615
rect 6963 18612 6975 18615
rect 7190 18612 7196 18624
rect 6963 18584 7196 18612
rect 6963 18581 6975 18584
rect 6917 18575 6975 18581
rect 7190 18572 7196 18584
rect 7248 18572 7254 18624
rect 9306 18612 9312 18624
rect 9267 18584 9312 18612
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 10870 18612 10876 18624
rect 10831 18584 10876 18612
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 12069 18615 12127 18621
rect 12069 18581 12081 18615
rect 12115 18612 12127 18615
rect 12158 18612 12164 18624
rect 12115 18584 12164 18612
rect 12115 18581 12127 18584
rect 12069 18575 12127 18581
rect 12158 18572 12164 18584
rect 12216 18572 12222 18624
rect 12437 18615 12495 18621
rect 12437 18581 12449 18615
rect 12483 18612 12495 18615
rect 12526 18612 12532 18624
rect 12483 18584 12532 18612
rect 12483 18581 12495 18584
rect 12437 18575 12495 18581
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 5994 18368 6000 18420
rect 6052 18408 6058 18420
rect 6181 18411 6239 18417
rect 6181 18408 6193 18411
rect 6052 18380 6193 18408
rect 6052 18368 6058 18380
rect 6181 18377 6193 18380
rect 6227 18408 6239 18411
rect 6546 18408 6552 18420
rect 6227 18380 6552 18408
rect 6227 18377 6239 18380
rect 6181 18371 6239 18377
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 10686 18408 10692 18420
rect 10647 18380 10692 18408
rect 10686 18368 10692 18380
rect 10744 18368 10750 18420
rect 10781 18411 10839 18417
rect 10781 18377 10793 18411
rect 10827 18408 10839 18411
rect 11330 18408 11336 18420
rect 10827 18380 11336 18408
rect 10827 18377 10839 18380
rect 10781 18371 10839 18377
rect 11330 18368 11336 18380
rect 11388 18368 11394 18420
rect 11885 18411 11943 18417
rect 11885 18377 11897 18411
rect 11931 18408 11943 18411
rect 11974 18408 11980 18420
rect 11931 18380 11980 18408
rect 11931 18377 11943 18380
rect 11885 18371 11943 18377
rect 11974 18368 11980 18380
rect 12032 18368 12038 18420
rect 15286 18408 15292 18420
rect 15247 18380 15292 18408
rect 15286 18368 15292 18380
rect 15344 18368 15350 18420
rect 15378 18368 15384 18420
rect 15436 18408 15442 18420
rect 16117 18411 16175 18417
rect 16117 18408 16129 18411
rect 15436 18380 16129 18408
rect 15436 18368 15442 18380
rect 16117 18377 16129 18380
rect 16163 18377 16175 18411
rect 16117 18371 16175 18377
rect 5629 18343 5687 18349
rect 5629 18309 5641 18343
rect 5675 18309 5687 18343
rect 5629 18303 5687 18309
rect 10321 18343 10379 18349
rect 10321 18309 10333 18343
rect 10367 18340 10379 18343
rect 10367 18312 11468 18340
rect 10367 18309 10379 18312
rect 10321 18303 10379 18309
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 5644 18272 5672 18303
rect 6362 18272 6368 18284
rect 1719 18244 1900 18272
rect 5644 18244 6368 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 1872 18204 1900 18244
rect 6362 18232 6368 18244
rect 6420 18272 6426 18284
rect 7469 18275 7527 18281
rect 7469 18272 7481 18275
rect 6420 18244 7481 18272
rect 6420 18232 6426 18244
rect 7469 18241 7481 18244
rect 7515 18272 7527 18275
rect 8205 18275 8263 18281
rect 8205 18272 8217 18275
rect 7515 18244 8217 18272
rect 7515 18241 7527 18244
rect 7469 18235 7527 18241
rect 8205 18241 8217 18244
rect 8251 18241 8263 18275
rect 8205 18235 8263 18241
rect 9306 18232 9312 18284
rect 9364 18272 9370 18284
rect 9674 18272 9680 18284
rect 9364 18244 9680 18272
rect 9364 18232 9370 18244
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 9861 18275 9919 18281
rect 9861 18241 9873 18275
rect 9907 18272 9919 18275
rect 11054 18272 11060 18284
rect 9907 18244 11060 18272
rect 9907 18241 9919 18244
rect 9861 18235 9919 18241
rect 2038 18213 2044 18216
rect 2032 18204 2044 18213
rect 1872 18176 2044 18204
rect 2032 18167 2044 18176
rect 2038 18164 2044 18167
rect 2096 18164 2102 18216
rect 4249 18207 4307 18213
rect 4249 18173 4261 18207
rect 4295 18204 4307 18207
rect 4338 18204 4344 18216
rect 4295 18176 4344 18204
rect 4295 18173 4307 18176
rect 4249 18167 4307 18173
rect 4338 18164 4344 18176
rect 4396 18204 4402 18216
rect 5626 18204 5632 18216
rect 4396 18176 5632 18204
rect 4396 18164 4402 18176
rect 5626 18164 5632 18176
rect 5684 18164 5690 18216
rect 7285 18207 7343 18213
rect 7285 18204 7297 18207
rect 6564 18176 7297 18204
rect 3789 18139 3847 18145
rect 3789 18105 3801 18139
rect 3835 18136 3847 18139
rect 4157 18139 4215 18145
rect 4157 18136 4169 18139
rect 3835 18108 4169 18136
rect 3835 18105 3847 18108
rect 3789 18099 3847 18105
rect 4157 18105 4169 18108
rect 4203 18136 4215 18139
rect 4516 18139 4574 18145
rect 4516 18136 4528 18139
rect 4203 18108 4528 18136
rect 4203 18105 4215 18108
rect 4157 18099 4215 18105
rect 4516 18105 4528 18108
rect 4562 18136 4574 18139
rect 4614 18136 4620 18148
rect 4562 18108 4620 18136
rect 4562 18105 4574 18108
rect 4516 18099 4574 18105
rect 3145 18071 3203 18077
rect 3145 18037 3157 18071
rect 3191 18068 3203 18071
rect 3804 18068 3832 18099
rect 4614 18096 4620 18108
rect 4672 18096 4678 18148
rect 5074 18096 5080 18148
rect 5132 18136 5138 18148
rect 6564 18145 6592 18176
rect 7285 18173 7297 18176
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 9125 18207 9183 18213
rect 9125 18173 9137 18207
rect 9171 18204 9183 18207
rect 9876 18204 9904 18235
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 11440 18281 11468 18312
rect 11425 18275 11483 18281
rect 11425 18241 11437 18275
rect 11471 18272 11483 18275
rect 15657 18275 15715 18281
rect 11471 18244 12572 18272
rect 11471 18241 11483 18244
rect 11425 18235 11483 18241
rect 12544 18216 12572 18244
rect 15657 18241 15669 18275
rect 15703 18272 15715 18275
rect 16114 18272 16120 18284
rect 15703 18244 16120 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 9171 18176 9904 18204
rect 9171 18173 9183 18176
rect 9125 18167 9183 18173
rect 10870 18164 10876 18216
rect 10928 18204 10934 18216
rect 11149 18207 11207 18213
rect 11149 18204 11161 18207
rect 10928 18176 11161 18204
rect 10928 18164 10934 18176
rect 11149 18173 11161 18176
rect 11195 18204 11207 18207
rect 11238 18204 11244 18216
rect 11195 18176 11244 18204
rect 11195 18173 11207 18176
rect 11149 18167 11207 18173
rect 11238 18164 11244 18176
rect 11296 18164 11302 18216
rect 12158 18164 12164 18216
rect 12216 18204 12222 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 12216 18176 12449 18204
rect 12216 18164 12222 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 12526 18164 12532 18216
rect 12584 18204 12590 18216
rect 12584 18176 13676 18204
rect 12584 18164 12590 18176
rect 6549 18139 6607 18145
rect 6549 18136 6561 18139
rect 5132 18108 6561 18136
rect 5132 18096 5138 18108
rect 6549 18105 6561 18108
rect 6595 18105 6607 18139
rect 6549 18099 6607 18105
rect 6638 18096 6644 18148
rect 6696 18136 6702 18148
rect 7190 18136 7196 18148
rect 6696 18108 7196 18136
rect 6696 18096 6702 18108
rect 7190 18096 7196 18108
rect 7248 18096 7254 18148
rect 8757 18139 8815 18145
rect 8757 18105 8769 18139
rect 8803 18136 8815 18139
rect 9398 18136 9404 18148
rect 8803 18108 9404 18136
rect 8803 18105 8815 18108
rect 8757 18099 8815 18105
rect 9398 18096 9404 18108
rect 9456 18136 9462 18148
rect 9585 18139 9643 18145
rect 9585 18136 9597 18139
rect 9456 18108 9597 18136
rect 9456 18096 9462 18108
rect 9585 18105 9597 18108
rect 9631 18105 9643 18139
rect 9585 18099 9643 18105
rect 12253 18139 12311 18145
rect 12253 18105 12265 18139
rect 12299 18136 12311 18139
rect 12682 18139 12740 18145
rect 12682 18136 12694 18139
rect 12299 18108 12694 18136
rect 12299 18105 12311 18108
rect 12253 18099 12311 18105
rect 12682 18105 12694 18108
rect 12728 18136 12740 18139
rect 13538 18136 13544 18148
rect 12728 18108 13544 18136
rect 12728 18105 12740 18108
rect 12682 18099 12740 18105
rect 13538 18096 13544 18108
rect 13596 18096 13602 18148
rect 3191 18040 3832 18068
rect 3191 18037 3203 18040
rect 3145 18031 3203 18037
rect 6730 18028 6736 18080
rect 6788 18068 6794 18080
rect 6825 18071 6883 18077
rect 6825 18068 6837 18071
rect 6788 18040 6837 18068
rect 6788 18028 6794 18040
rect 6825 18037 6837 18040
rect 6871 18037 6883 18071
rect 6825 18031 6883 18037
rect 7929 18071 7987 18077
rect 7929 18037 7941 18071
rect 7975 18068 7987 18071
rect 8202 18068 8208 18080
rect 7975 18040 8208 18068
rect 7975 18037 7987 18040
rect 7929 18031 7987 18037
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 9214 18068 9220 18080
rect 9175 18040 9220 18068
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 10686 18028 10692 18080
rect 10744 18068 10750 18080
rect 11241 18071 11299 18077
rect 11241 18068 11253 18071
rect 10744 18040 11253 18068
rect 10744 18028 10750 18040
rect 11241 18037 11253 18040
rect 11287 18068 11299 18071
rect 11514 18068 11520 18080
rect 11287 18040 11520 18068
rect 11287 18037 11299 18040
rect 11241 18031 11299 18037
rect 11514 18028 11520 18040
rect 11572 18028 11578 18080
rect 13648 18068 13676 18176
rect 15286 18164 15292 18216
rect 15344 18204 15350 18216
rect 15381 18207 15439 18213
rect 15381 18204 15393 18207
rect 15344 18176 15393 18204
rect 15344 18164 15350 18176
rect 15381 18173 15393 18176
rect 15427 18173 15439 18207
rect 15381 18167 15439 18173
rect 13817 18071 13875 18077
rect 13817 18068 13829 18071
rect 13648 18040 13829 18068
rect 13817 18037 13829 18040
rect 13863 18037 13875 18071
rect 14366 18068 14372 18080
rect 14327 18040 14372 18068
rect 13817 18031 13875 18037
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1762 17824 1768 17876
rect 1820 17824 1826 17876
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 3789 17867 3847 17873
rect 3789 17864 3801 17867
rect 2832 17836 3801 17864
rect 2832 17824 2838 17836
rect 3789 17833 3801 17836
rect 3835 17864 3847 17867
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 3835 17836 4077 17864
rect 3835 17833 3847 17836
rect 3789 17827 3847 17833
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 4706 17824 4712 17876
rect 4764 17864 4770 17876
rect 5077 17867 5135 17873
rect 5077 17864 5089 17867
rect 4764 17836 5089 17864
rect 4764 17824 4770 17836
rect 5077 17833 5089 17836
rect 5123 17833 5135 17867
rect 5626 17864 5632 17876
rect 5587 17836 5632 17864
rect 5077 17827 5135 17833
rect 5626 17824 5632 17836
rect 5684 17824 5690 17876
rect 11422 17824 11428 17876
rect 11480 17864 11486 17876
rect 11609 17867 11667 17873
rect 11609 17864 11621 17867
rect 11480 17836 11621 17864
rect 11480 17824 11486 17836
rect 11609 17833 11621 17836
rect 11655 17833 11667 17867
rect 13538 17864 13544 17876
rect 13499 17836 13544 17864
rect 11609 17827 11667 17833
rect 13538 17824 13544 17836
rect 13596 17824 13602 17876
rect 14366 17864 14372 17876
rect 14327 17836 14372 17864
rect 14366 17824 14372 17836
rect 14424 17824 14430 17876
rect 1780 17796 1808 17824
rect 1504 17768 1808 17796
rect 1504 17737 1532 17768
rect 3602 17756 3608 17808
rect 3660 17796 3666 17808
rect 4430 17796 4436 17808
rect 3660 17768 4436 17796
rect 3660 17756 3666 17768
rect 4430 17756 4436 17768
rect 4488 17756 4494 17808
rect 5828 17768 6408 17796
rect 1489 17731 1547 17737
rect 1489 17697 1501 17731
rect 1535 17697 1547 17731
rect 1489 17691 1547 17697
rect 1756 17731 1814 17737
rect 1756 17697 1768 17731
rect 1802 17728 1814 17731
rect 2038 17728 2044 17740
rect 1802 17700 2044 17728
rect 1802 17697 1814 17700
rect 1756 17691 1814 17697
rect 2038 17688 2044 17700
rect 2096 17688 2102 17740
rect 5828 17737 5856 17768
rect 6270 17737 6276 17740
rect 5813 17731 5871 17737
rect 5813 17697 5825 17731
rect 5859 17697 5871 17731
rect 6264 17728 6276 17737
rect 5813 17691 5871 17697
rect 5920 17700 6276 17728
rect 4246 17620 4252 17672
rect 4304 17660 4310 17672
rect 4525 17663 4583 17669
rect 4525 17660 4537 17663
rect 4304 17632 4537 17660
rect 4304 17620 4310 17632
rect 4525 17629 4537 17632
rect 4571 17629 4583 17663
rect 4706 17660 4712 17672
rect 4667 17632 4712 17660
rect 4525 17623 4583 17629
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 5537 17663 5595 17669
rect 5537 17629 5549 17663
rect 5583 17660 5595 17663
rect 5920 17660 5948 17700
rect 6264 17691 6276 17700
rect 6270 17688 6276 17691
rect 6328 17688 6334 17740
rect 6380 17728 6408 17768
rect 7374 17728 7380 17740
rect 6380 17700 7380 17728
rect 7374 17688 7380 17700
rect 7432 17728 7438 17740
rect 8018 17728 8024 17740
rect 7432 17700 8024 17728
rect 7432 17688 7438 17700
rect 8018 17688 8024 17700
rect 8076 17688 8082 17740
rect 9950 17737 9956 17740
rect 9493 17731 9551 17737
rect 9493 17697 9505 17731
rect 9539 17728 9551 17731
rect 9944 17728 9956 17737
rect 9539 17700 9956 17728
rect 9539 17697 9551 17700
rect 9493 17691 9551 17697
rect 9944 17691 9956 17700
rect 9950 17688 9956 17691
rect 10008 17688 10014 17740
rect 11054 17728 11060 17740
rect 10967 17700 11060 17728
rect 11054 17688 11060 17700
rect 11112 17728 11118 17740
rect 12428 17731 12486 17737
rect 12428 17728 12440 17731
rect 11112 17700 12440 17728
rect 11112 17688 11118 17700
rect 12428 17697 12440 17700
rect 12474 17728 12486 17731
rect 13538 17728 13544 17740
rect 12474 17700 13544 17728
rect 12474 17697 12486 17700
rect 12428 17691 12486 17697
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 5583 17632 5948 17660
rect 5997 17663 6055 17669
rect 5583 17629 5595 17632
rect 5537 17623 5595 17629
rect 5997 17629 6009 17663
rect 6043 17629 6055 17663
rect 7926 17660 7932 17672
rect 7887 17632 7932 17660
rect 5997 17623 6055 17629
rect 2869 17595 2927 17601
rect 2869 17561 2881 17595
rect 2915 17592 2927 17595
rect 2958 17592 2964 17604
rect 2915 17564 2964 17592
rect 2915 17561 2927 17564
rect 2869 17555 2927 17561
rect 2958 17552 2964 17564
rect 3016 17592 3022 17604
rect 3421 17595 3479 17601
rect 3421 17592 3433 17595
rect 3016 17564 3433 17592
rect 3016 17552 3022 17564
rect 3421 17561 3433 17564
rect 3467 17561 3479 17595
rect 3421 17555 3479 17561
rect 5626 17552 5632 17604
rect 5684 17592 5690 17604
rect 6012 17592 6040 17623
rect 7926 17620 7932 17632
rect 7984 17620 7990 17672
rect 8570 17660 8576 17672
rect 8531 17632 8576 17660
rect 8570 17620 8576 17632
rect 8628 17620 8634 17672
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 5684 17564 6040 17592
rect 5684 17552 5690 17564
rect 6012 17524 6040 17564
rect 6362 17524 6368 17536
rect 6012 17496 6368 17524
rect 6362 17484 6368 17496
rect 6420 17484 6426 17536
rect 7374 17524 7380 17536
rect 7335 17496 7380 17524
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 8294 17524 8300 17536
rect 8255 17496 8300 17524
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 9030 17524 9036 17536
rect 8991 17496 9036 17524
rect 9030 17484 9036 17496
rect 9088 17484 9094 17536
rect 9692 17524 9720 17623
rect 11072 17601 11100 17688
rect 12158 17660 12164 17672
rect 11992 17632 12164 17660
rect 11057 17595 11115 17601
rect 11057 17561 11069 17595
rect 11103 17561 11115 17595
rect 11057 17555 11115 17561
rect 11146 17524 11152 17536
rect 9692 17496 11152 17524
rect 11146 17484 11152 17496
rect 11204 17524 11210 17536
rect 11992 17533 12020 17632
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 11977 17527 12035 17533
rect 11977 17524 11989 17527
rect 11204 17496 11989 17524
rect 11204 17484 11210 17496
rect 11977 17493 11989 17496
rect 12023 17493 12035 17527
rect 11977 17487 12035 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2866 17320 2872 17332
rect 2827 17292 2872 17320
rect 2866 17280 2872 17292
rect 2924 17280 2930 17332
rect 4157 17323 4215 17329
rect 4157 17289 4169 17323
rect 4203 17320 4215 17323
rect 4246 17320 4252 17332
rect 4203 17292 4252 17320
rect 4203 17289 4215 17292
rect 4157 17283 4215 17289
rect 4246 17280 4252 17292
rect 4304 17280 4310 17332
rect 4430 17320 4436 17332
rect 4391 17292 4436 17320
rect 4430 17280 4436 17292
rect 4488 17280 4494 17332
rect 5166 17320 5172 17332
rect 5127 17292 5172 17320
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 6270 17320 6276 17332
rect 6231 17292 6276 17320
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 6362 17280 6368 17332
rect 6420 17320 6426 17332
rect 9398 17320 9404 17332
rect 6420 17292 6868 17320
rect 9359 17292 9404 17320
rect 6420 17280 6426 17292
rect 6730 17252 6736 17264
rect 5644 17224 6736 17252
rect 2038 17184 2044 17196
rect 1951 17156 2044 17184
rect 2038 17144 2044 17156
rect 2096 17184 2102 17196
rect 2409 17187 2467 17193
rect 2409 17184 2421 17187
rect 2096 17156 2421 17184
rect 2096 17144 2102 17156
rect 2409 17153 2421 17156
rect 2455 17184 2467 17187
rect 3513 17187 3571 17193
rect 3513 17184 3525 17187
rect 2455 17156 3525 17184
rect 2455 17153 2467 17156
rect 2409 17147 2467 17153
rect 3513 17153 3525 17156
rect 3559 17153 3571 17187
rect 3513 17147 3571 17153
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 3326 17116 3332 17128
rect 1443 17088 3332 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 3326 17076 3332 17088
rect 3384 17076 3390 17128
rect 3418 17076 3424 17128
rect 3476 17116 3482 17128
rect 3528 17116 3556 17147
rect 4614 17144 4620 17196
rect 4672 17184 4678 17196
rect 5644 17193 5672 17224
rect 6730 17212 6736 17224
rect 6788 17212 6794 17264
rect 6840 17193 6868 17292
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 11057 17323 11115 17329
rect 11057 17289 11069 17323
rect 11103 17320 11115 17323
rect 11330 17320 11336 17332
rect 11103 17292 11336 17320
rect 11103 17289 11115 17292
rect 11057 17283 11115 17289
rect 11330 17280 11336 17292
rect 11388 17280 11394 17332
rect 13538 17320 13544 17332
rect 13499 17292 13544 17320
rect 13538 17280 13544 17292
rect 13596 17280 13602 17332
rect 11885 17255 11943 17261
rect 11885 17221 11897 17255
rect 11931 17252 11943 17255
rect 12437 17255 12495 17261
rect 12437 17252 12449 17255
rect 11931 17224 12449 17252
rect 11931 17221 11943 17224
rect 11885 17215 11943 17221
rect 12437 17221 12449 17224
rect 12483 17221 12495 17255
rect 12437 17215 12495 17221
rect 5629 17187 5687 17193
rect 5629 17184 5641 17187
rect 4672 17156 5641 17184
rect 4672 17144 4678 17156
rect 5629 17153 5641 17156
rect 5675 17153 5687 17187
rect 5629 17147 5687 17153
rect 5813 17187 5871 17193
rect 5813 17153 5825 17187
rect 5859 17184 5871 17187
rect 6549 17187 6607 17193
rect 6549 17184 6561 17187
rect 5859 17156 6561 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 6549 17153 6561 17156
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17153 6883 17187
rect 9306 17184 9312 17196
rect 9219 17156 9312 17184
rect 6825 17147 6883 17153
rect 4706 17116 4712 17128
rect 3476 17088 4712 17116
rect 3476 17076 3482 17088
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 5534 17116 5540 17128
rect 5495 17088 5540 17116
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 2314 17008 2320 17060
rect 2372 17048 2378 17060
rect 2777 17051 2835 17057
rect 2777 17048 2789 17051
rect 2372 17020 2789 17048
rect 2372 17008 2378 17020
rect 2777 17017 2789 17020
rect 2823 17048 2835 17051
rect 6564 17048 6592 17147
rect 6840 17116 6868 17147
rect 9306 17144 9312 17156
rect 9364 17184 9370 17196
rect 9766 17184 9772 17196
rect 9364 17156 9772 17184
rect 9364 17144 9370 17156
rect 9766 17144 9772 17156
rect 9824 17184 9830 17196
rect 9861 17187 9919 17193
rect 9861 17184 9873 17187
rect 9824 17156 9873 17184
rect 9824 17144 9830 17156
rect 9861 17153 9873 17156
rect 9907 17153 9919 17187
rect 9861 17147 9919 17153
rect 8757 17119 8815 17125
rect 8757 17116 8769 17119
rect 6840 17088 8769 17116
rect 8757 17085 8769 17088
rect 8803 17116 8815 17119
rect 9030 17116 9036 17128
rect 8803 17088 9036 17116
rect 8803 17085 8815 17088
rect 8757 17079 8815 17085
rect 9030 17076 9036 17088
rect 9088 17076 9094 17128
rect 7092 17051 7150 17057
rect 7092 17048 7104 17051
rect 2823 17020 3372 17048
rect 6564 17020 7104 17048
rect 2823 17017 2835 17020
rect 2777 17011 2835 17017
rect 1578 16980 1584 16992
rect 1539 16952 1584 16980
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 3234 16980 3240 16992
rect 3195 16952 3240 16980
rect 3234 16940 3240 16952
rect 3292 16940 3298 16992
rect 3344 16989 3372 17020
rect 7092 17017 7104 17020
rect 7138 17048 7150 17051
rect 7374 17048 7380 17060
rect 7138 17020 7380 17048
rect 7138 17017 7150 17020
rect 7092 17011 7150 17017
rect 7374 17008 7380 17020
rect 7432 17008 7438 17060
rect 9876 17048 9904 17147
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 10045 17187 10103 17193
rect 10045 17184 10057 17187
rect 10008 17156 10057 17184
rect 10008 17144 10014 17156
rect 10045 17153 10057 17156
rect 10091 17184 10103 17187
rect 10091 17156 10548 17184
rect 10091 17153 10103 17156
rect 10045 17147 10103 17153
rect 10042 17048 10048 17060
rect 9876 17020 10048 17048
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 3329 16983 3387 16989
rect 3329 16949 3341 16983
rect 3375 16949 3387 16983
rect 3329 16943 3387 16949
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 4893 16983 4951 16989
rect 4893 16980 4905 16983
rect 4764 16952 4905 16980
rect 4764 16940 4770 16952
rect 4893 16949 4905 16952
rect 4939 16980 4951 16983
rect 5994 16980 6000 16992
rect 4939 16952 6000 16980
rect 4939 16949 4951 16952
rect 4893 16943 4951 16949
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 8202 16980 8208 16992
rect 8163 16952 8208 16980
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 9766 16980 9772 16992
rect 9727 16952 9772 16980
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 10520 16989 10548 17156
rect 11238 17144 11244 17196
rect 11296 17184 11302 17196
rect 11333 17187 11391 17193
rect 11333 17184 11345 17187
rect 11296 17156 11345 17184
rect 11296 17144 11302 17156
rect 11333 17153 11345 17156
rect 11379 17153 11391 17187
rect 11333 17147 11391 17153
rect 12253 17187 12311 17193
rect 12253 17153 12265 17187
rect 12299 17184 12311 17187
rect 12986 17184 12992 17196
rect 12299 17156 12992 17184
rect 12299 17153 12311 17156
rect 12253 17147 12311 17153
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 13173 17187 13231 17193
rect 13173 17153 13185 17187
rect 13219 17184 13231 17187
rect 13446 17184 13452 17196
rect 13219 17156 13452 17184
rect 13219 17153 13231 17156
rect 13173 17147 13231 17153
rect 13446 17144 13452 17156
rect 13504 17144 13510 17196
rect 14366 17184 14372 17196
rect 14327 17156 14372 17184
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 12437 17051 12495 17057
rect 12437 17017 12449 17051
rect 12483 17048 12495 17051
rect 14614 17051 14672 17057
rect 14614 17048 14626 17051
rect 12483 17020 12940 17048
rect 12483 17017 12495 17020
rect 12437 17011 12495 17017
rect 10505 16983 10563 16989
rect 10505 16949 10517 16983
rect 10551 16980 10563 16983
rect 10686 16980 10692 16992
rect 10551 16952 10692 16980
rect 10551 16949 10563 16952
rect 10505 16943 10563 16949
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 12526 16980 12532 16992
rect 12487 16952 12532 16980
rect 12526 16940 12532 16952
rect 12584 16940 12590 16992
rect 12912 16989 12940 17020
rect 14200 17020 14626 17048
rect 14200 16992 14228 17020
rect 14614 17017 14626 17020
rect 14660 17017 14672 17051
rect 14614 17011 14672 17017
rect 12897 16983 12955 16989
rect 12897 16949 12909 16983
rect 12943 16980 12955 16983
rect 13170 16980 13176 16992
rect 12943 16952 13176 16980
rect 12943 16949 12955 16952
rect 12897 16943 12955 16949
rect 13170 16940 13176 16952
rect 13228 16940 13234 16992
rect 14182 16980 14188 16992
rect 14143 16952 14188 16980
rect 14182 16940 14188 16952
rect 14240 16940 14246 16992
rect 15746 16980 15752 16992
rect 15707 16952 15752 16980
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1857 16779 1915 16785
rect 1857 16745 1869 16779
rect 1903 16776 1915 16779
rect 2498 16776 2504 16788
rect 1903 16748 2504 16776
rect 1903 16745 1915 16748
rect 1857 16739 1915 16745
rect 2498 16736 2504 16748
rect 2556 16736 2562 16788
rect 3326 16776 3332 16788
rect 3287 16748 3332 16776
rect 3326 16736 3332 16748
rect 3384 16736 3390 16788
rect 3694 16736 3700 16788
rect 3752 16776 3758 16788
rect 4065 16779 4123 16785
rect 4065 16776 4077 16779
rect 3752 16748 4077 16776
rect 3752 16736 3758 16748
rect 4065 16745 4077 16748
rect 4111 16745 4123 16779
rect 4614 16776 4620 16788
rect 4575 16748 4620 16776
rect 4065 16739 4123 16745
rect 4614 16736 4620 16748
rect 4672 16736 4678 16788
rect 5074 16776 5080 16788
rect 5035 16748 5080 16776
rect 5074 16736 5080 16748
rect 5132 16736 5138 16788
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 6089 16779 6147 16785
rect 6089 16776 6101 16779
rect 5592 16748 6101 16776
rect 5592 16736 5598 16748
rect 6089 16745 6101 16748
rect 6135 16745 6147 16779
rect 6638 16776 6644 16788
rect 6599 16748 6644 16776
rect 6089 16739 6147 16745
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7009 16779 7067 16785
rect 7009 16776 7021 16779
rect 6972 16748 7021 16776
rect 6972 16736 6978 16748
rect 7009 16745 7021 16748
rect 7055 16745 7067 16779
rect 8018 16776 8024 16788
rect 7979 16748 8024 16776
rect 7009 16739 7067 16745
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 8570 16736 8576 16788
rect 8628 16776 8634 16788
rect 9401 16779 9459 16785
rect 9401 16776 9413 16779
rect 8628 16748 9413 16776
rect 8628 16736 8634 16748
rect 9401 16745 9413 16748
rect 9447 16776 9459 16779
rect 9766 16776 9772 16788
rect 9447 16748 9772 16776
rect 9447 16745 9459 16748
rect 9401 16739 9459 16745
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 10137 16779 10195 16785
rect 10137 16745 10149 16779
rect 10183 16745 10195 16779
rect 10137 16739 10195 16745
rect 2225 16711 2283 16717
rect 2225 16677 2237 16711
rect 2271 16708 2283 16711
rect 2590 16708 2596 16720
rect 2271 16680 2596 16708
rect 2271 16677 2283 16680
rect 2225 16671 2283 16677
rect 2590 16668 2596 16680
rect 2648 16668 2654 16720
rect 2682 16668 2688 16720
rect 2740 16708 2746 16720
rect 3605 16711 3663 16717
rect 3605 16708 3617 16711
rect 2740 16680 3617 16708
rect 2740 16668 2746 16680
rect 3605 16677 3617 16680
rect 3651 16677 3663 16711
rect 7101 16711 7159 16717
rect 7101 16708 7113 16711
rect 3605 16671 3663 16677
rect 6932 16680 7113 16708
rect 2130 16600 2136 16652
rect 2188 16640 2194 16652
rect 2317 16643 2375 16649
rect 2317 16640 2329 16643
rect 2188 16612 2329 16640
rect 2188 16600 2194 16612
rect 2317 16609 2329 16612
rect 2363 16609 2375 16643
rect 2317 16603 2375 16609
rect 2406 16600 2412 16652
rect 2464 16640 2470 16652
rect 2869 16643 2927 16649
rect 2869 16640 2881 16643
rect 2464 16612 2881 16640
rect 2464 16600 2470 16612
rect 2869 16609 2881 16612
rect 2915 16640 2927 16643
rect 3234 16640 3240 16652
rect 2915 16612 3240 16640
rect 2915 16609 2927 16612
rect 2869 16603 2927 16609
rect 3234 16600 3240 16612
rect 3292 16600 3298 16652
rect 5442 16640 5448 16652
rect 5403 16612 5448 16640
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16640 6607 16643
rect 6822 16640 6828 16652
rect 6595 16612 6828 16640
rect 6595 16609 6607 16612
rect 6549 16603 6607 16609
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 2501 16575 2559 16581
rect 2501 16541 2513 16575
rect 2547 16572 2559 16575
rect 3418 16572 3424 16584
rect 2547 16544 3424 16572
rect 2547 16541 2559 16544
rect 2501 16535 2559 16541
rect 3418 16532 3424 16544
rect 3476 16532 3482 16584
rect 5074 16532 5080 16584
rect 5132 16572 5138 16584
rect 5537 16575 5595 16581
rect 5537 16572 5549 16575
rect 5132 16544 5549 16572
rect 5132 16532 5138 16544
rect 5537 16541 5549 16544
rect 5583 16541 5595 16575
rect 5537 16535 5595 16541
rect 5629 16575 5687 16581
rect 5629 16541 5641 16575
rect 5675 16541 5687 16575
rect 6932 16572 6960 16680
rect 7101 16677 7113 16680
rect 7147 16677 7159 16711
rect 7101 16671 7159 16677
rect 9030 16668 9036 16720
rect 9088 16708 9094 16720
rect 9088 16680 9628 16708
rect 9088 16668 9094 16680
rect 8297 16643 8355 16649
rect 8297 16609 8309 16643
rect 8343 16640 8355 16643
rect 8570 16640 8576 16652
rect 8343 16612 8576 16640
rect 8343 16609 8355 16612
rect 8297 16603 8355 16609
rect 8570 16600 8576 16612
rect 8628 16640 8634 16652
rect 9214 16640 9220 16652
rect 8628 16612 9220 16640
rect 8628 16600 8634 16612
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 9600 16640 9628 16680
rect 9674 16668 9680 16720
rect 9732 16708 9738 16720
rect 10152 16708 10180 16739
rect 11422 16736 11428 16788
rect 11480 16776 11486 16788
rect 12069 16779 12127 16785
rect 12069 16776 12081 16779
rect 11480 16748 12081 16776
rect 11480 16736 11486 16748
rect 12069 16745 12081 16748
rect 12115 16745 12127 16779
rect 12069 16739 12127 16745
rect 13814 16736 13820 16788
rect 13872 16776 13878 16788
rect 14093 16779 14151 16785
rect 14093 16776 14105 16779
rect 13872 16748 14105 16776
rect 13872 16736 13878 16748
rect 14093 16745 14105 16748
rect 14139 16776 14151 16779
rect 14826 16776 14832 16788
rect 14139 16748 14832 16776
rect 14139 16745 14151 16748
rect 14093 16739 14151 16745
rect 14826 16736 14832 16748
rect 14884 16736 14890 16788
rect 9732 16680 10180 16708
rect 10597 16711 10655 16717
rect 9732 16668 9738 16680
rect 10597 16677 10609 16711
rect 10643 16708 10655 16711
rect 10778 16708 10784 16720
rect 10643 16680 10784 16708
rect 10643 16677 10655 16680
rect 10597 16671 10655 16677
rect 10778 16668 10784 16680
rect 10836 16708 10842 16720
rect 13173 16711 13231 16717
rect 10836 16680 13032 16708
rect 10836 16668 10842 16680
rect 9861 16643 9919 16649
rect 9861 16640 9873 16643
rect 9600 16612 9873 16640
rect 9861 16609 9873 16612
rect 9907 16609 9919 16643
rect 9861 16603 9919 16609
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16640 10563 16643
rect 10962 16640 10968 16652
rect 10551 16612 10968 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 11112 16612 11161 16640
rect 11112 16600 11118 16612
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 11606 16640 11612 16652
rect 11567 16612 11612 16640
rect 11149 16603 11207 16609
rect 11606 16600 11612 16612
rect 11664 16640 11670 16652
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 11664 16612 11897 16640
rect 11664 16600 11670 16612
rect 11885 16609 11897 16612
rect 11931 16609 11943 16643
rect 12437 16643 12495 16649
rect 12437 16640 12449 16643
rect 11885 16603 11943 16609
rect 12360 16612 12449 16640
rect 7282 16572 7288 16584
rect 5629 16535 5687 16541
rect 6564 16544 6960 16572
rect 7195 16544 7288 16572
rect 5644 16504 5672 16535
rect 6564 16516 6592 16544
rect 7282 16532 7288 16544
rect 7340 16572 7346 16584
rect 8478 16572 8484 16584
rect 7340 16544 7788 16572
rect 8439 16544 8484 16572
rect 7340 16532 7346 16544
rect 5000 16476 5672 16504
rect 5000 16448 5028 16476
rect 6546 16464 6552 16516
rect 6604 16464 6610 16516
rect 7760 16448 7788 16544
rect 8478 16532 8484 16544
rect 8536 16532 8542 16584
rect 10686 16572 10692 16584
rect 10647 16544 10692 16572
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 12158 16572 12164 16584
rect 11756 16544 12164 16572
rect 11756 16532 11762 16544
rect 12158 16532 12164 16544
rect 12216 16572 12222 16584
rect 12360 16572 12388 16612
rect 12437 16609 12449 16612
rect 12483 16609 12495 16643
rect 13004 16640 13032 16680
rect 13173 16677 13185 16711
rect 13219 16708 13231 16711
rect 13446 16708 13452 16720
rect 13219 16680 13452 16708
rect 13219 16677 13231 16680
rect 13173 16671 13231 16677
rect 13446 16668 13452 16680
rect 13504 16668 13510 16720
rect 13630 16668 13636 16720
rect 13688 16708 13694 16720
rect 14001 16711 14059 16717
rect 14001 16708 14013 16711
rect 13688 16680 14013 16708
rect 13688 16668 13694 16680
rect 14001 16677 14013 16680
rect 14047 16677 14059 16711
rect 14001 16671 14059 16677
rect 13004 16612 13676 16640
rect 12437 16603 12495 16609
rect 12526 16572 12532 16584
rect 12216 16544 12388 16572
rect 12487 16544 12532 16572
rect 12216 16532 12222 16544
rect 12526 16532 12532 16544
rect 12584 16532 12590 16584
rect 12618 16532 12624 16584
rect 12676 16572 12682 16584
rect 12676 16544 12721 16572
rect 12676 16532 12682 16544
rect 13648 16513 13676 16612
rect 14182 16532 14188 16584
rect 14240 16572 14246 16584
rect 14240 16544 14285 16572
rect 14240 16532 14246 16544
rect 13633 16507 13691 16513
rect 13633 16473 13645 16507
rect 13679 16473 13691 16507
rect 13633 16467 13691 16473
rect 1673 16439 1731 16445
rect 1673 16405 1685 16439
rect 1719 16436 1731 16439
rect 2038 16436 2044 16448
rect 1719 16408 2044 16436
rect 1719 16405 1731 16408
rect 1673 16399 1731 16405
rect 2038 16396 2044 16408
rect 2096 16396 2102 16448
rect 4982 16436 4988 16448
rect 4943 16408 4988 16436
rect 4982 16396 4988 16408
rect 5040 16396 5046 16448
rect 7742 16436 7748 16448
rect 7703 16408 7748 16436
rect 7742 16396 7748 16408
rect 7800 16396 7806 16448
rect 9122 16436 9128 16448
rect 9083 16408 9128 16436
rect 9122 16396 9128 16408
rect 9180 16396 9186 16448
rect 11054 16396 11060 16448
rect 11112 16436 11118 16448
rect 11701 16439 11759 16445
rect 11701 16436 11713 16439
rect 11112 16408 11713 16436
rect 11112 16396 11118 16408
rect 11701 16405 11713 16408
rect 11747 16436 11759 16439
rect 12250 16436 12256 16448
rect 11747 16408 12256 16436
rect 11747 16405 11759 16408
rect 11701 16399 11759 16405
rect 12250 16396 12256 16408
rect 12308 16396 12314 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2961 16235 3019 16241
rect 2961 16201 2973 16235
rect 3007 16232 3019 16235
rect 3418 16232 3424 16244
rect 3007 16204 3424 16232
rect 3007 16201 3019 16204
rect 2961 16195 3019 16201
rect 3418 16192 3424 16204
rect 3476 16192 3482 16244
rect 6273 16235 6331 16241
rect 6273 16201 6285 16235
rect 6319 16232 6331 16235
rect 6730 16232 6736 16244
rect 6319 16204 6736 16232
rect 6319 16201 6331 16204
rect 6273 16195 6331 16201
rect 6730 16192 6736 16204
rect 6788 16192 6794 16244
rect 7742 16192 7748 16244
rect 7800 16232 7806 16244
rect 7837 16235 7895 16241
rect 7837 16232 7849 16235
rect 7800 16204 7849 16232
rect 7800 16192 7806 16204
rect 7837 16201 7849 16204
rect 7883 16201 7895 16235
rect 7837 16195 7895 16201
rect 10597 16235 10655 16241
rect 10597 16201 10609 16235
rect 10643 16232 10655 16235
rect 10686 16232 10692 16244
rect 10643 16204 10692 16232
rect 10643 16201 10655 16204
rect 10597 16195 10655 16201
rect 10686 16192 10692 16204
rect 10744 16192 10750 16244
rect 12989 16235 13047 16241
rect 12989 16201 13001 16235
rect 13035 16232 13047 16235
rect 14182 16232 14188 16244
rect 13035 16204 14188 16232
rect 13035 16201 13047 16204
rect 12989 16195 13047 16201
rect 14182 16192 14188 16204
rect 14240 16232 14246 16244
rect 15289 16235 15347 16241
rect 15289 16232 15301 16235
rect 14240 16204 15301 16232
rect 14240 16192 14246 16204
rect 15289 16201 15301 16204
rect 15335 16201 15347 16235
rect 15289 16195 15347 16201
rect 13722 16164 13728 16176
rect 13683 16136 13728 16164
rect 13722 16124 13728 16136
rect 13780 16124 13786 16176
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 5442 16056 5448 16108
rect 5500 16096 5506 16108
rect 5537 16099 5595 16105
rect 5537 16096 5549 16099
rect 5500 16068 5549 16096
rect 5500 16056 5506 16068
rect 5537 16065 5549 16068
rect 5583 16065 5595 16099
rect 7374 16096 7380 16108
rect 7335 16068 7380 16096
rect 5537 16059 5595 16065
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 9398 16096 9404 16108
rect 9359 16068 9404 16096
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 11146 16056 11152 16108
rect 11204 16096 11210 16108
rect 11241 16099 11299 16105
rect 11241 16096 11253 16099
rect 11204 16068 11253 16096
rect 11204 16056 11210 16068
rect 11241 16065 11253 16068
rect 11287 16065 11299 16099
rect 11241 16059 11299 16065
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16096 13415 16099
rect 13630 16096 13636 16108
rect 13403 16068 13636 16096
rect 13403 16065 13415 16068
rect 13357 16059 13415 16065
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 16669 16099 16727 16105
rect 16669 16065 16681 16099
rect 16715 16096 16727 16099
rect 16758 16096 16764 16108
rect 16715 16068 16764 16096
rect 16715 16065 16727 16068
rect 16669 16059 16727 16065
rect 16758 16056 16764 16068
rect 16816 16056 16822 16108
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 16028 2007 16031
rect 2130 16028 2136 16040
rect 1995 16000 2136 16028
rect 1995 15997 2007 16000
rect 1949 15991 2007 15997
rect 2130 15988 2136 16000
rect 2188 16028 2194 16040
rect 2682 16028 2688 16040
rect 2188 16000 2688 16028
rect 2188 15988 2194 16000
rect 2682 15988 2688 16000
rect 2740 15988 2746 16040
rect 3053 16031 3111 16037
rect 3053 15997 3065 16031
rect 3099 15997 3111 16031
rect 3053 15991 3111 15997
rect 3068 15960 3096 15991
rect 3142 15988 3148 16040
rect 3200 16028 3206 16040
rect 3309 16031 3367 16037
rect 3309 16028 3321 16031
rect 3200 16000 3321 16028
rect 3200 15988 3206 16000
rect 3309 15997 3321 16000
rect 3355 15997 3367 16031
rect 7190 16028 7196 16040
rect 7151 16000 7196 16028
rect 3309 15991 3367 15997
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 8757 16031 8815 16037
rect 8757 15997 8769 16031
rect 8803 16028 8815 16031
rect 9214 16028 9220 16040
rect 8803 16000 9220 16028
rect 8803 15997 8815 16000
rect 8757 15991 8815 15997
rect 9214 15988 9220 16000
rect 9272 15988 9278 16040
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 16028 11023 16031
rect 11057 16031 11115 16037
rect 11057 16028 11069 16031
rect 11011 16000 11069 16028
rect 11011 15997 11023 16000
rect 10965 15991 11023 15997
rect 11057 15997 11069 16000
rect 11103 16028 11115 16031
rect 11330 16028 11336 16040
rect 11103 16000 11336 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 11330 15988 11336 16000
rect 11388 15988 11394 16040
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 16028 13967 16031
rect 13955 16000 14412 16028
rect 13955 15997 13967 16000
rect 13909 15991 13967 15997
rect 14384 15972 14412 16000
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 16393 16031 16451 16037
rect 16393 16028 16405 16031
rect 16356 16000 16405 16028
rect 16356 15988 16362 16000
rect 16393 15997 16405 16000
rect 16439 16028 16451 16031
rect 17129 16031 17187 16037
rect 17129 16028 17141 16031
rect 16439 16000 17141 16028
rect 16439 15997 16451 16000
rect 16393 15991 16451 15997
rect 17129 15997 17141 16000
rect 17175 15997 17187 16031
rect 17129 15991 17187 15997
rect 5258 15960 5264 15972
rect 3068 15932 5264 15960
rect 5258 15920 5264 15932
rect 5316 15920 5322 15972
rect 6914 15920 6920 15972
rect 6972 15960 6978 15972
rect 14182 15969 14188 15972
rect 7285 15963 7343 15969
rect 7285 15960 7297 15963
rect 6972 15932 7297 15960
rect 6972 15920 6978 15932
rect 7285 15929 7297 15932
rect 7331 15929 7343 15963
rect 9309 15963 9367 15969
rect 9309 15960 9321 15963
rect 7285 15923 7343 15929
rect 8312 15932 9321 15960
rect 8312 15904 8340 15932
rect 9309 15929 9321 15932
rect 9355 15929 9367 15963
rect 14176 15960 14188 15969
rect 14143 15932 14188 15960
rect 9309 15923 9367 15929
rect 14176 15923 14188 15932
rect 14182 15920 14188 15923
rect 14240 15920 14246 15972
rect 14366 15920 14372 15972
rect 14424 15920 14430 15972
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 1854 15892 1860 15904
rect 1815 15864 1860 15892
rect 1854 15852 1860 15864
rect 1912 15852 1918 15904
rect 2593 15895 2651 15901
rect 2593 15861 2605 15895
rect 2639 15892 2651 15895
rect 2682 15892 2688 15904
rect 2639 15864 2688 15892
rect 2639 15861 2651 15864
rect 2593 15855 2651 15861
rect 2682 15852 2688 15864
rect 2740 15852 2746 15904
rect 3510 15852 3516 15904
rect 3568 15892 3574 15904
rect 4433 15895 4491 15901
rect 4433 15892 4445 15895
rect 3568 15864 4445 15892
rect 3568 15852 3574 15864
rect 4433 15861 4445 15864
rect 4479 15861 4491 15895
rect 5074 15892 5080 15904
rect 5035 15864 5080 15892
rect 4433 15855 4491 15861
rect 5074 15852 5080 15864
rect 5132 15852 5138 15904
rect 6546 15892 6552 15904
rect 6507 15864 6552 15892
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 6822 15892 6828 15904
rect 6783 15864 6828 15892
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 8294 15892 8300 15904
rect 8255 15864 8300 15892
rect 8294 15852 8300 15864
rect 8352 15852 8358 15904
rect 8846 15892 8852 15904
rect 8807 15864 8852 15892
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 9214 15892 9220 15904
rect 9175 15864 9220 15892
rect 9214 15852 9220 15864
rect 9272 15892 9278 15904
rect 10137 15895 10195 15901
rect 10137 15892 10149 15895
rect 9272 15864 10149 15892
rect 9272 15852 9278 15864
rect 10137 15861 10149 15864
rect 10183 15892 10195 15895
rect 10962 15892 10968 15904
rect 10183 15864 10968 15892
rect 10183 15861 10195 15864
rect 10137 15855 10195 15861
rect 10962 15852 10968 15864
rect 11020 15852 11026 15904
rect 12158 15892 12164 15904
rect 12119 15864 12164 15892
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2041 15691 2099 15697
rect 2041 15657 2053 15691
rect 2087 15688 2099 15691
rect 2130 15688 2136 15700
rect 2087 15660 2136 15688
rect 2087 15657 2099 15660
rect 2041 15651 2099 15657
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 3142 15688 3148 15700
rect 3103 15660 3148 15688
rect 3142 15648 3148 15660
rect 3200 15648 3206 15700
rect 3510 15688 3516 15700
rect 3471 15660 3516 15688
rect 3510 15648 3516 15660
rect 3568 15648 3574 15700
rect 4249 15691 4307 15697
rect 4249 15657 4261 15691
rect 4295 15688 4307 15691
rect 4522 15688 4528 15700
rect 4295 15660 4528 15688
rect 4295 15657 4307 15660
rect 4249 15651 4307 15657
rect 4522 15648 4528 15660
rect 4580 15648 4586 15700
rect 5169 15691 5227 15697
rect 5169 15657 5181 15691
rect 5215 15688 5227 15691
rect 5442 15688 5448 15700
rect 5215 15660 5448 15688
rect 5215 15657 5227 15660
rect 5169 15651 5227 15657
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 5994 15648 6000 15700
rect 6052 15688 6058 15700
rect 6641 15691 6699 15697
rect 6641 15688 6653 15691
rect 6052 15660 6653 15688
rect 6052 15648 6058 15660
rect 6641 15657 6653 15660
rect 6687 15657 6699 15691
rect 6641 15651 6699 15657
rect 6730 15648 6736 15700
rect 6788 15688 6794 15700
rect 7285 15691 7343 15697
rect 7285 15688 7297 15691
rect 6788 15660 7297 15688
rect 6788 15648 6794 15660
rect 7285 15657 7297 15660
rect 7331 15688 7343 15691
rect 7374 15688 7380 15700
rect 7331 15660 7380 15688
rect 7331 15657 7343 15660
rect 7285 15651 7343 15657
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 8570 15688 8576 15700
rect 8531 15660 8576 15688
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 8941 15691 8999 15697
rect 8941 15657 8953 15691
rect 8987 15688 8999 15691
rect 9398 15688 9404 15700
rect 8987 15660 9404 15688
rect 8987 15657 8999 15660
rect 8941 15651 8999 15657
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 10042 15648 10048 15700
rect 10100 15688 10106 15700
rect 10137 15691 10195 15697
rect 10137 15688 10149 15691
rect 10100 15660 10149 15688
rect 10100 15648 10106 15660
rect 10137 15657 10149 15660
rect 10183 15657 10195 15691
rect 10778 15688 10784 15700
rect 10739 15660 10784 15688
rect 10137 15651 10195 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 11330 15688 11336 15700
rect 11291 15660 11336 15688
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 12713 15691 12771 15697
rect 12713 15688 12725 15691
rect 12584 15660 12725 15688
rect 12584 15648 12590 15660
rect 12713 15657 12725 15660
rect 12759 15657 12771 15691
rect 12713 15651 12771 15657
rect 13078 15648 13084 15700
rect 13136 15688 13142 15700
rect 13357 15691 13415 15697
rect 13357 15688 13369 15691
rect 13136 15660 13369 15688
rect 13136 15648 13142 15660
rect 13357 15657 13369 15660
rect 13403 15657 13415 15691
rect 13357 15651 13415 15657
rect 14366 15648 14372 15700
rect 14424 15688 14430 15700
rect 14645 15691 14703 15697
rect 14645 15688 14657 15691
rect 14424 15660 14657 15688
rect 14424 15648 14430 15660
rect 14645 15657 14657 15660
rect 14691 15657 14703 15691
rect 14645 15651 14703 15657
rect 1854 15580 1860 15632
rect 1912 15620 1918 15632
rect 3789 15623 3847 15629
rect 3789 15620 3801 15623
rect 1912 15592 3801 15620
rect 1912 15580 1918 15592
rect 3789 15589 3801 15592
rect 3835 15589 3847 15623
rect 3789 15583 3847 15589
rect 12437 15623 12495 15629
rect 12437 15589 12449 15623
rect 12483 15620 12495 15623
rect 12618 15620 12624 15632
rect 12483 15592 12624 15620
rect 12483 15589 12495 15592
rect 12437 15583 12495 15589
rect 12618 15580 12624 15592
rect 12676 15580 12682 15632
rect 15470 15580 15476 15632
rect 15528 15620 15534 15632
rect 15565 15623 15623 15629
rect 15565 15620 15577 15623
rect 15528 15592 15577 15620
rect 15528 15580 15534 15592
rect 15565 15589 15577 15592
rect 15611 15589 15623 15623
rect 15565 15583 15623 15589
rect 2222 15552 2228 15564
rect 2135 15524 2228 15552
rect 2222 15512 2228 15524
rect 2280 15552 2286 15564
rect 2409 15555 2467 15561
rect 2409 15552 2421 15555
rect 2280 15524 2421 15552
rect 2280 15512 2286 15524
rect 2409 15521 2421 15524
rect 2455 15521 2467 15555
rect 4062 15552 4068 15564
rect 4023 15524 4068 15552
rect 2409 15515 2467 15521
rect 4062 15512 4068 15524
rect 4120 15552 4126 15564
rect 4246 15552 4252 15564
rect 4120 15524 4252 15552
rect 4120 15512 4126 15524
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 5534 15561 5540 15564
rect 5528 15552 5540 15561
rect 5495 15524 5540 15552
rect 5528 15515 5540 15524
rect 5534 15512 5540 15515
rect 5592 15512 5598 15564
rect 7742 15552 7748 15564
rect 7703 15524 7748 15552
rect 7742 15512 7748 15524
rect 7800 15512 7806 15564
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9732 15524 10057 15552
rect 9732 15512 9738 15524
rect 10045 15521 10057 15524
rect 10091 15552 10103 15555
rect 10870 15552 10876 15564
rect 10091 15524 10876 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 11698 15552 11704 15564
rect 11659 15524 11704 15552
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 13262 15552 13268 15564
rect 13223 15524 13268 15552
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 15286 15552 15292 15564
rect 15247 15524 15292 15552
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 1949 15351 2007 15357
rect 1949 15317 1961 15351
rect 1995 15348 2007 15351
rect 2240 15348 2268 15512
rect 2314 15444 2320 15496
rect 2372 15484 2378 15496
rect 2501 15487 2559 15493
rect 2501 15484 2513 15487
rect 2372 15456 2513 15484
rect 2372 15444 2378 15456
rect 2501 15453 2513 15456
rect 2547 15484 2559 15487
rect 2590 15484 2596 15496
rect 2547 15456 2596 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15484 2743 15487
rect 3510 15484 3516 15496
rect 2731 15456 3516 15484
rect 2731 15453 2743 15456
rect 2685 15447 2743 15453
rect 3510 15444 3516 15456
rect 3568 15444 3574 15496
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15484 4767 15487
rect 5258 15484 5264 15496
rect 4755 15456 5264 15484
rect 4755 15453 4767 15456
rect 4709 15447 4767 15453
rect 5258 15444 5264 15456
rect 5316 15444 5322 15496
rect 7926 15484 7932 15496
rect 7887 15456 7932 15484
rect 7926 15444 7932 15456
rect 7984 15444 7990 15496
rect 9398 15444 9404 15496
rect 9456 15484 9462 15496
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 9456 15456 10241 15484
rect 9456 15444 9462 15456
rect 10229 15453 10241 15456
rect 10275 15484 10287 15487
rect 10502 15484 10508 15496
rect 10275 15456 10508 15484
rect 10275 15453 10287 15456
rect 10229 15447 10287 15453
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 11790 15484 11796 15496
rect 11751 15456 11796 15484
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 11882 15444 11888 15496
rect 11940 15484 11946 15496
rect 11940 15456 11985 15484
rect 11940 15444 11946 15456
rect 13354 15444 13360 15496
rect 13412 15484 13418 15496
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 13412 15456 13461 15484
rect 13412 15444 13418 15456
rect 13449 15453 13461 15456
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 11900 15416 11928 15444
rect 14001 15419 14059 15425
rect 14001 15416 14013 15419
rect 11900 15388 14013 15416
rect 14001 15385 14013 15388
rect 14047 15416 14059 15419
rect 14182 15416 14188 15428
rect 14047 15388 14188 15416
rect 14047 15385 14059 15388
rect 14001 15379 14059 15385
rect 14182 15376 14188 15388
rect 14240 15376 14246 15428
rect 3418 15348 3424 15360
rect 1995 15320 3424 15348
rect 1995 15317 2007 15320
rect 1949 15311 2007 15317
rect 3418 15308 3424 15320
rect 3476 15308 3482 15360
rect 7653 15351 7711 15357
rect 7653 15317 7665 15351
rect 7699 15348 7711 15351
rect 8110 15348 8116 15360
rect 7699 15320 8116 15348
rect 7699 15317 7711 15320
rect 7653 15311 7711 15317
rect 8110 15308 8116 15320
rect 8168 15308 8174 15360
rect 9214 15348 9220 15360
rect 9175 15320 9220 15348
rect 9214 15308 9220 15320
rect 9272 15308 9278 15360
rect 9677 15351 9735 15357
rect 9677 15317 9689 15351
rect 9723 15348 9735 15351
rect 9766 15348 9772 15360
rect 9723 15320 9772 15348
rect 9723 15317 9735 15320
rect 9677 15311 9735 15317
rect 9766 15308 9772 15320
rect 9824 15308 9830 15360
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 11149 15351 11207 15357
rect 11149 15348 11161 15351
rect 11112 15320 11161 15348
rect 11112 15308 11118 15320
rect 11149 15317 11161 15320
rect 11195 15348 11207 15351
rect 12250 15348 12256 15360
rect 11195 15320 12256 15348
rect 11195 15317 11207 15320
rect 11149 15311 11207 15317
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 12894 15348 12900 15360
rect 12855 15320 12900 15348
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 14274 15348 14280 15360
rect 14235 15320 14280 15348
rect 14274 15308 14280 15320
rect 14332 15308 14338 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 5534 15104 5540 15156
rect 5592 15144 5598 15156
rect 5629 15147 5687 15153
rect 5629 15144 5641 15147
rect 5592 15116 5641 15144
rect 5592 15104 5598 15116
rect 5629 15113 5641 15116
rect 5675 15144 5687 15147
rect 6273 15147 6331 15153
rect 6273 15144 6285 15147
rect 5675 15116 6285 15144
rect 5675 15113 5687 15116
rect 5629 15107 5687 15113
rect 6273 15113 6285 15116
rect 6319 15144 6331 15147
rect 6730 15144 6736 15156
rect 6319 15116 6736 15144
rect 6319 15113 6331 15116
rect 6273 15107 6331 15113
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 7101 15147 7159 15153
rect 7101 15113 7113 15147
rect 7147 15144 7159 15147
rect 7190 15144 7196 15156
rect 7147 15116 7196 15144
rect 7147 15113 7159 15116
rect 7101 15107 7159 15113
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 7561 15147 7619 15153
rect 7561 15113 7573 15147
rect 7607 15144 7619 15147
rect 8202 15144 8208 15156
rect 7607 15116 8208 15144
rect 7607 15113 7619 15116
rect 7561 15107 7619 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 9033 15147 9091 15153
rect 9033 15113 9045 15147
rect 9079 15144 9091 15147
rect 9490 15144 9496 15156
rect 9079 15116 9496 15144
rect 9079 15113 9091 15116
rect 9033 15107 9091 15113
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 10502 15144 10508 15156
rect 10463 15116 10508 15144
rect 10502 15104 10508 15116
rect 10560 15144 10566 15156
rect 10686 15144 10692 15156
rect 10560 15116 10692 15144
rect 10560 15104 10566 15116
rect 10686 15104 10692 15116
rect 10744 15144 10750 15156
rect 11057 15147 11115 15153
rect 11057 15144 11069 15147
rect 10744 15116 11069 15144
rect 10744 15104 10750 15116
rect 11057 15113 11069 15116
rect 11103 15113 11115 15147
rect 11057 15107 11115 15113
rect 11517 15147 11575 15153
rect 11517 15113 11529 15147
rect 11563 15144 11575 15147
rect 11882 15144 11888 15156
rect 11563 15116 11888 15144
rect 11563 15113 11575 15116
rect 11517 15107 11575 15113
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 13078 15144 13084 15156
rect 13039 15116 13084 15144
rect 13078 15104 13084 15116
rect 13136 15104 13142 15156
rect 14182 15104 14188 15156
rect 14240 15144 14246 15156
rect 14921 15147 14979 15153
rect 14921 15144 14933 15147
rect 14240 15116 14933 15144
rect 14240 15104 14246 15116
rect 14921 15113 14933 15116
rect 14967 15113 14979 15147
rect 14921 15107 14979 15113
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 15473 15147 15531 15153
rect 15473 15144 15485 15147
rect 15344 15116 15485 15144
rect 15344 15104 15350 15116
rect 15473 15113 15485 15116
rect 15519 15113 15531 15147
rect 21818 15144 21824 15156
rect 21779 15116 21824 15144
rect 15473 15107 15531 15113
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 7374 15008 7380 15020
rect 7335 14980 7380 15008
rect 7374 14968 7380 14980
rect 7432 15008 7438 15020
rect 8021 15011 8079 15017
rect 8021 15008 8033 15011
rect 7432 14980 8033 15008
rect 7432 14968 7438 14980
rect 8021 14977 8033 14980
rect 8067 14977 8079 15011
rect 8021 14971 8079 14977
rect 8110 14968 8116 15020
rect 8168 15008 8174 15020
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 8168 14980 8217 15008
rect 8168 14968 8174 14980
rect 8205 14977 8217 14980
rect 8251 15008 8263 15011
rect 8251 14980 8800 15008
rect 8251 14977 8263 14980
rect 8205 14971 8263 14977
rect 1486 14940 1492 14952
rect 1447 14912 1492 14940
rect 1486 14900 1492 14912
rect 1544 14900 1550 14952
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4249 14943 4307 14949
rect 4249 14940 4261 14943
rect 4120 14912 4261 14940
rect 4120 14900 4126 14912
rect 4249 14909 4261 14912
rect 4295 14940 4307 14943
rect 5258 14940 5264 14952
rect 4295 14912 5264 14940
rect 4295 14909 4307 14912
rect 4249 14903 4307 14909
rect 5258 14900 5264 14912
rect 5316 14900 5322 14952
rect 1756 14875 1814 14881
rect 1756 14841 1768 14875
rect 1802 14872 1814 14875
rect 1946 14872 1952 14884
rect 1802 14844 1952 14872
rect 1802 14841 1814 14844
rect 1756 14835 1814 14841
rect 1946 14832 1952 14844
rect 2004 14832 2010 14884
rect 4157 14875 4215 14881
rect 4157 14841 4169 14875
rect 4203 14872 4215 14875
rect 4516 14875 4574 14881
rect 4516 14872 4528 14875
rect 4203 14844 4528 14872
rect 4203 14841 4215 14844
rect 4157 14835 4215 14841
rect 4516 14841 4528 14844
rect 4562 14872 4574 14875
rect 4982 14872 4988 14884
rect 4562 14844 4988 14872
rect 4562 14841 4574 14844
rect 4516 14835 4574 14841
rect 4982 14832 4988 14844
rect 5040 14872 5046 14884
rect 6270 14872 6276 14884
rect 5040 14844 6276 14872
rect 5040 14832 5046 14844
rect 6270 14832 6276 14844
rect 6328 14832 6334 14884
rect 6641 14875 6699 14881
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 6730 14872 6736 14884
rect 6687 14844 6736 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 6730 14832 6736 14844
rect 6788 14832 6794 14884
rect 7742 14832 7748 14884
rect 7800 14872 7806 14884
rect 8573 14875 8631 14881
rect 8573 14872 8585 14875
rect 7800 14844 8585 14872
rect 7800 14832 7806 14844
rect 8573 14841 8585 14844
rect 8619 14841 8631 14875
rect 8772 14872 8800 14980
rect 9122 14940 9128 14952
rect 9083 14912 9128 14940
rect 9122 14900 9128 14912
rect 9180 14900 9186 14952
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13808 14943 13866 14949
rect 13808 14909 13820 14943
rect 13854 14940 13866 14943
rect 14274 14940 14280 14952
rect 13854 14912 14280 14940
rect 13854 14909 13866 14912
rect 13808 14903 13866 14909
rect 9398 14881 9404 14884
rect 9392 14872 9404 14881
rect 8772 14844 9404 14872
rect 8573 14835 8631 14841
rect 9392 14835 9404 14844
rect 9398 14832 9404 14835
rect 9456 14832 9462 14884
rect 11790 14832 11796 14884
rect 11848 14872 11854 14884
rect 11885 14875 11943 14881
rect 11885 14872 11897 14875
rect 11848 14844 11897 14872
rect 11848 14832 11854 14844
rect 11885 14841 11897 14844
rect 11931 14872 11943 14875
rect 12342 14872 12348 14884
rect 11931 14844 12348 14872
rect 11931 14841 11943 14844
rect 11885 14835 11943 14841
rect 12342 14832 12348 14844
rect 12400 14832 12406 14884
rect 12618 14832 12624 14884
rect 12676 14872 12682 14884
rect 13556 14872 13584 14903
rect 14274 14900 14280 14912
rect 14332 14900 14338 14952
rect 20990 14900 20996 14952
rect 21048 14940 21054 14952
rect 21637 14943 21695 14949
rect 21637 14940 21649 14943
rect 21048 14912 21649 14940
rect 21048 14900 21054 14912
rect 21637 14909 21649 14912
rect 21683 14940 21695 14943
rect 22189 14943 22247 14949
rect 22189 14940 22201 14943
rect 21683 14912 22201 14940
rect 21683 14909 21695 14912
rect 21637 14903 21695 14909
rect 22189 14909 22201 14912
rect 22235 14909 22247 14943
rect 22189 14903 22247 14909
rect 14366 14872 14372 14884
rect 12676 14844 14372 14872
rect 12676 14832 12682 14844
rect 14366 14832 14372 14844
rect 14424 14832 14430 14884
rect 2038 14764 2044 14816
rect 2096 14804 2102 14816
rect 2869 14807 2927 14813
rect 2869 14804 2881 14807
rect 2096 14776 2881 14804
rect 2096 14764 2102 14776
rect 2869 14773 2881 14776
rect 2915 14804 2927 14807
rect 3050 14804 3056 14816
rect 2915 14776 3056 14804
rect 2915 14773 2927 14776
rect 2869 14767 2927 14773
rect 3050 14764 3056 14776
rect 3108 14764 3114 14816
rect 3418 14804 3424 14816
rect 3379 14776 3424 14804
rect 3418 14764 3424 14776
rect 3476 14764 3482 14816
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 7929 14807 7987 14813
rect 7929 14804 7941 14807
rect 7524 14776 7941 14804
rect 7524 14764 7530 14776
rect 7929 14773 7941 14776
rect 7975 14773 7987 14807
rect 7929 14767 7987 14773
rect 12066 14764 12072 14816
rect 12124 14804 12130 14816
rect 12161 14807 12219 14813
rect 12161 14804 12173 14807
rect 12124 14776 12173 14804
rect 12124 14764 12130 14776
rect 12161 14773 12173 14776
rect 12207 14773 12219 14807
rect 12526 14804 12532 14816
rect 12487 14776 12532 14804
rect 12161 14767 12219 14773
rect 12526 14764 12532 14776
rect 12584 14764 12590 14816
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 13262 14804 13268 14816
rect 12860 14776 13268 14804
rect 12860 14764 12866 14776
rect 13262 14764 13268 14776
rect 13320 14804 13326 14816
rect 13357 14807 13415 14813
rect 13357 14804 13369 14807
rect 13320 14776 13369 14804
rect 13320 14764 13326 14776
rect 13357 14773 13369 14776
rect 13403 14773 13415 14807
rect 13357 14767 13415 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1397 14603 1455 14609
rect 1397 14569 1409 14603
rect 1443 14600 1455 14603
rect 1854 14600 1860 14612
rect 1443 14572 1860 14600
rect 1443 14569 1455 14572
rect 1397 14563 1455 14569
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 3510 14600 3516 14612
rect 3471 14572 3516 14600
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 4246 14560 4252 14612
rect 4304 14600 4310 14612
rect 4617 14603 4675 14609
rect 4617 14600 4629 14603
rect 4304 14572 4629 14600
rect 4304 14560 4310 14572
rect 4617 14569 4629 14572
rect 4663 14569 4675 14603
rect 4617 14563 4675 14569
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 8021 14603 8079 14609
rect 8021 14600 8033 14603
rect 7800 14572 8033 14600
rect 7800 14560 7806 14572
rect 8021 14569 8033 14572
rect 8067 14569 8079 14603
rect 8021 14563 8079 14569
rect 8202 14560 8208 14612
rect 8260 14600 8266 14612
rect 8481 14603 8539 14609
rect 8481 14600 8493 14603
rect 8260 14572 8493 14600
rect 8260 14560 8266 14572
rect 8481 14569 8493 14572
rect 8527 14600 8539 14603
rect 8846 14600 8852 14612
rect 8527 14572 8852 14600
rect 8527 14569 8539 14572
rect 8481 14563 8539 14569
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 9953 14603 10011 14609
rect 9953 14569 9965 14603
rect 9999 14600 10011 14603
rect 10042 14600 10048 14612
rect 9999 14572 10048 14600
rect 9999 14569 10011 14572
rect 9953 14563 10011 14569
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 11698 14560 11704 14612
rect 11756 14600 11762 14612
rect 12161 14603 12219 14609
rect 12161 14600 12173 14603
rect 11756 14572 12173 14600
rect 11756 14560 11762 14572
rect 12161 14569 12173 14572
rect 12207 14600 12219 14603
rect 12342 14600 12348 14612
rect 12207 14572 12348 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 12618 14600 12624 14612
rect 12579 14572 12624 14600
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13872 14572 14105 14600
rect 13872 14560 13878 14572
rect 14093 14569 14105 14572
rect 14139 14600 14151 14603
rect 14274 14600 14280 14612
rect 14139 14572 14280 14600
rect 14139 14569 14151 14572
rect 14093 14563 14151 14569
rect 14274 14560 14280 14572
rect 14332 14560 14338 14612
rect 14366 14560 14372 14612
rect 14424 14600 14430 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 14424 14572 14657 14600
rect 14424 14560 14430 14572
rect 14645 14569 14657 14572
rect 14691 14569 14703 14603
rect 14645 14563 14703 14569
rect 5258 14532 5264 14544
rect 5171 14504 5264 14532
rect 1765 14467 1823 14473
rect 1765 14433 1777 14467
rect 1811 14464 1823 14467
rect 2774 14464 2780 14476
rect 1811 14436 2780 14464
rect 1811 14433 1823 14436
rect 1765 14427 1823 14433
rect 2774 14424 2780 14436
rect 2832 14464 2838 14476
rect 2961 14467 3019 14473
rect 2961 14464 2973 14467
rect 2832 14436 2973 14464
rect 2832 14424 2838 14436
rect 2961 14433 2973 14436
rect 3007 14433 3019 14467
rect 2961 14427 3019 14433
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 5184 14473 5212 14504
rect 5258 14492 5264 14504
rect 5316 14532 5322 14544
rect 6730 14532 6736 14544
rect 5316 14504 6736 14532
rect 5316 14492 5322 14504
rect 6730 14492 6736 14504
rect 6788 14492 6794 14544
rect 8110 14492 8116 14544
rect 8168 14532 8174 14544
rect 8389 14535 8447 14541
rect 8389 14532 8401 14535
rect 8168 14504 8401 14532
rect 8168 14492 8174 14504
rect 8389 14501 8401 14504
rect 8435 14532 8447 14535
rect 9582 14532 9588 14544
rect 8435 14504 9588 14532
rect 8435 14501 8447 14504
rect 8389 14495 8447 14501
rect 9582 14492 9588 14504
rect 9640 14492 9646 14544
rect 10496 14535 10554 14541
rect 10496 14501 10508 14535
rect 10542 14532 10554 14535
rect 10686 14532 10692 14544
rect 10542 14504 10692 14532
rect 10542 14501 10554 14504
rect 10496 14495 10554 14501
rect 10686 14492 10692 14504
rect 10744 14492 10750 14544
rect 12066 14492 12072 14544
rect 12124 14532 12130 14544
rect 12124 14504 12940 14532
rect 12124 14492 12130 14504
rect 4065 14467 4123 14473
rect 4065 14464 4077 14467
rect 4028 14436 4077 14464
rect 4028 14424 4034 14436
rect 4065 14433 4077 14436
rect 4111 14433 4123 14467
rect 4065 14427 4123 14433
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14433 5227 14467
rect 5169 14427 5227 14433
rect 5436 14467 5494 14473
rect 5436 14433 5448 14467
rect 5482 14464 5494 14467
rect 5994 14464 6000 14476
rect 5482 14436 6000 14464
rect 5482 14433 5494 14436
rect 5436 14427 5494 14433
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 9122 14424 9128 14476
rect 9180 14464 9186 14476
rect 10229 14467 10287 14473
rect 10229 14464 10241 14467
rect 9180 14436 10241 14464
rect 9180 14424 9186 14436
rect 10229 14433 10241 14436
rect 10275 14464 10287 14467
rect 10962 14464 10968 14476
rect 10275 14436 10968 14464
rect 10275 14433 10287 14436
rect 10229 14427 10287 14433
rect 10962 14424 10968 14436
rect 11020 14424 11026 14476
rect 12250 14424 12256 14476
rect 12308 14464 12314 14476
rect 12618 14464 12624 14476
rect 12308 14436 12624 14464
rect 12308 14424 12314 14436
rect 12618 14424 12624 14436
rect 12676 14464 12682 14476
rect 12713 14467 12771 14473
rect 12713 14464 12725 14467
rect 12676 14436 12725 14464
rect 12676 14424 12682 14436
rect 12713 14433 12725 14436
rect 12759 14433 12771 14467
rect 12912 14464 12940 14504
rect 12980 14467 13038 14473
rect 12980 14464 12992 14467
rect 12912 14436 12992 14464
rect 12713 14427 12771 14433
rect 12980 14433 12992 14436
rect 13026 14464 13038 14467
rect 13354 14464 13360 14476
rect 13026 14436 13360 14464
rect 13026 14433 13038 14436
rect 12980 14427 13038 14433
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 1854 14396 1860 14408
rect 1815 14368 1860 14396
rect 1854 14356 1860 14368
rect 1912 14356 1918 14408
rect 1946 14356 1952 14408
rect 2004 14396 2010 14408
rect 2041 14399 2099 14405
rect 2041 14396 2053 14399
rect 2004 14368 2053 14396
rect 2004 14356 2010 14368
rect 2041 14365 2053 14368
rect 2087 14396 2099 14399
rect 3510 14396 3516 14408
rect 2087 14368 3516 14396
rect 2087 14365 2099 14368
rect 2041 14359 2099 14365
rect 3510 14356 3516 14368
rect 3568 14356 3574 14408
rect 8570 14356 8576 14408
rect 8628 14396 8634 14408
rect 8628 14368 8673 14396
rect 8628 14356 8634 14368
rect 1872 14328 1900 14356
rect 2409 14331 2467 14337
rect 2409 14328 2421 14331
rect 1872 14300 2421 14328
rect 2409 14297 2421 14300
rect 2455 14297 2467 14331
rect 2409 14291 2467 14297
rect 4249 14331 4307 14337
rect 4249 14297 4261 14331
rect 4295 14328 4307 14331
rect 4430 14328 4436 14340
rect 4295 14300 4436 14328
rect 4295 14297 4307 14300
rect 4249 14291 4307 14297
rect 4430 14288 4436 14300
rect 4488 14288 4494 14340
rect 6270 14288 6276 14340
rect 6328 14328 6334 14340
rect 6549 14331 6607 14337
rect 6549 14328 6561 14331
rect 6328 14300 6561 14328
rect 6328 14288 6334 14300
rect 6549 14297 6561 14300
rect 6595 14328 6607 14331
rect 6914 14328 6920 14340
rect 6595 14300 6920 14328
rect 6595 14297 6607 14300
rect 6549 14291 6607 14297
rect 6914 14288 6920 14300
rect 6972 14288 6978 14340
rect 2590 14220 2596 14272
rect 2648 14260 2654 14272
rect 2777 14263 2835 14269
rect 2777 14260 2789 14263
rect 2648 14232 2789 14260
rect 2648 14220 2654 14232
rect 2777 14229 2789 14232
rect 2823 14229 2835 14263
rect 2777 14223 2835 14229
rect 3602 14220 3608 14272
rect 3660 14260 3666 14272
rect 3789 14263 3847 14269
rect 3789 14260 3801 14263
rect 3660 14232 3801 14260
rect 3660 14220 3666 14232
rect 3789 14229 3801 14232
rect 3835 14229 3847 14263
rect 4982 14260 4988 14272
rect 4943 14232 4988 14260
rect 3789 14223 3847 14229
rect 4982 14220 4988 14232
rect 5040 14220 5046 14272
rect 7190 14260 7196 14272
rect 7151 14232 7196 14260
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 7466 14220 7472 14272
rect 7524 14260 7530 14272
rect 7561 14263 7619 14269
rect 7561 14260 7573 14263
rect 7524 14232 7573 14260
rect 7524 14220 7530 14232
rect 7561 14229 7573 14232
rect 7607 14229 7619 14263
rect 7561 14223 7619 14229
rect 9217 14263 9275 14269
rect 9217 14229 9229 14263
rect 9263 14260 9275 14263
rect 9398 14260 9404 14272
rect 9263 14232 9404 14260
rect 9263 14229 9275 14232
rect 9217 14223 9275 14229
rect 9398 14220 9404 14232
rect 9456 14260 9462 14272
rect 9582 14260 9588 14272
rect 9456 14232 9588 14260
rect 9456 14220 9462 14232
rect 9582 14220 9588 14232
rect 9640 14220 9646 14272
rect 11606 14260 11612 14272
rect 11567 14232 11612 14260
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 3510 14016 3516 14068
rect 3568 14056 3574 14068
rect 3605 14059 3663 14065
rect 3605 14056 3617 14059
rect 3568 14028 3617 14056
rect 3568 14016 3574 14028
rect 3605 14025 3617 14028
rect 3651 14025 3663 14059
rect 3970 14056 3976 14068
rect 3931 14028 3976 14056
rect 3605 14019 3663 14025
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 6822 14056 6828 14068
rect 6783 14028 6828 14056
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 7929 14059 7987 14065
rect 7929 14025 7941 14059
rect 7975 14056 7987 14059
rect 8570 14056 8576 14068
rect 7975 14028 8576 14056
rect 7975 14025 7987 14028
rect 7929 14019 7987 14025
rect 8570 14016 8576 14028
rect 8628 14016 8634 14068
rect 8754 14016 8760 14068
rect 8812 14056 8818 14068
rect 9677 14059 9735 14065
rect 9677 14056 9689 14059
rect 8812 14028 9689 14056
rect 8812 14016 8818 14028
rect 9677 14025 9689 14028
rect 9723 14025 9735 14059
rect 9677 14019 9735 14025
rect 10505 14059 10563 14065
rect 10505 14025 10517 14059
rect 10551 14056 10563 14059
rect 10686 14056 10692 14068
rect 10551 14028 10692 14056
rect 10551 14025 10563 14028
rect 10505 14019 10563 14025
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 11330 14056 11336 14068
rect 11291 14028 11336 14056
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 11664 14028 12173 14056
rect 11664 14016 11670 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 5169 13991 5227 13997
rect 5169 13957 5181 13991
rect 5215 13988 5227 13991
rect 11885 13991 11943 13997
rect 5215 13960 7236 13988
rect 5215 13957 5227 13960
rect 5169 13951 5227 13957
rect 7208 13932 7236 13960
rect 11885 13957 11897 13991
rect 11931 13988 11943 13991
rect 12066 13988 12072 14000
rect 11931 13960 12072 13988
rect 11931 13957 11943 13960
rect 11885 13951 11943 13957
rect 12066 13948 12072 13960
rect 12124 13948 12130 14000
rect 4890 13880 4896 13932
rect 4948 13920 4954 13932
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 4948 13892 5089 13920
rect 4948 13880 4954 13892
rect 5077 13889 5089 13892
rect 5123 13920 5135 13923
rect 5442 13920 5448 13932
rect 5123 13892 5448 13920
rect 5123 13889 5135 13892
rect 5077 13883 5135 13889
rect 5442 13880 5448 13892
rect 5500 13920 5506 13932
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 5500 13892 5641 13920
rect 5500 13880 5506 13892
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13920 5871 13923
rect 5994 13920 6000 13932
rect 5859 13892 6000 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 5994 13880 6000 13892
rect 6052 13880 6058 13932
rect 7190 13880 7196 13932
rect 7248 13920 7254 13932
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 7248 13892 7297 13920
rect 7248 13880 7254 13892
rect 7285 13889 7297 13892
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13889 7435 13923
rect 12176 13920 12204 14019
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 13817 14059 13875 14065
rect 13817 14056 13829 14059
rect 13412 14028 13829 14056
rect 13412 14016 13418 14028
rect 13817 14025 13829 14028
rect 13863 14025 13875 14059
rect 13817 14019 13875 14025
rect 16390 13920 16396 13932
rect 12176 13892 12572 13920
rect 16351 13892 16396 13920
rect 7377 13883 7435 13889
rect 1486 13812 1492 13864
rect 1544 13852 1550 13864
rect 1673 13855 1731 13861
rect 1673 13852 1685 13855
rect 1544 13824 1685 13852
rect 1544 13812 1550 13824
rect 1673 13821 1685 13824
rect 1719 13852 1731 13855
rect 1762 13852 1768 13864
rect 1719 13824 1768 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 1940 13855 1998 13861
rect 1940 13821 1952 13855
rect 1986 13852 1998 13855
rect 3050 13852 3056 13864
rect 1986 13824 3056 13852
rect 1986 13821 1998 13824
rect 1940 13815 1998 13821
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 4709 13855 4767 13861
rect 4709 13821 4721 13855
rect 4755 13852 4767 13855
rect 4755 13824 5488 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 4154 13784 4160 13796
rect 4115 13756 4160 13784
rect 4154 13744 4160 13756
rect 4212 13744 4218 13796
rect 5460 13784 5488 13824
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 7392 13852 7420 13883
rect 6972 13824 7420 13852
rect 8297 13855 8355 13861
rect 6972 13812 6978 13824
rect 8297 13821 8309 13855
rect 8343 13852 8355 13855
rect 8386 13852 8392 13864
rect 8343 13824 8392 13852
rect 8343 13821 8355 13824
rect 8297 13815 8355 13821
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 12437 13855 12495 13861
rect 12437 13821 12449 13855
rect 12483 13821 12495 13855
rect 12544 13852 12572 13892
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 20990 13920 20996 13932
rect 20951 13892 20996 13920
rect 20990 13880 20996 13892
rect 21048 13880 21054 13932
rect 12693 13855 12751 13861
rect 12693 13852 12705 13855
rect 12544 13824 12705 13852
rect 12437 13815 12495 13821
rect 12693 13821 12705 13824
rect 12739 13821 12751 13855
rect 16114 13852 16120 13864
rect 16075 13824 16120 13852
rect 12693 13815 12751 13821
rect 5537 13787 5595 13793
rect 5537 13784 5549 13787
rect 5460 13756 5549 13784
rect 5537 13753 5549 13756
rect 5583 13784 5595 13787
rect 6454 13784 6460 13796
rect 5583 13756 6460 13784
rect 5583 13753 5595 13756
rect 5537 13747 5595 13753
rect 6454 13744 6460 13756
rect 6512 13744 6518 13796
rect 10870 13784 10876 13796
rect 10831 13756 10876 13784
rect 10870 13744 10876 13756
rect 10928 13744 10934 13796
rect 12452 13784 12480 13815
rect 16114 13812 16120 13824
rect 16172 13852 16178 13864
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 16172 13824 16865 13852
rect 16172 13812 16178 13824
rect 16853 13821 16865 13824
rect 16899 13821 16911 13855
rect 20714 13852 20720 13864
rect 20675 13824 20720 13852
rect 16853 13815 16911 13821
rect 20714 13812 20720 13824
rect 20772 13852 20778 13864
rect 21453 13855 21511 13861
rect 21453 13852 21465 13855
rect 20772 13824 21465 13852
rect 20772 13812 20778 13824
rect 21453 13821 21465 13824
rect 21499 13821 21511 13855
rect 21453 13815 21511 13821
rect 12452 13756 12664 13784
rect 12636 13728 12664 13756
rect 2314 13676 2320 13728
rect 2372 13716 2378 13728
rect 3053 13719 3111 13725
rect 3053 13716 3065 13719
rect 2372 13688 3065 13716
rect 2372 13676 2378 13688
rect 3053 13685 3065 13688
rect 3099 13685 3111 13719
rect 3053 13679 3111 13685
rect 5994 13676 6000 13728
rect 6052 13716 6058 13728
rect 6181 13719 6239 13725
rect 6181 13716 6193 13719
rect 6052 13688 6193 13716
rect 6052 13676 6058 13688
rect 6181 13685 6193 13688
rect 6227 13716 6239 13719
rect 6549 13719 6607 13725
rect 6549 13716 6561 13719
rect 6227 13688 6561 13716
rect 6227 13685 6239 13688
rect 6181 13679 6239 13685
rect 6549 13685 6561 13688
rect 6595 13685 6607 13719
rect 7190 13716 7196 13728
rect 7151 13688 7196 13716
rect 6549 13679 6607 13685
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 12618 13676 12624 13728
rect 12676 13676 12682 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2774 13512 2780 13524
rect 2735 13484 2780 13512
rect 2774 13472 2780 13484
rect 2832 13472 2838 13524
rect 3050 13512 3056 13524
rect 3011 13484 3056 13512
rect 3050 13472 3056 13484
rect 3108 13472 3114 13524
rect 3421 13515 3479 13521
rect 3421 13481 3433 13515
rect 3467 13512 3479 13515
rect 3878 13512 3884 13524
rect 3467 13484 3884 13512
rect 3467 13481 3479 13484
rect 3421 13475 3479 13481
rect 3878 13472 3884 13484
rect 3936 13512 3942 13524
rect 4062 13512 4068 13524
rect 3936 13484 4068 13512
rect 3936 13472 3942 13484
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 5721 13515 5779 13521
rect 5721 13481 5733 13515
rect 5767 13512 5779 13515
rect 6362 13512 6368 13524
rect 5767 13484 6368 13512
rect 5767 13481 5779 13484
rect 5721 13475 5779 13481
rect 6362 13472 6368 13484
rect 6420 13472 6426 13524
rect 7190 13512 7196 13524
rect 6472 13484 7196 13512
rect 4706 13404 4712 13456
rect 4764 13444 4770 13456
rect 5629 13447 5687 13453
rect 5629 13444 5641 13447
rect 4764 13416 5641 13444
rect 4764 13404 4770 13416
rect 5629 13413 5641 13416
rect 5675 13444 5687 13447
rect 6086 13444 6092 13456
rect 5675 13416 6092 13444
rect 5675 13413 5687 13416
rect 5629 13407 5687 13413
rect 6086 13404 6092 13416
rect 6144 13404 6150 13456
rect 1670 13336 1676 13388
rect 1728 13376 1734 13388
rect 2041 13379 2099 13385
rect 2041 13376 2053 13379
rect 1728 13348 2053 13376
rect 1728 13336 1734 13348
rect 2041 13345 2053 13348
rect 2087 13345 2099 13379
rect 3602 13376 3608 13388
rect 3563 13348 3608 13376
rect 2041 13339 2099 13345
rect 3602 13336 3608 13348
rect 3660 13336 3666 13388
rect 2130 13308 2136 13320
rect 2091 13280 2136 13308
rect 2130 13268 2136 13280
rect 2188 13268 2194 13320
rect 2314 13308 2320 13320
rect 2275 13280 2320 13308
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13308 4123 13311
rect 4801 13311 4859 13317
rect 4801 13308 4813 13311
rect 4111 13280 4813 13308
rect 4111 13277 4123 13280
rect 4065 13271 4123 13277
rect 4801 13277 4813 13280
rect 4847 13308 4859 13311
rect 5166 13308 5172 13320
rect 4847 13280 5172 13308
rect 4847 13277 4859 13280
rect 4801 13271 4859 13277
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13308 5963 13311
rect 5994 13308 6000 13320
rect 5951 13280 6000 13308
rect 5951 13277 5963 13280
rect 5905 13271 5963 13277
rect 5994 13268 6000 13280
rect 6052 13268 6058 13320
rect 6472 13249 6500 13484
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7929 13515 7987 13521
rect 7929 13481 7941 13515
rect 7975 13512 7987 13515
rect 8202 13512 8208 13524
rect 7975 13484 8208 13512
rect 7975 13481 7987 13484
rect 7929 13475 7987 13481
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 10134 13512 10140 13524
rect 10095 13484 10140 13512
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12894 13512 12900 13524
rect 12492 13484 12537 13512
rect 12855 13484 12900 13512
rect 12492 13472 12498 13484
rect 12894 13472 12900 13484
rect 12952 13472 12958 13524
rect 6914 13404 6920 13456
rect 6972 13444 6978 13456
rect 7561 13447 7619 13453
rect 6972 13416 7017 13444
rect 6972 13404 6978 13416
rect 7561 13413 7573 13447
rect 7607 13444 7619 13447
rect 8110 13444 8116 13456
rect 7607 13416 8116 13444
rect 7607 13413 7619 13416
rect 7561 13407 7619 13413
rect 8110 13404 8116 13416
rect 8168 13404 8174 13456
rect 9493 13447 9551 13453
rect 9493 13413 9505 13447
rect 9539 13444 9551 13447
rect 9582 13444 9588 13456
rect 9539 13416 9588 13444
rect 9539 13413 9551 13416
rect 9493 13407 9551 13413
rect 9582 13404 9588 13416
rect 9640 13444 9646 13456
rect 9640 13416 10272 13444
rect 9640 13404 9646 13416
rect 8389 13379 8447 13385
rect 8389 13376 8401 13379
rect 7944 13348 8401 13376
rect 7944 13320 7972 13348
rect 8389 13345 8401 13348
rect 8435 13345 8447 13379
rect 10042 13376 10048 13388
rect 10003 13348 10048 13376
rect 8389 13339 8447 13345
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13308 7067 13311
rect 7926 13308 7932 13320
rect 7055 13280 7932 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 7926 13268 7932 13280
rect 7984 13268 7990 13320
rect 8478 13308 8484 13320
rect 8439 13280 8484 13308
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 10244 13317 10272 13416
rect 12618 13404 12624 13456
rect 12676 13444 12682 13456
rect 13449 13447 13507 13453
rect 13449 13444 13461 13447
rect 12676 13416 13461 13444
rect 12676 13404 12682 13416
rect 13449 13413 13461 13416
rect 13495 13413 13507 13447
rect 13449 13407 13507 13413
rect 17586 13404 17592 13456
rect 17644 13444 17650 13456
rect 17681 13447 17739 13453
rect 17681 13444 17693 13447
rect 17644 13416 17693 13444
rect 17644 13404 17650 13416
rect 17681 13413 17693 13416
rect 17727 13413 17739 13447
rect 17681 13407 17739 13413
rect 11882 13336 11888 13388
rect 11940 13376 11946 13388
rect 12158 13376 12164 13388
rect 11940 13348 12164 13376
rect 11940 13336 11946 13348
rect 12158 13336 12164 13348
rect 12216 13376 12222 13388
rect 12805 13379 12863 13385
rect 12805 13376 12817 13379
rect 12216 13348 12817 13376
rect 12216 13336 12222 13348
rect 12805 13345 12817 13348
rect 12851 13345 12863 13379
rect 17402 13376 17408 13388
rect 17363 13348 17408 13376
rect 12805 13339 12863 13345
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 10229 13311 10287 13317
rect 8711 13280 9168 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 5261 13243 5319 13249
rect 5261 13209 5273 13243
rect 5307 13240 5319 13243
rect 6457 13243 6515 13249
rect 6457 13240 6469 13243
rect 5307 13212 6469 13240
rect 5307 13209 5319 13212
rect 5261 13203 5319 13209
rect 6457 13209 6469 13212
rect 6503 13209 6515 13243
rect 8018 13240 8024 13252
rect 7979 13212 8024 13240
rect 6457 13203 6515 13209
rect 8018 13200 8024 13212
rect 8076 13200 8082 13252
rect 1673 13175 1731 13181
rect 1673 13141 1685 13175
rect 1719 13172 1731 13175
rect 2682 13172 2688 13184
rect 1719 13144 2688 13172
rect 1719 13141 1731 13144
rect 1673 13135 1731 13141
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 9140 13181 9168 13280
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13308 13139 13311
rect 13722 13308 13728 13320
rect 13127 13280 13728 13308
rect 13127 13277 13139 13280
rect 13081 13271 13139 13277
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 9677 13243 9735 13249
rect 9677 13209 9689 13243
rect 9723 13240 9735 13243
rect 10870 13240 10876 13252
rect 9723 13212 10876 13240
rect 9723 13209 9735 13212
rect 9677 13203 9735 13209
rect 10870 13200 10876 13212
rect 10928 13240 10934 13252
rect 11057 13243 11115 13249
rect 11057 13240 11069 13243
rect 10928 13212 11069 13240
rect 10928 13200 10934 13212
rect 11057 13209 11069 13212
rect 11103 13209 11115 13243
rect 11057 13203 11115 13209
rect 11885 13243 11943 13249
rect 11885 13209 11897 13243
rect 11931 13240 11943 13243
rect 12618 13240 12624 13252
rect 11931 13212 12624 13240
rect 11931 13209 11943 13212
rect 11885 13203 11943 13209
rect 12618 13200 12624 13212
rect 12676 13200 12682 13252
rect 9125 13175 9183 13181
rect 9125 13141 9137 13175
rect 9171 13172 9183 13175
rect 9214 13172 9220 13184
rect 9171 13144 9220 13172
rect 9171 13141 9183 13144
rect 9125 13135 9183 13141
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 10781 13175 10839 13181
rect 10781 13141 10793 13175
rect 10827 13172 10839 13175
rect 10962 13172 10968 13184
rect 10827 13144 10968 13172
rect 10827 13141 10839 13144
rect 10781 13135 10839 13141
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 11422 13172 11428 13184
rect 11383 13144 11428 13172
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1670 12968 1676 12980
rect 1631 12940 1676 12968
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 2130 12968 2136 12980
rect 2091 12940 2136 12968
rect 2130 12928 2136 12940
rect 2188 12928 2194 12980
rect 3878 12968 3884 12980
rect 2332 12940 3884 12968
rect 1762 12860 1768 12912
rect 1820 12900 1826 12912
rect 2332 12900 2360 12940
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 4798 12968 4804 12980
rect 4759 12940 4804 12968
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 6362 12968 6368 12980
rect 5951 12940 6368 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 6362 12928 6368 12940
rect 6420 12928 6426 12980
rect 7926 12968 7932 12980
rect 7887 12940 7932 12968
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 9769 12971 9827 12977
rect 9769 12968 9781 12971
rect 9732 12940 9781 12968
rect 9732 12928 9738 12940
rect 9769 12937 9781 12940
rect 9815 12937 9827 12971
rect 9769 12931 9827 12937
rect 10134 12928 10140 12980
rect 10192 12968 10198 12980
rect 11425 12971 11483 12977
rect 11425 12968 11437 12971
rect 10192 12940 11437 12968
rect 10192 12928 10198 12940
rect 11425 12937 11437 12940
rect 11471 12937 11483 12971
rect 11882 12968 11888 12980
rect 11843 12940 11888 12968
rect 11425 12931 11483 12937
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12492 12940 12537 12968
rect 12492 12928 12498 12940
rect 12894 12928 12900 12980
rect 12952 12968 12958 12980
rect 13817 12971 13875 12977
rect 13817 12968 13829 12971
rect 12952 12940 13829 12968
rect 12952 12928 12958 12940
rect 13817 12937 13829 12940
rect 13863 12937 13875 12971
rect 13817 12931 13875 12937
rect 15473 12971 15531 12977
rect 15473 12937 15485 12971
rect 15519 12968 15531 12971
rect 16206 12968 16212 12980
rect 15519 12940 16212 12968
rect 15519 12937 15531 12940
rect 15473 12931 15531 12937
rect 16206 12928 16212 12940
rect 16264 12928 16270 12980
rect 4706 12900 4712 12912
rect 1820 12872 2360 12900
rect 4667 12872 4712 12900
rect 1820 12860 1826 12872
rect 2332 12841 2360 12872
rect 4706 12860 4712 12872
rect 4764 12860 4770 12912
rect 6549 12903 6607 12909
rect 6549 12900 6561 12903
rect 5276 12872 6561 12900
rect 5276 12844 5304 12872
rect 6549 12869 6561 12872
rect 6595 12869 6607 12903
rect 10410 12900 10416 12912
rect 10371 12872 10416 12900
rect 6549 12863 6607 12869
rect 10410 12860 10416 12872
rect 10468 12860 10474 12912
rect 13541 12903 13599 12909
rect 13541 12869 13553 12903
rect 13587 12900 13599 12903
rect 13722 12900 13728 12912
rect 13587 12872 13728 12900
rect 13587 12869 13599 12872
rect 13541 12863 13599 12869
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12801 2375 12835
rect 5258 12832 5264 12844
rect 5219 12804 5264 12832
rect 2317 12795 2375 12801
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12801 5411 12835
rect 5353 12795 5411 12801
rect 2406 12724 2412 12776
rect 2464 12764 2470 12776
rect 2573 12767 2631 12773
rect 2573 12764 2585 12767
rect 2464 12736 2585 12764
rect 2464 12724 2470 12736
rect 2573 12733 2585 12736
rect 2619 12733 2631 12767
rect 5166 12764 5172 12776
rect 5127 12736 5172 12764
rect 2573 12727 2631 12733
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 4341 12699 4399 12705
rect 4341 12696 4353 12699
rect 3712 12668 4353 12696
rect 3712 12637 3740 12668
rect 4341 12665 4353 12668
rect 4387 12696 4399 12699
rect 4706 12696 4712 12708
rect 4387 12668 4712 12696
rect 4387 12665 4399 12668
rect 4341 12659 4399 12665
rect 4706 12656 4712 12668
rect 4764 12696 4770 12708
rect 5368 12696 5396 12795
rect 7834 12792 7840 12844
rect 7892 12832 7898 12844
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 7892 12804 8401 12832
rect 7892 12792 7898 12804
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 10870 12832 10876 12844
rect 10831 12804 10876 12832
rect 8389 12795 8447 12801
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 10962 12792 10968 12844
rect 11020 12832 11026 12844
rect 12897 12835 12955 12841
rect 12897 12832 12909 12835
rect 11020 12804 11065 12832
rect 12176 12804 12909 12832
rect 11020 12792 11026 12804
rect 12176 12776 12204 12804
rect 12897 12801 12909 12804
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12832 13047 12835
rect 13078 12832 13084 12844
rect 13035 12804 13084 12832
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 13078 12792 13084 12804
rect 13136 12832 13142 12844
rect 13556 12832 13584 12863
rect 13722 12860 13728 12872
rect 13780 12860 13786 12912
rect 16758 12860 16764 12912
rect 16816 12900 16822 12912
rect 17402 12900 17408 12912
rect 16816 12872 17408 12900
rect 16816 12860 16822 12872
rect 17402 12860 17408 12872
rect 17460 12900 17466 12912
rect 17773 12903 17831 12909
rect 17773 12900 17785 12903
rect 17460 12872 17785 12900
rect 17460 12860 17466 12872
rect 17773 12869 17785 12872
rect 17819 12869 17831 12903
rect 17773 12863 17831 12869
rect 13136 12804 13584 12832
rect 14277 12835 14335 12841
rect 13136 12792 13142 12804
rect 14277 12801 14289 12835
rect 14323 12832 14335 12835
rect 16942 12832 16948 12844
rect 14323 12804 15332 12832
rect 16903 12804 16948 12832
rect 14323 12801 14335 12804
rect 14277 12795 14335 12801
rect 8294 12764 8300 12776
rect 8255 12736 8300 12764
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 12158 12764 12164 12776
rect 12119 12736 12164 12764
rect 12158 12724 12164 12736
rect 12216 12724 12222 12776
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12584 12736 12817 12764
rect 12584 12724 12590 12736
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 13998 12764 14004 12776
rect 13911 12736 14004 12764
rect 12805 12727 12863 12733
rect 13998 12724 14004 12736
rect 14056 12764 14062 12776
rect 15304 12773 15332 12804
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 18322 12832 18328 12844
rect 18283 12804 18328 12832
rect 18322 12792 18328 12804
rect 18380 12792 18386 12844
rect 14737 12767 14795 12773
rect 14737 12764 14749 12767
rect 14056 12736 14749 12764
rect 14056 12724 14062 12736
rect 14737 12733 14749 12736
rect 14783 12733 14795 12767
rect 14737 12727 14795 12733
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12764 15347 12767
rect 15841 12767 15899 12773
rect 15841 12764 15853 12767
rect 15335 12736 15853 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 15841 12733 15853 12736
rect 15887 12733 15899 12767
rect 16666 12764 16672 12776
rect 16579 12736 16672 12764
rect 15841 12727 15899 12733
rect 16666 12724 16672 12736
rect 16724 12764 16730 12776
rect 17405 12767 17463 12773
rect 17405 12764 17417 12767
rect 16724 12736 17417 12764
rect 16724 12724 16730 12736
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 18046 12764 18052 12776
rect 18007 12736 18052 12764
rect 17405 12727 17463 12733
rect 18046 12724 18052 12736
rect 18104 12764 18110 12776
rect 18785 12767 18843 12773
rect 18785 12764 18797 12767
rect 18104 12736 18797 12764
rect 18104 12724 18110 12736
rect 18785 12733 18797 12736
rect 18831 12733 18843 12767
rect 18785 12727 18843 12733
rect 4764 12668 5396 12696
rect 4764 12656 4770 12668
rect 5534 12656 5540 12708
rect 5592 12696 5598 12708
rect 5994 12696 6000 12708
rect 5592 12668 6000 12696
rect 5592 12656 5598 12668
rect 5994 12656 6000 12668
rect 6052 12696 6058 12708
rect 6181 12699 6239 12705
rect 6181 12696 6193 12699
rect 6052 12668 6193 12696
rect 6052 12656 6058 12668
rect 6181 12665 6193 12668
rect 6227 12665 6239 12699
rect 6181 12659 6239 12665
rect 7653 12699 7711 12705
rect 7653 12665 7665 12699
rect 7699 12696 7711 12699
rect 8656 12699 8714 12705
rect 8656 12696 8668 12699
rect 7699 12668 8668 12696
rect 7699 12665 7711 12668
rect 7653 12659 7711 12665
rect 8656 12665 8668 12668
rect 8702 12696 8714 12699
rect 9214 12696 9220 12708
rect 8702 12668 9220 12696
rect 8702 12665 8714 12668
rect 8656 12659 8714 12665
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 3697 12631 3755 12637
rect 3697 12597 3709 12631
rect 3743 12597 3755 12631
rect 6822 12628 6828 12640
rect 6783 12600 6828 12628
rect 3697 12591 3755 12597
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7834 12588 7840 12640
rect 7892 12628 7898 12640
rect 8113 12631 8171 12637
rect 8113 12628 8125 12631
rect 7892 12600 8125 12628
rect 7892 12588 7898 12600
rect 8113 12597 8125 12600
rect 8159 12597 8171 12631
rect 10778 12628 10784 12640
rect 10739 12600 10784 12628
rect 8113 12591 8171 12597
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1673 12427 1731 12433
rect 1673 12393 1685 12427
rect 1719 12424 1731 12427
rect 2406 12424 2412 12436
rect 1719 12396 2412 12424
rect 1719 12393 1731 12396
rect 1673 12387 1731 12393
rect 2406 12384 2412 12396
rect 2464 12424 2470 12436
rect 2777 12427 2835 12433
rect 2777 12424 2789 12427
rect 2464 12396 2789 12424
rect 2464 12384 2470 12396
rect 2777 12393 2789 12396
rect 2823 12393 2835 12427
rect 2777 12387 2835 12393
rect 7009 12427 7067 12433
rect 7009 12393 7021 12427
rect 7055 12393 7067 12427
rect 7466 12424 7472 12436
rect 7427 12396 7472 12424
rect 7009 12387 7067 12393
rect 6546 12356 6552 12368
rect 6507 12328 6552 12356
rect 6546 12316 6552 12328
rect 6604 12316 6610 12368
rect 6914 12356 6920 12368
rect 6656 12328 6920 12356
rect 1946 12248 1952 12300
rect 2004 12288 2010 12300
rect 2133 12291 2191 12297
rect 2133 12288 2145 12291
rect 2004 12260 2145 12288
rect 2004 12248 2010 12260
rect 2133 12257 2145 12260
rect 2179 12288 2191 12291
rect 3513 12291 3571 12297
rect 3513 12288 3525 12291
rect 2179 12260 3525 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 3513 12257 3525 12260
rect 3559 12257 3571 12291
rect 3513 12251 3571 12257
rect 3878 12248 3884 12300
rect 3936 12288 3942 12300
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 3936 12260 4077 12288
rect 3936 12248 3942 12260
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 4065 12251 4123 12257
rect 4332 12291 4390 12297
rect 4332 12257 4344 12291
rect 4378 12288 4390 12291
rect 4706 12288 4712 12300
rect 4378 12260 4712 12288
rect 4378 12257 4390 12260
rect 4332 12251 4390 12257
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 5994 12248 6000 12300
rect 6052 12288 6058 12300
rect 6656 12288 6684 12328
rect 6914 12316 6920 12328
rect 6972 12316 6978 12368
rect 7024 12356 7052 12387
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 9214 12424 9220 12436
rect 9175 12396 9220 12424
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 9769 12427 9827 12433
rect 9769 12393 9781 12427
rect 9815 12424 9827 12427
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 9815 12396 10701 12424
rect 9815 12393 9827 12396
rect 9769 12387 9827 12393
rect 10689 12393 10701 12396
rect 10735 12424 10747 12427
rect 10778 12424 10784 12436
rect 10735 12396 10784 12424
rect 10735 12393 10747 12396
rect 10689 12387 10747 12393
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12713 12427 12771 12433
rect 12713 12424 12725 12427
rect 12584 12396 12725 12424
rect 12584 12384 12590 12396
rect 12713 12393 12725 12396
rect 12759 12393 12771 12427
rect 13078 12424 13084 12436
rect 13039 12396 13084 12424
rect 12713 12387 12771 12393
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 13262 12424 13268 12436
rect 13223 12396 13268 12424
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 8478 12356 8484 12368
rect 7024 12328 8484 12356
rect 8478 12316 8484 12328
rect 8536 12316 8542 12368
rect 10962 12316 10968 12368
rect 11020 12365 11026 12368
rect 11020 12359 11084 12365
rect 11020 12325 11038 12359
rect 11072 12325 11084 12359
rect 11020 12319 11084 12325
rect 11020 12316 11026 12319
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 6052 12260 6684 12288
rect 6748 12260 7389 12288
rect 6052 12248 6058 12260
rect 1670 12180 1676 12232
rect 1728 12220 1734 12232
rect 2225 12223 2283 12229
rect 2225 12220 2237 12223
rect 1728 12192 2237 12220
rect 1728 12180 1734 12192
rect 2225 12189 2237 12192
rect 2271 12189 2283 12223
rect 2406 12220 2412 12232
rect 2367 12192 2412 12220
rect 2225 12183 2283 12189
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 6546 12180 6552 12232
rect 6604 12220 6610 12232
rect 6748 12220 6776 12260
rect 7377 12257 7389 12260
rect 7423 12257 7435 12291
rect 8104 12291 8162 12297
rect 8104 12288 8116 12291
rect 7377 12251 7435 12257
rect 7576 12260 8116 12288
rect 7576 12229 7604 12260
rect 8104 12257 8116 12260
rect 8150 12288 8162 12291
rect 9030 12288 9036 12300
rect 8150 12260 9036 12288
rect 8150 12257 8162 12260
rect 8104 12251 8162 12257
rect 9030 12248 9036 12260
rect 9088 12248 9094 12300
rect 11422 12288 11428 12300
rect 10796 12260 11428 12288
rect 10796 12232 10824 12260
rect 11422 12248 11428 12260
rect 11480 12248 11486 12300
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 14366 12288 14372 12300
rect 13679 12260 14372 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 14366 12248 14372 12260
rect 14424 12248 14430 12300
rect 6604 12192 6776 12220
rect 7561 12223 7619 12229
rect 6604 12180 6610 12192
rect 7561 12189 7573 12223
rect 7607 12189 7619 12223
rect 7834 12220 7840 12232
rect 7795 12192 7840 12220
rect 7561 12183 7619 12189
rect 1762 12152 1768 12164
rect 1723 12124 1768 12152
rect 1762 12112 1768 12124
rect 1820 12112 1826 12164
rect 6270 12112 6276 12164
rect 6328 12152 6334 12164
rect 7576 12152 7604 12183
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 10778 12220 10784 12232
rect 9180 12192 10784 12220
rect 9180 12180 9186 12192
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 12434 12220 12440 12232
rect 11940 12192 12440 12220
rect 11940 12180 11946 12192
rect 12434 12180 12440 12192
rect 12492 12220 12498 12232
rect 13725 12223 13783 12229
rect 13725 12220 13737 12223
rect 12492 12192 13737 12220
rect 12492 12180 12498 12192
rect 13725 12189 13737 12192
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 13872 12192 13917 12220
rect 13872 12180 13878 12192
rect 6328 12124 7604 12152
rect 6328 12112 6334 12124
rect 3142 12084 3148 12096
rect 3103 12056 3148 12084
rect 3142 12044 3148 12056
rect 3200 12044 3206 12096
rect 5442 12084 5448 12096
rect 5403 12056 5448 12084
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 5994 12084 6000 12096
rect 5955 12056 6000 12084
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 6972 12056 7017 12084
rect 6972 12044 6978 12056
rect 10134 12044 10140 12096
rect 10192 12084 10198 12096
rect 10229 12087 10287 12093
rect 10229 12084 10241 12087
rect 10192 12056 10241 12084
rect 10192 12044 10198 12056
rect 10229 12053 10241 12056
rect 10275 12053 10287 12087
rect 12158 12084 12164 12096
rect 12119 12056 12164 12084
rect 10229 12047 10287 12053
rect 12158 12044 12164 12056
rect 12216 12044 12222 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 2685 11883 2743 11889
rect 2685 11880 2697 11883
rect 2464 11852 2697 11880
rect 2464 11840 2470 11852
rect 2685 11849 2697 11852
rect 2731 11880 2743 11883
rect 3234 11880 3240 11892
rect 2731 11852 3240 11880
rect 2731 11849 2743 11852
rect 2685 11843 2743 11849
rect 3234 11840 3240 11852
rect 3292 11880 3298 11892
rect 3513 11883 3571 11889
rect 3513 11880 3525 11883
rect 3292 11852 3525 11880
rect 3292 11840 3298 11852
rect 3513 11849 3525 11852
rect 3559 11849 3571 11883
rect 5350 11880 5356 11892
rect 5311 11852 5356 11880
rect 3513 11843 3571 11849
rect 2222 11744 2228 11756
rect 2183 11716 2228 11744
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 3528 11744 3556 11843
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 6270 11880 6276 11892
rect 6231 11852 6276 11880
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 7834 11880 7840 11892
rect 6840 11852 7840 11880
rect 6840 11753 6868 11852
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 10689 11883 10747 11889
rect 10689 11849 10701 11883
rect 10735 11880 10747 11883
rect 10962 11880 10968 11892
rect 10735 11852 10968 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 10962 11840 10968 11852
rect 11020 11880 11026 11892
rect 11241 11883 11299 11889
rect 11241 11880 11253 11883
rect 11020 11852 11253 11880
rect 11020 11840 11026 11852
rect 11241 11849 11253 11852
rect 11287 11849 11299 11883
rect 11882 11880 11888 11892
rect 11843 11852 11888 11880
rect 11241 11843 11299 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12158 11880 12164 11892
rect 12119 11852 12164 11880
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 14366 11880 14372 11892
rect 14327 11852 14372 11880
rect 14366 11840 14372 11852
rect 14424 11880 14430 11892
rect 14424 11852 14964 11880
rect 14424 11840 14430 11852
rect 8205 11815 8263 11821
rect 8205 11781 8217 11815
rect 8251 11781 8263 11815
rect 8205 11775 8263 11781
rect 6825 11747 6883 11753
rect 3528 11716 4108 11744
rect 2041 11679 2099 11685
rect 2041 11645 2053 11679
rect 2087 11676 2099 11679
rect 2314 11676 2320 11688
rect 2087 11648 2320 11676
rect 2087 11645 2099 11648
rect 2041 11639 2099 11645
rect 2314 11636 2320 11648
rect 2372 11676 2378 11688
rect 3142 11676 3148 11688
rect 2372 11648 3148 11676
rect 2372 11636 2378 11648
rect 3142 11636 3148 11648
rect 3200 11636 3206 11688
rect 3878 11676 3884 11688
rect 3839 11648 3884 11676
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11645 4031 11679
rect 4080 11676 4108 11716
rect 6825 11713 6837 11747
rect 6871 11713 6883 11747
rect 8220 11744 8248 11775
rect 9217 11747 9275 11753
rect 9217 11744 9229 11747
rect 8220 11716 9229 11744
rect 6825 11707 6883 11713
rect 9217 11713 9229 11716
rect 9263 11744 9275 11747
rect 12176 11744 12204 11840
rect 14936 11753 14964 11852
rect 14921 11747 14979 11753
rect 9263 11716 9444 11744
rect 12176 11716 12572 11744
rect 9263 11713 9275 11716
rect 9217 11707 9275 11713
rect 4229 11679 4287 11685
rect 4229 11676 4241 11679
rect 4080 11648 4241 11676
rect 3973 11639 4031 11645
rect 4229 11645 4241 11648
rect 4275 11645 4287 11679
rect 4229 11639 4287 11645
rect 3988 11608 4016 11639
rect 6914 11636 6920 11688
rect 6972 11676 6978 11688
rect 7081 11679 7139 11685
rect 7081 11676 7093 11679
rect 6972 11648 7093 11676
rect 6972 11636 6978 11648
rect 7081 11645 7093 11648
rect 7127 11645 7139 11679
rect 7081 11639 7139 11645
rect 7834 11636 7840 11688
rect 7892 11676 7898 11688
rect 9122 11676 9128 11688
rect 7892 11648 9128 11676
rect 7892 11636 7898 11648
rect 9122 11636 9128 11648
rect 9180 11676 9186 11688
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 9180 11648 9321 11676
rect 9180 11636 9186 11648
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9416 11676 9444 11716
rect 12544 11688 12572 11716
rect 14921 11713 14933 11747
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 9582 11685 9588 11688
rect 9576 11676 9588 11685
rect 9416 11648 9588 11676
rect 9309 11639 9367 11645
rect 9576 11639 9588 11648
rect 4982 11608 4988 11620
rect 3988 11580 4988 11608
rect 4982 11568 4988 11580
rect 5040 11568 5046 11620
rect 9324 11608 9352 11639
rect 9582 11636 9588 11639
rect 9640 11636 9646 11688
rect 12342 11636 12348 11688
rect 12400 11676 12406 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 12400 11648 12449 11676
rect 12400 11636 12406 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 12693 11679 12751 11685
rect 12693 11676 12705 11679
rect 12584 11648 12705 11676
rect 12584 11636 12590 11648
rect 12693 11645 12705 11648
rect 12739 11645 12751 11679
rect 12693 11639 12751 11645
rect 9674 11608 9680 11620
rect 9324 11580 9680 11608
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 1670 11540 1676 11552
rect 1631 11512 1676 11540
rect 1670 11500 1676 11512
rect 1728 11500 1734 11552
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 3050 11540 3056 11552
rect 2188 11512 2233 11540
rect 3011 11512 3056 11540
rect 2188 11500 2194 11512
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 3697 11543 3755 11549
rect 3697 11540 3709 11543
rect 3660 11512 3709 11540
rect 3660 11500 3666 11512
rect 3697 11509 3709 11512
rect 3743 11509 3755 11543
rect 6546 11540 6552 11552
rect 6507 11512 6552 11540
rect 3697 11503 3755 11509
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 8849 11543 8907 11549
rect 8849 11509 8861 11543
rect 8895 11540 8907 11543
rect 9030 11540 9036 11552
rect 8895 11512 9036 11540
rect 8895 11509 8907 11512
rect 8849 11503 8907 11509
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 13814 11540 13820 11552
rect 13727 11512 13820 11540
rect 13814 11500 13820 11512
rect 13872 11540 13878 11552
rect 14737 11543 14795 11549
rect 14737 11540 14749 11543
rect 13872 11512 14749 11540
rect 13872 11500 13878 11512
rect 14737 11509 14749 11512
rect 14783 11509 14795 11543
rect 14737 11503 14795 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1765 11339 1823 11345
rect 1765 11305 1777 11339
rect 1811 11336 1823 11339
rect 2130 11336 2136 11348
rect 1811 11308 2136 11336
rect 1811 11305 1823 11308
rect 1765 11299 1823 11305
rect 2130 11296 2136 11308
rect 2188 11336 2194 11348
rect 3145 11339 3203 11345
rect 3145 11336 3157 11339
rect 2188 11308 3157 11336
rect 2188 11296 2194 11308
rect 3145 11305 3157 11308
rect 3191 11305 3203 11339
rect 4706 11336 4712 11348
rect 4667 11308 4712 11336
rect 3145 11299 3203 11305
rect 4706 11296 4712 11308
rect 4764 11296 4770 11348
rect 6270 11296 6276 11348
rect 6328 11336 6334 11348
rect 6365 11339 6423 11345
rect 6365 11336 6377 11339
rect 6328 11308 6377 11336
rect 6328 11296 6334 11308
rect 6365 11305 6377 11308
rect 6411 11336 6423 11339
rect 6914 11336 6920 11348
rect 6411 11308 6920 11336
rect 6411 11305 6423 11308
rect 6365 11299 6423 11305
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 7101 11339 7159 11345
rect 7101 11305 7113 11339
rect 7147 11336 7159 11339
rect 7466 11336 7472 11348
rect 7147 11308 7472 11336
rect 7147 11305 7159 11308
rect 7101 11299 7159 11305
rect 7466 11296 7472 11308
rect 7524 11296 7530 11348
rect 8478 11336 8484 11348
rect 8439 11308 8484 11336
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 8938 11336 8944 11348
rect 8899 11308 8944 11336
rect 8938 11296 8944 11308
rect 8996 11296 9002 11348
rect 10778 11296 10784 11348
rect 10836 11336 10842 11348
rect 11241 11339 11299 11345
rect 11241 11336 11253 11339
rect 10836 11308 11253 11336
rect 10836 11296 10842 11308
rect 11241 11305 11253 11308
rect 11287 11336 11299 11339
rect 11609 11339 11667 11345
rect 11609 11336 11621 11339
rect 11287 11308 11621 11336
rect 11287 11305 11299 11308
rect 11241 11299 11299 11305
rect 11609 11305 11621 11308
rect 11655 11336 11667 11339
rect 11977 11339 12035 11345
rect 11977 11336 11989 11339
rect 11655 11308 11989 11336
rect 11655 11305 11667 11308
rect 11609 11299 11667 11305
rect 11977 11305 11989 11308
rect 12023 11336 12035 11339
rect 12342 11336 12348 11348
rect 12023 11308 12348 11336
rect 12023 11305 12035 11308
rect 11977 11299 12035 11305
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 12526 11336 12532 11348
rect 12487 11308 12532 11336
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 14090 11336 14096 11348
rect 14051 11308 14096 11336
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 1670 11228 1676 11280
rect 1728 11268 1734 11280
rect 3513 11271 3571 11277
rect 3513 11268 3525 11271
rect 1728 11240 3525 11268
rect 1728 11228 1734 11240
rect 3513 11237 3525 11240
rect 3559 11237 3571 11271
rect 3513 11231 3571 11237
rect 5252 11271 5310 11277
rect 5252 11237 5264 11271
rect 5298 11268 5310 11271
rect 5442 11268 5448 11280
rect 5298 11240 5448 11268
rect 5298 11237 5310 11240
rect 5252 11231 5310 11237
rect 5442 11228 5448 11240
rect 5500 11228 5506 11280
rect 1854 11160 1860 11212
rect 1912 11200 1918 11212
rect 2133 11203 2191 11209
rect 2133 11200 2145 11203
rect 1912 11172 2145 11200
rect 1912 11160 1918 11172
rect 2133 11169 2145 11172
rect 2179 11200 2191 11203
rect 2498 11200 2504 11212
rect 2179 11172 2504 11200
rect 2179 11169 2191 11172
rect 2133 11163 2191 11169
rect 2498 11160 2504 11172
rect 2556 11200 2562 11212
rect 4341 11203 4399 11209
rect 4341 11200 4353 11203
rect 2556 11172 4353 11200
rect 2556 11160 2562 11172
rect 4341 11169 4353 11172
rect 4387 11200 4399 11203
rect 4522 11200 4528 11212
rect 4387 11172 4528 11200
rect 4387 11169 4399 11172
rect 4341 11163 4399 11169
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 4982 11200 4988 11212
rect 4943 11172 4988 11200
rect 4982 11160 4988 11172
rect 5040 11200 5046 11212
rect 5534 11200 5540 11212
rect 5040 11172 5540 11200
rect 5040 11160 5046 11172
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11200 7895 11203
rect 8478 11200 8484 11212
rect 7883 11172 8484 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 8754 11160 8760 11212
rect 8812 11200 8818 11212
rect 9217 11203 9275 11209
rect 9217 11200 9229 11203
rect 8812 11172 9229 11200
rect 8812 11160 8818 11172
rect 9217 11169 9229 11172
rect 9263 11169 9275 11203
rect 9217 11163 9275 11169
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11200 10655 11203
rect 10962 11200 10968 11212
rect 10643 11172 10968 11200
rect 10643 11169 10655 11172
rect 10597 11163 10655 11169
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 12360 11200 12388 11296
rect 12980 11271 13038 11277
rect 12980 11237 12992 11271
rect 13026 11268 13038 11271
rect 13722 11268 13728 11280
rect 13026 11240 13728 11268
rect 13026 11237 13038 11240
rect 12980 11231 13038 11237
rect 13722 11228 13728 11240
rect 13780 11228 13786 11280
rect 12713 11203 12771 11209
rect 12713 11200 12725 11203
rect 12360 11172 12725 11200
rect 12713 11169 12725 11172
rect 12759 11200 12771 11203
rect 12802 11200 12808 11212
rect 12759 11172 12808 11200
rect 12759 11169 12771 11172
rect 12713 11163 12771 11169
rect 12802 11160 12808 11172
rect 12860 11160 12866 11212
rect 18506 11200 18512 11212
rect 18467 11172 18512 11200
rect 18506 11160 18512 11172
rect 18564 11160 18570 11212
rect 18782 11200 18788 11212
rect 18743 11172 18788 11200
rect 18782 11160 18788 11172
rect 18840 11160 18846 11212
rect 1762 11092 1768 11144
rect 1820 11132 1826 11144
rect 2225 11135 2283 11141
rect 2225 11132 2237 11135
rect 1820 11104 2237 11132
rect 1820 11092 1826 11104
rect 2225 11101 2237 11104
rect 2271 11101 2283 11135
rect 2406 11132 2412 11144
rect 2367 11104 2412 11132
rect 2225 11095 2283 11101
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 7282 11092 7288 11144
rect 7340 11132 7346 11144
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 7340 11104 7941 11132
rect 7340 11092 7346 11104
rect 7929 11101 7941 11104
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11132 8171 11135
rect 8202 11132 8208 11144
rect 8159 11104 8208 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 10686 11132 10692 11144
rect 10647 11104 10692 11132
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 10778 11092 10784 11144
rect 10836 11132 10842 11144
rect 10836 11104 10881 11132
rect 10836 11092 10842 11104
rect 2130 11024 2136 11076
rect 2188 11064 2194 11076
rect 2777 11067 2835 11073
rect 2777 11064 2789 11067
rect 2188 11036 2789 11064
rect 2188 11024 2194 11036
rect 2777 11033 2789 11036
rect 2823 11064 2835 11067
rect 3050 11064 3056 11076
rect 2823 11036 3056 11064
rect 2823 11033 2835 11036
rect 2777 11027 2835 11033
rect 3050 11024 3056 11036
rect 3108 11024 3114 11076
rect 7466 11064 7472 11076
rect 7427 11036 7472 11064
rect 7466 11024 7472 11036
rect 7524 11024 7530 11076
rect 8294 11024 8300 11076
rect 8352 11064 8358 11076
rect 8570 11064 8576 11076
rect 8352 11036 8576 11064
rect 8352 11024 8358 11036
rect 8570 11024 8576 11036
rect 8628 11064 8634 11076
rect 9033 11067 9091 11073
rect 9033 11064 9045 11067
rect 8628 11036 9045 11064
rect 8628 11024 8634 11036
rect 9033 11033 9045 11036
rect 9079 11033 9091 11067
rect 10226 11064 10232 11076
rect 10187 11036 10232 11064
rect 9033 11027 9091 11033
rect 10226 11024 10232 11036
rect 10284 11024 10290 11076
rect 1673 10999 1731 11005
rect 1673 10965 1685 10999
rect 1719 10996 1731 10999
rect 2222 10996 2228 11008
rect 1719 10968 2228 10996
rect 1719 10965 1731 10968
rect 1673 10959 1731 10965
rect 2222 10956 2228 10968
rect 2280 10996 2286 11008
rect 2406 10996 2412 11008
rect 2280 10968 2412 10996
rect 2280 10956 2286 10968
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 10137 10999 10195 11005
rect 10137 10965 10149 10999
rect 10183 10996 10195 10999
rect 10870 10996 10876 11008
rect 10183 10968 10876 10996
rect 10183 10965 10195 10968
rect 10137 10959 10195 10965
rect 10870 10956 10876 10968
rect 10928 10956 10934 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 3234 10792 3240 10804
rect 3195 10764 3240 10792
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 4154 10792 4160 10804
rect 4115 10764 4160 10792
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 5442 10792 5448 10804
rect 5403 10764 5448 10792
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5721 10795 5779 10801
rect 5721 10792 5733 10795
rect 5592 10764 5733 10792
rect 5592 10752 5598 10764
rect 5721 10761 5733 10764
rect 5767 10792 5779 10795
rect 6089 10795 6147 10801
rect 6089 10792 6101 10795
rect 5767 10764 6101 10792
rect 5767 10761 5779 10764
rect 5721 10755 5779 10761
rect 6089 10761 6101 10764
rect 6135 10761 6147 10795
rect 9030 10792 9036 10804
rect 8991 10764 9036 10792
rect 6089 10755 6147 10761
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 9677 10795 9735 10801
rect 9677 10761 9689 10795
rect 9723 10792 9735 10795
rect 9766 10792 9772 10804
rect 9723 10764 9772 10792
rect 9723 10761 9735 10764
rect 9677 10755 9735 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10137 10795 10195 10801
rect 10137 10792 10149 10795
rect 10100 10764 10149 10792
rect 10100 10752 10106 10764
rect 10137 10761 10149 10764
rect 10183 10792 10195 10795
rect 10686 10792 10692 10804
rect 10183 10764 10692 10792
rect 10183 10761 10195 10764
rect 10137 10755 10195 10761
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 12434 10792 12440 10804
rect 12395 10764 12440 10792
rect 12434 10752 12440 10764
rect 12492 10752 12498 10804
rect 13541 10795 13599 10801
rect 13541 10761 13553 10795
rect 13587 10792 13599 10795
rect 13722 10792 13728 10804
rect 13587 10764 13728 10792
rect 13587 10761 13599 10764
rect 13541 10755 13599 10761
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 18506 10792 18512 10804
rect 18467 10764 18512 10792
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10656 3939 10659
rect 4985 10659 5043 10665
rect 4985 10656 4997 10659
rect 3927 10628 4997 10656
rect 3927 10625 3939 10628
rect 3881 10619 3939 10625
rect 4985 10625 4997 10628
rect 5031 10656 5043 10659
rect 5460 10656 5488 10752
rect 5031 10628 5488 10656
rect 5031 10625 5043 10628
rect 4985 10619 5043 10625
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 7653 10659 7711 10665
rect 7653 10656 7665 10659
rect 7616 10628 7665 10656
rect 7616 10616 7622 10628
rect 7653 10625 7665 10628
rect 7699 10625 7711 10659
rect 9784 10656 9812 10752
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 9784 10628 10609 10656
rect 7653 10619 7711 10625
rect 10597 10625 10609 10628
rect 10643 10625 10655 10659
rect 10597 10619 10655 10625
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10656 10839 10659
rect 10870 10656 10876 10668
rect 10827 10628 10876 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 12526 10616 12532 10668
rect 12584 10656 12590 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12584 10628 13001 10656
rect 12584 10616 12590 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 20441 10659 20499 10665
rect 20441 10625 20453 10659
rect 20487 10656 20499 10659
rect 21358 10656 21364 10668
rect 20487 10628 21364 10656
rect 20487 10625 20499 10628
rect 20441 10619 20499 10625
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 2406 10588 2412 10600
rect 1903 10560 2412 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 4154 10548 4160 10600
rect 4212 10588 4218 10600
rect 4709 10591 4767 10597
rect 4709 10588 4721 10591
rect 4212 10560 4721 10588
rect 4212 10548 4218 10560
rect 4709 10557 4721 10560
rect 4755 10557 4767 10591
rect 20162 10588 20168 10600
rect 20123 10560 20168 10588
rect 4709 10551 4767 10557
rect 20162 10548 20168 10560
rect 20220 10588 20226 10600
rect 20901 10591 20959 10597
rect 20901 10588 20913 10591
rect 20220 10560 20913 10588
rect 20220 10548 20226 10560
rect 20901 10557 20913 10560
rect 20947 10557 20959 10591
rect 20901 10551 20959 10557
rect 2130 10529 2136 10532
rect 2124 10520 2136 10529
rect 2091 10492 2136 10520
rect 2124 10483 2136 10492
rect 2130 10480 2136 10483
rect 2188 10480 2194 10532
rect 4522 10480 4528 10532
rect 4580 10520 4586 10532
rect 4801 10523 4859 10529
rect 4801 10520 4813 10523
rect 4580 10492 4813 10520
rect 4580 10480 4586 10492
rect 4801 10489 4813 10492
rect 4847 10489 4859 10523
rect 4801 10483 4859 10489
rect 6641 10523 6699 10529
rect 6641 10489 6653 10523
rect 6687 10520 6699 10523
rect 7282 10520 7288 10532
rect 6687 10492 7288 10520
rect 6687 10489 6699 10492
rect 6641 10483 6699 10489
rect 7282 10480 7288 10492
rect 7340 10480 7346 10532
rect 7561 10523 7619 10529
rect 7561 10489 7573 10523
rect 7607 10520 7619 10523
rect 7920 10523 7978 10529
rect 7920 10520 7932 10523
rect 7607 10492 7932 10520
rect 7607 10489 7619 10492
rect 7561 10483 7619 10489
rect 7920 10489 7932 10492
rect 7966 10520 7978 10523
rect 8202 10520 8208 10532
rect 7966 10492 8208 10520
rect 7966 10489 7978 10492
rect 7920 10483 7978 10489
rect 1762 10452 1768 10464
rect 1723 10424 1768 10452
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 4341 10455 4399 10461
rect 4341 10421 4353 10455
rect 4387 10452 4399 10455
rect 4614 10452 4620 10464
rect 4387 10424 4620 10452
rect 4387 10421 4399 10424
rect 4341 10415 4399 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 7193 10455 7251 10461
rect 7193 10421 7205 10455
rect 7239 10452 7251 10455
rect 7576 10452 7604 10483
rect 8202 10480 8208 10492
rect 8260 10480 8266 10532
rect 10505 10523 10563 10529
rect 10505 10520 10517 10523
rect 9968 10492 10517 10520
rect 9968 10464 9996 10492
rect 10505 10489 10517 10492
rect 10551 10489 10563 10523
rect 12158 10520 12164 10532
rect 12119 10492 12164 10520
rect 10505 10483 10563 10489
rect 12158 10480 12164 10492
rect 12216 10520 12222 10532
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 12216 10492 12817 10520
rect 12216 10480 12222 10492
rect 12805 10489 12817 10492
rect 12851 10489 12863 10523
rect 12805 10483 12863 10489
rect 9950 10452 9956 10464
rect 7239 10424 7604 10452
rect 9911 10424 9956 10452
rect 7239 10421 7251 10424
rect 7193 10415 7251 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11149 10455 11207 10461
rect 11149 10452 11161 10455
rect 11112 10424 11161 10452
rect 11112 10412 11118 10424
rect 11149 10421 11161 10424
rect 11195 10421 11207 10455
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 11149 10415 11207 10421
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 12897 10455 12955 10461
rect 12897 10452 12909 10455
rect 12768 10424 12909 10452
rect 12768 10412 12774 10424
rect 12897 10421 12909 10424
rect 12943 10421 12955 10455
rect 12897 10415 12955 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 2225 10251 2283 10257
rect 2225 10217 2237 10251
rect 2271 10248 2283 10251
rect 2314 10248 2320 10260
rect 2271 10220 2320 10248
rect 2271 10217 2283 10220
rect 2225 10211 2283 10217
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 2593 10251 2651 10257
rect 2593 10217 2605 10251
rect 2639 10248 2651 10251
rect 2682 10248 2688 10260
rect 2639 10220 2688 10248
rect 2639 10217 2651 10220
rect 2593 10211 2651 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 4614 10208 4620 10260
rect 4672 10248 4678 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 4672 10220 5457 10248
rect 4672 10208 4678 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 5626 10248 5632 10260
rect 5587 10220 5632 10248
rect 5445 10211 5503 10217
rect 5460 10180 5488 10211
rect 5626 10208 5632 10220
rect 5684 10208 5690 10260
rect 5994 10248 6000 10260
rect 5907 10220 6000 10248
rect 5994 10208 6000 10220
rect 6052 10248 6058 10260
rect 6822 10248 6828 10260
rect 6052 10220 6828 10248
rect 6052 10208 6058 10220
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7282 10248 7288 10260
rect 7243 10220 7288 10248
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 7742 10248 7748 10260
rect 7703 10220 7748 10248
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 8754 10208 8760 10260
rect 8812 10248 8818 10260
rect 9033 10251 9091 10257
rect 9033 10248 9045 10251
rect 8812 10220 9045 10248
rect 8812 10208 8818 10220
rect 9033 10217 9045 10220
rect 9079 10217 9091 10251
rect 10042 10248 10048 10260
rect 10003 10220 10048 10248
rect 9033 10211 9091 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 12710 10248 12716 10260
rect 12575 10220 12716 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 13173 10251 13231 10257
rect 13173 10248 13185 10251
rect 12860 10220 13185 10248
rect 12860 10208 12866 10220
rect 13173 10217 13185 10220
rect 13219 10217 13231 10251
rect 13173 10211 13231 10217
rect 6089 10183 6147 10189
rect 6089 10180 6101 10183
rect 5460 10152 6101 10180
rect 6089 10149 6101 10152
rect 6135 10149 6147 10183
rect 6089 10143 6147 10149
rect 10226 10140 10232 10192
rect 10284 10180 10290 10192
rect 10404 10183 10462 10189
rect 10404 10180 10416 10183
rect 10284 10152 10416 10180
rect 10284 10140 10290 10152
rect 10404 10149 10416 10152
rect 10450 10180 10462 10183
rect 10870 10180 10876 10192
rect 10450 10152 10876 10180
rect 10450 10149 10462 10152
rect 10404 10143 10462 10149
rect 10870 10140 10876 10152
rect 10928 10140 10934 10192
rect 1578 10072 1584 10124
rect 1636 10112 1642 10124
rect 2498 10112 2504 10124
rect 1636 10084 2504 10112
rect 1636 10072 1642 10084
rect 2498 10072 2504 10084
rect 2556 10112 2562 10124
rect 2682 10112 2688 10124
rect 2556 10084 2688 10112
rect 2556 10072 2562 10084
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 4430 10112 4436 10124
rect 4391 10084 4436 10112
rect 4430 10072 4436 10084
rect 4488 10072 4494 10124
rect 7650 10112 7656 10124
rect 7611 10084 7656 10112
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 18874 10112 18880 10124
rect 18835 10084 18880 10112
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 19150 10112 19156 10124
rect 19111 10084 19156 10112
rect 19150 10072 19156 10084
rect 19208 10072 19214 10124
rect 2222 10004 2228 10056
rect 2280 10044 2286 10056
rect 2777 10047 2835 10053
rect 2777 10044 2789 10047
rect 2280 10016 2789 10044
rect 2280 10004 2286 10016
rect 2777 10013 2789 10016
rect 2823 10044 2835 10047
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 2823 10016 3249 10044
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 3237 10013 3249 10016
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4212 10016 4537 10044
rect 4212 10004 4218 10016
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4706 10044 4712 10056
rect 4667 10016 4712 10044
rect 4525 10007 4583 10013
rect 4062 9976 4068 9988
rect 4023 9948 4068 9976
rect 4062 9936 4068 9948
rect 4120 9936 4126 9988
rect 4540 9976 4568 10007
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 6270 10044 6276 10056
rect 6231 10016 6276 10044
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 7837 10047 7895 10053
rect 7837 10044 7849 10047
rect 7239 10016 7849 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 7837 10013 7849 10016
rect 7883 10044 7895 10047
rect 7926 10044 7932 10056
rect 7883 10016 7932 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 7926 10004 7932 10016
rect 7984 10044 7990 10056
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 7984 10016 8309 10044
rect 7984 10004 7990 10016
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 10134 10044 10140 10056
rect 8297 10007 8355 10013
rect 9416 10016 10140 10044
rect 5077 9979 5135 9985
rect 5077 9976 5089 9979
rect 4540 9948 5089 9976
rect 5077 9945 5089 9948
rect 5123 9945 5135 9979
rect 5077 9939 5135 9945
rect 3878 9908 3884 9920
rect 3839 9880 3884 9908
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 6822 9908 6828 9920
rect 6783 9880 6828 9908
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 9416 9917 9444 10016
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 8665 9911 8723 9917
rect 8665 9908 8677 9911
rect 7616 9880 8677 9908
rect 7616 9868 7622 9880
rect 8665 9877 8677 9880
rect 8711 9908 8723 9911
rect 9401 9911 9459 9917
rect 9401 9908 9413 9911
rect 8711 9880 9413 9908
rect 8711 9877 8723 9880
rect 8665 9871 8723 9877
rect 9401 9877 9413 9880
rect 9447 9877 9459 9911
rect 9401 9871 9459 9877
rect 10778 9868 10784 9920
rect 10836 9908 10842 9920
rect 11514 9908 11520 9920
rect 10836 9880 11520 9908
rect 10836 9868 10842 9880
rect 11514 9868 11520 9880
rect 11572 9868 11578 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 4430 9704 4436 9716
rect 4080 9676 4436 9704
rect 3973 9639 4031 9645
rect 3973 9605 3985 9639
rect 4019 9636 4031 9639
rect 4080 9636 4108 9676
rect 4430 9664 4436 9676
rect 4488 9664 4494 9716
rect 5994 9704 6000 9716
rect 5955 9676 6000 9704
rect 5994 9664 6000 9676
rect 6052 9664 6058 9716
rect 7650 9704 7656 9716
rect 6932 9676 7656 9704
rect 6638 9636 6644 9648
rect 4019 9608 4108 9636
rect 6551 9608 6644 9636
rect 4019 9605 4031 9608
rect 3973 9599 4031 9605
rect 6638 9596 6644 9608
rect 6696 9636 6702 9648
rect 6932 9636 6960 9676
rect 7650 9664 7656 9676
rect 7708 9664 7714 9716
rect 10226 9704 10232 9716
rect 10187 9676 10232 9704
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 18874 9704 18880 9716
rect 18835 9676 18880 9704
rect 18874 9664 18880 9676
rect 18932 9664 18938 9716
rect 9674 9636 9680 9648
rect 6696 9608 6960 9636
rect 9635 9608 9680 9636
rect 6696 9596 6702 9608
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 10962 9568 10968 9580
rect 10459 9540 10968 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 19613 9571 19671 9577
rect 19613 9537 19625 9571
rect 19659 9568 19671 9571
rect 20622 9568 20628 9580
rect 19659 9540 20628 9568
rect 19659 9537 19671 9540
rect 19613 9531 19671 9537
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 1581 9503 1639 9509
rect 1581 9469 1593 9503
rect 1627 9500 1639 9503
rect 2590 9500 2596 9512
rect 1627 9472 2596 9500
rect 1627 9469 1639 9472
rect 1581 9463 1639 9469
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9500 4123 9503
rect 4154 9500 4160 9512
rect 4111 9472 4160 9500
rect 4111 9469 4123 9472
rect 4065 9463 4123 9469
rect 4154 9460 4160 9472
rect 4212 9500 4218 9512
rect 5442 9500 5448 9512
rect 4212 9472 5448 9500
rect 4212 9460 4218 9472
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 7558 9500 7564 9512
rect 6972 9472 7564 9500
rect 6972 9460 6978 9472
rect 7558 9460 7564 9472
rect 7616 9500 7622 9512
rect 7926 9509 7932 9512
rect 7653 9503 7711 9509
rect 7653 9500 7665 9503
rect 7616 9472 7665 9500
rect 7616 9460 7622 9472
rect 7653 9469 7665 9472
rect 7699 9469 7711 9503
rect 7920 9500 7932 9509
rect 7887 9472 7932 9500
rect 7653 9463 7711 9469
rect 7920 9463 7932 9472
rect 7926 9460 7932 9463
rect 7984 9460 7990 9512
rect 19334 9460 19340 9512
rect 19392 9500 19398 9512
rect 20073 9503 20131 9509
rect 20073 9500 20085 9503
rect 19392 9472 20085 9500
rect 19392 9460 19398 9472
rect 20073 9469 20085 9472
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 1848 9435 1906 9441
rect 1848 9401 1860 9435
rect 1894 9432 1906 9435
rect 2222 9432 2228 9444
rect 1894 9404 2228 9432
rect 1894 9401 1906 9404
rect 1848 9395 1906 9401
rect 2222 9392 2228 9404
rect 2280 9432 2286 9444
rect 3513 9435 3571 9441
rect 3513 9432 3525 9435
rect 2280 9404 3525 9432
rect 2280 9392 2286 9404
rect 3513 9401 3525 9404
rect 3559 9401 3571 9435
rect 3513 9395 3571 9401
rect 3878 9392 3884 9444
rect 3936 9432 3942 9444
rect 4332 9435 4390 9441
rect 4332 9432 4344 9435
rect 3936 9404 4344 9432
rect 3936 9392 3942 9404
rect 4332 9401 4344 9404
rect 4378 9432 4390 9435
rect 5074 9432 5080 9444
rect 4378 9404 5080 9432
rect 4378 9401 4390 9404
rect 4332 9395 4390 9401
rect 5074 9392 5080 9404
rect 5132 9392 5138 9444
rect 7377 9435 7435 9441
rect 7377 9401 7389 9435
rect 7423 9432 7435 9435
rect 7742 9432 7748 9444
rect 7423 9404 7748 9432
rect 7423 9401 7435 9404
rect 7377 9395 7435 9401
rect 7742 9392 7748 9404
rect 7800 9392 7806 9444
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 2961 9367 3019 9373
rect 2961 9364 2973 9367
rect 2188 9336 2973 9364
rect 2188 9324 2194 9336
rect 2961 9333 2973 9336
rect 3007 9333 3019 9367
rect 5442 9364 5448 9376
rect 5403 9336 5448 9364
rect 2961 9327 3019 9333
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 9033 9367 9091 9373
rect 9033 9364 9045 9367
rect 8352 9336 9045 9364
rect 8352 9324 8358 9336
rect 9033 9333 9045 9336
rect 9079 9333 9091 9367
rect 9033 9327 9091 9333
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10873 9367 10931 9373
rect 10873 9364 10885 9367
rect 10192 9336 10885 9364
rect 10192 9324 10198 9336
rect 10873 9333 10885 9336
rect 10919 9333 10931 9367
rect 10873 9327 10931 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2682 9160 2688 9172
rect 2643 9132 2688 9160
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2924 9132 2973 9160
rect 2924 9120 2930 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 2961 9123 3019 9129
rect 3421 9163 3479 9169
rect 3421 9129 3433 9163
rect 3467 9160 3479 9163
rect 4154 9160 4160 9172
rect 3467 9132 4160 9160
rect 3467 9129 3479 9132
rect 3421 9123 3479 9129
rect 1949 9095 2007 9101
rect 1949 9061 1961 9095
rect 1995 9092 2007 9095
rect 2038 9092 2044 9104
rect 1995 9064 2044 9092
rect 1995 9061 2007 9064
rect 1949 9055 2007 9061
rect 2038 9052 2044 9064
rect 2096 9052 2102 9104
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 3436 9092 3464 9123
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 6270 9120 6276 9172
rect 6328 9160 6334 9172
rect 6365 9163 6423 9169
rect 6365 9160 6377 9163
rect 6328 9132 6377 9160
rect 6328 9120 6334 9132
rect 6365 9129 6377 9132
rect 6411 9129 6423 9163
rect 6365 9123 6423 9129
rect 7926 9120 7932 9172
rect 7984 9160 7990 9172
rect 8297 9163 8355 9169
rect 8297 9160 8309 9163
rect 7984 9132 8309 9160
rect 7984 9120 7990 9132
rect 8297 9129 8309 9132
rect 8343 9160 8355 9163
rect 8938 9160 8944 9172
rect 8343 9132 8944 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 11882 9160 11888 9172
rect 11843 9132 11888 9160
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 4706 9101 4712 9104
rect 2556 9064 3464 9092
rect 4341 9095 4399 9101
rect 2556 9052 2562 9064
rect 4341 9061 4353 9095
rect 4387 9092 4399 9095
rect 4700 9092 4712 9101
rect 4387 9064 4712 9092
rect 4387 9061 4399 9064
rect 4341 9055 4399 9061
rect 4700 9055 4712 9064
rect 4764 9092 4770 9104
rect 5442 9092 5448 9104
rect 4764 9064 5448 9092
rect 4706 9052 4712 9055
rect 4764 9052 4770 9064
rect 5442 9052 5448 9064
rect 5500 9052 5506 9104
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 3605 9027 3663 9033
rect 3605 9024 3617 9027
rect 3568 8996 3617 9024
rect 3568 8984 3574 8996
rect 3605 8993 3617 8996
rect 3651 8993 3663 9027
rect 3605 8987 3663 8993
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 4433 9027 4491 9033
rect 4433 9024 4445 9027
rect 4212 8996 4445 9024
rect 4212 8984 4218 8996
rect 4433 8993 4445 8996
rect 4479 9024 4491 9027
rect 4522 9024 4528 9036
rect 4479 8996 4528 9024
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 7184 9027 7242 9033
rect 7184 8993 7196 9027
rect 7230 9024 7242 9027
rect 7466 9024 7472 9036
rect 7230 8996 7472 9024
rect 7230 8993 7242 8996
rect 7184 8987 7242 8993
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 10134 8984 10140 9036
rect 10192 9024 10198 9036
rect 10505 9027 10563 9033
rect 10505 9024 10517 9027
rect 10192 8996 10517 9024
rect 10192 8984 10198 8996
rect 10505 8993 10517 8996
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 10594 8984 10600 9036
rect 10652 9024 10658 9036
rect 10778 9033 10784 9036
rect 10761 9027 10784 9033
rect 10761 9024 10773 9027
rect 10652 8996 10773 9024
rect 10652 8984 10658 8996
rect 10761 8993 10773 8996
rect 10836 9024 10842 9036
rect 10836 8996 10909 9024
rect 10761 8987 10784 8993
rect 10778 8984 10784 8987
rect 10836 8984 10842 8996
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8925 2099 8959
rect 2222 8956 2228 8968
rect 2183 8928 2228 8956
rect 2041 8919 2099 8925
rect 2056 8888 2084 8919
rect 2222 8916 2228 8928
rect 2280 8916 2286 8968
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 6972 8928 7017 8956
rect 6972 8916 6978 8928
rect 2682 8888 2688 8900
rect 2056 8860 2688 8888
rect 2682 8848 2688 8860
rect 2740 8848 2746 8900
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 5592 8792 5825 8820
rect 5592 8780 5598 8792
rect 5813 8789 5825 8792
rect 5859 8789 5871 8823
rect 6730 8820 6736 8832
rect 6691 8792 6736 8820
rect 5813 8783 5871 8789
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 1946 8616 1952 8628
rect 1627 8588 1952 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 2682 8616 2688 8628
rect 2643 8588 2688 8616
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 2958 8616 2964 8628
rect 2919 8588 2964 8616
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 3145 8619 3203 8625
rect 3145 8585 3157 8619
rect 3191 8616 3203 8619
rect 4062 8616 4068 8628
rect 3191 8588 4068 8616
rect 3191 8585 3203 8588
rect 3145 8579 3203 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 4706 8616 4712 8628
rect 4571 8588 4712 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 4890 8616 4896 8628
rect 4851 8588 4896 8616
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 6730 8616 6736 8628
rect 5123 8588 6736 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 6730 8576 6736 8588
rect 6788 8616 6794 8628
rect 8294 8616 8300 8628
rect 6788 8588 7328 8616
rect 8255 8588 8300 8616
rect 6788 8576 6794 8588
rect 6822 8548 6828 8560
rect 6783 8520 6828 8548
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 1636 8452 2053 8480
rect 1636 8440 1642 8452
rect 2041 8449 2053 8452
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2056 8412 2084 8443
rect 2130 8440 2136 8492
rect 2188 8480 2194 8492
rect 2188 8452 2233 8480
rect 2188 8440 2194 8452
rect 2866 8440 2872 8492
rect 2924 8480 2930 8492
rect 3605 8483 3663 8489
rect 3605 8480 3617 8483
rect 2924 8452 3617 8480
rect 2924 8440 2930 8452
rect 3605 8449 3617 8452
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 3789 8483 3847 8489
rect 3789 8449 3801 8483
rect 3835 8480 3847 8483
rect 3878 8480 3884 8492
rect 3835 8452 3884 8480
rect 3835 8449 3847 8452
rect 3789 8443 3847 8449
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 7300 8489 7328 8588
rect 8294 8576 8300 8588
rect 8352 8616 8358 8628
rect 10594 8616 10600 8628
rect 8352 8588 8892 8616
rect 10555 8588 10600 8616
rect 8352 8576 8358 8588
rect 8389 8551 8447 8557
rect 8389 8517 8401 8551
rect 8435 8548 8447 8551
rect 8478 8548 8484 8560
rect 8435 8520 8484 8548
rect 8435 8517 8447 8520
rect 8389 8511 8447 8517
rect 8478 8508 8484 8520
rect 8536 8508 8542 8560
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 5592 8452 5641 8480
rect 5592 8440 5598 8452
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7466 8480 7472 8492
rect 7427 8452 7472 8480
rect 7285 8443 7343 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 8864 8489 8892 8588
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 10134 8508 10140 8560
rect 10192 8548 10198 8560
rect 10873 8551 10931 8557
rect 10873 8548 10885 8551
rect 10192 8520 10885 8548
rect 10192 8508 10198 8520
rect 10873 8517 10885 8520
rect 10919 8517 10931 8551
rect 10873 8511 10931 8517
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 8996 8452 9041 8480
rect 8996 8440 9002 8452
rect 2774 8412 2780 8424
rect 2056 8384 2780 8412
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 2958 8372 2964 8424
rect 3016 8412 3022 8424
rect 3513 8415 3571 8421
rect 3513 8412 3525 8415
rect 3016 8384 3525 8412
rect 3016 8372 3022 8384
rect 3513 8381 3525 8384
rect 3559 8381 3571 8415
rect 3513 8375 3571 8381
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 5445 8415 5503 8421
rect 5445 8412 5457 8415
rect 4948 8384 5457 8412
rect 4948 8372 4954 8384
rect 5445 8381 5457 8384
rect 5491 8381 5503 8415
rect 5445 8375 5503 8381
rect 6273 8415 6331 8421
rect 6273 8381 6285 8415
rect 6319 8412 6331 8415
rect 7484 8412 7512 8440
rect 6319 8384 7512 8412
rect 6319 8381 6331 8384
rect 6273 8375 6331 8381
rect 4798 8304 4804 8356
rect 4856 8344 4862 8356
rect 5537 8347 5595 8353
rect 5537 8344 5549 8347
rect 4856 8316 5549 8344
rect 4856 8304 4862 8316
rect 5537 8313 5549 8316
rect 5583 8313 5595 8347
rect 5537 8307 5595 8313
rect 6641 8347 6699 8353
rect 6641 8313 6653 8347
rect 6687 8344 6699 8347
rect 6730 8344 6736 8356
rect 6687 8316 6736 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 6730 8304 6736 8316
rect 6788 8344 6794 8356
rect 7193 8347 7251 8353
rect 7193 8344 7205 8347
rect 6788 8316 7205 8344
rect 6788 8304 6794 8316
rect 7193 8313 7205 8316
rect 7239 8313 7251 8347
rect 8757 8347 8815 8353
rect 8757 8344 8769 8347
rect 7193 8307 7251 8313
rect 8128 8316 8769 8344
rect 8128 8288 8156 8316
rect 8757 8313 8769 8316
rect 8803 8313 8815 8347
rect 8757 8307 8815 8313
rect 1946 8276 1952 8288
rect 1907 8248 1952 8276
rect 1946 8236 1952 8248
rect 2004 8236 2010 8288
rect 7929 8279 7987 8285
rect 7929 8245 7941 8279
rect 7975 8276 7987 8279
rect 8110 8276 8116 8288
rect 7975 8248 8116 8276
rect 7975 8245 7987 8248
rect 7929 8239 7987 8245
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 1946 8072 1952 8084
rect 1627 8044 1952 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 1946 8032 1952 8044
rect 2004 8072 2010 8084
rect 2409 8075 2467 8081
rect 2409 8072 2421 8075
rect 2004 8044 2421 8072
rect 2004 8032 2010 8044
rect 2409 8041 2421 8044
rect 2455 8041 2467 8075
rect 2774 8072 2780 8084
rect 2735 8044 2780 8072
rect 2409 8035 2467 8041
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 3145 8075 3203 8081
rect 3145 8072 3157 8075
rect 2924 8044 3157 8072
rect 2924 8032 2930 8044
rect 3145 8041 3157 8044
rect 3191 8041 3203 8075
rect 3145 8035 3203 8041
rect 3605 8075 3663 8081
rect 3605 8041 3617 8075
rect 3651 8072 3663 8075
rect 3878 8072 3884 8084
rect 3651 8044 3884 8072
rect 3651 8041 3663 8044
rect 3605 8035 3663 8041
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 4157 8075 4215 8081
rect 4157 8041 4169 8075
rect 4203 8072 4215 8075
rect 4430 8072 4436 8084
rect 4203 8044 4436 8072
rect 4203 8041 4215 8044
rect 4157 8035 4215 8041
rect 4430 8032 4436 8044
rect 4488 8032 4494 8084
rect 4522 8032 4528 8084
rect 4580 8072 4586 8084
rect 4617 8075 4675 8081
rect 4617 8072 4629 8075
rect 4580 8044 4629 8072
rect 4580 8032 4586 8044
rect 4617 8041 4629 8044
rect 4663 8041 4675 8075
rect 4617 8035 4675 8041
rect 4798 8032 4804 8084
rect 4856 8072 4862 8084
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 4856 8044 5089 8072
rect 4856 8032 4862 8044
rect 5077 8041 5089 8044
rect 5123 8041 5135 8075
rect 5534 8072 5540 8084
rect 5495 8044 5540 8072
rect 5077 8035 5135 8041
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 7009 8075 7067 8081
rect 7009 8041 7021 8075
rect 7055 8072 7067 8075
rect 7466 8072 7472 8084
rect 7055 8044 7472 8072
rect 7055 8041 7067 8044
rect 7009 8035 7067 8041
rect 7466 8032 7472 8044
rect 7524 8072 7530 8084
rect 7561 8075 7619 8081
rect 7561 8072 7573 8075
rect 7524 8044 7573 8072
rect 7524 8032 7530 8044
rect 7561 8041 7573 8044
rect 7607 8041 7619 8075
rect 8110 8072 8116 8084
rect 8071 8044 8116 8072
rect 7561 8035 7619 8041
rect 8110 8032 8116 8044
rect 8168 8032 8174 8084
rect 8665 8075 8723 8081
rect 8665 8041 8677 8075
rect 8711 8072 8723 8075
rect 8938 8072 8944 8084
rect 8711 8044 8944 8072
rect 8711 8041 8723 8044
rect 8665 8035 8723 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 2038 8004 2044 8016
rect 1999 7976 2044 8004
rect 2038 7964 2044 7976
rect 2096 7964 2102 8016
rect 5552 8004 5580 8032
rect 5874 8007 5932 8013
rect 5874 8004 5886 8007
rect 5552 7976 5886 8004
rect 5874 7973 5886 7976
rect 5920 8004 5932 8007
rect 5994 8004 6000 8016
rect 5920 7976 6000 8004
rect 5920 7973 5932 7976
rect 5874 7967 5932 7973
rect 5994 7964 6000 7976
rect 6052 7964 6058 8016
rect 5534 7828 5540 7880
rect 5592 7868 5598 7880
rect 5629 7871 5687 7877
rect 5629 7868 5641 7871
rect 5592 7840 5641 7868
rect 5592 7828 5598 7840
rect 5629 7837 5641 7840
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2041 7531 2099 7537
rect 2041 7497 2053 7531
rect 2087 7528 2099 7531
rect 2130 7528 2136 7540
rect 2087 7500 2136 7528
rect 2087 7497 2099 7500
rect 2041 7491 2099 7497
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 2314 7488 2320 7540
rect 2372 7528 2378 7540
rect 2409 7531 2467 7537
rect 2409 7528 2421 7531
rect 2372 7500 2421 7528
rect 2372 7488 2378 7500
rect 2409 7497 2421 7500
rect 2455 7528 2467 7531
rect 2498 7528 2504 7540
rect 2455 7500 2504 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 3510 7528 3516 7540
rect 3471 7500 3516 7528
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 4522 7528 4528 7540
rect 4483 7500 4528 7528
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 5997 7531 6055 7537
rect 5997 7528 6009 7531
rect 5592 7500 6009 7528
rect 5592 7488 5598 7500
rect 5997 7497 6009 7500
rect 6043 7528 6055 7531
rect 6914 7528 6920 7540
rect 6043 7500 6920 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6914 7488 6920 7500
rect 6972 7528 6978 7540
rect 7285 7531 7343 7537
rect 7285 7528 7297 7531
rect 6972 7500 7297 7528
rect 6972 7488 6978 7500
rect 7285 7497 7297 7500
rect 7331 7528 7343 7531
rect 8113 7531 8171 7537
rect 8113 7528 8125 7531
rect 7331 7500 8125 7528
rect 7331 7497 7343 7500
rect 7285 7491 7343 7497
rect 8113 7497 8125 7500
rect 8159 7497 8171 7531
rect 8570 7528 8576 7540
rect 8531 7500 8576 7528
rect 8113 7491 8171 7497
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 22465 7531 22523 7537
rect 22465 7497 22477 7531
rect 22511 7528 22523 7531
rect 23566 7528 23572 7540
rect 22511 7500 23572 7528
rect 22511 7497 22523 7500
rect 22465 7491 22523 7497
rect 23566 7488 23572 7500
rect 23624 7488 23630 7540
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7392 5779 7395
rect 5994 7392 6000 7404
rect 5767 7364 6000 7392
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 6825 7395 6883 7401
rect 6825 7392 6837 7395
rect 6788 7364 6837 7392
rect 6788 7352 6794 7364
rect 6825 7361 6837 7364
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 8297 7327 8355 7333
rect 8297 7293 8309 7327
rect 8343 7324 8355 7327
rect 8570 7324 8576 7336
rect 8343 7296 8576 7324
rect 8343 7293 8355 7296
rect 8297 7287 8355 7293
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 22278 7324 22284 7336
rect 22239 7296 22284 7324
rect 22278 7284 22284 7296
rect 22336 7324 22342 7336
rect 22833 7327 22891 7333
rect 22833 7324 22845 7327
rect 22336 7296 22845 7324
rect 22336 7284 22342 7296
rect 22833 7293 22845 7296
rect 22879 7293 22891 7327
rect 22833 7287 22891 7293
rect 1673 7191 1731 7197
rect 1673 7157 1685 7191
rect 1719 7188 1731 7191
rect 2222 7188 2228 7200
rect 1719 7160 2228 7188
rect 1719 7157 1731 7160
rect 1673 7151 1731 7157
rect 2222 7148 2228 7160
rect 2280 7188 2286 7200
rect 2682 7188 2688 7200
rect 2280 7160 2688 7188
rect 2280 7148 2286 7160
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 22738 6848 22744 6860
rect 22699 6820 22744 6848
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 22925 6715 22983 6721
rect 22925 6681 22937 6715
rect 22971 6712 22983 6715
rect 23382 6712 23388 6724
rect 22971 6684 23388 6712
rect 22971 6681 22983 6684
rect 22925 6675 22983 6681
rect 23382 6672 23388 6684
rect 23440 6672 23446 6724
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 22738 6440 22744 6452
rect 22699 6412 22744 6440
rect 22738 6400 22744 6412
rect 22796 6400 22802 6452
rect 23842 6440 23848 6452
rect 23803 6412 23848 6440
rect 23842 6400 23848 6412
rect 23900 6400 23906 6452
rect 23658 6236 23664 6248
rect 23619 6208 23664 6236
rect 23658 6196 23664 6208
rect 23716 6236 23722 6248
rect 24213 6239 24271 6245
rect 24213 6236 24225 6239
rect 23716 6208 24225 6236
rect 23716 6196 23722 6208
rect 24213 6205 24225 6208
rect 24259 6205 24271 6239
rect 24213 6199 24271 6205
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 24213 5899 24271 5905
rect 24213 5865 24225 5899
rect 24259 5896 24271 5899
rect 24854 5896 24860 5908
rect 24259 5868 24860 5896
rect 24259 5865 24271 5868
rect 24213 5859 24271 5865
rect 24854 5856 24860 5868
rect 24912 5856 24918 5908
rect 24026 5760 24032 5772
rect 23987 5732 24032 5760
rect 24026 5720 24032 5732
rect 24084 5720 24090 5772
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 24026 5352 24032 5364
rect 23987 5324 24032 5352
rect 24026 5312 24032 5324
rect 24084 5312 24090 5364
rect 24762 5352 24768 5364
rect 24723 5324 24768 5352
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 24578 5148 24584 5160
rect 24539 5120 24584 5148
rect 24578 5108 24584 5120
rect 24636 5148 24642 5160
rect 25133 5151 25191 5157
rect 25133 5148 25145 5151
rect 24636 5120 25145 5148
rect 24636 5108 24642 5120
rect 25133 5117 25145 5120
rect 25179 5117 25191 5151
rect 25133 5111 25191 5117
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 24762 4808 24768 4820
rect 24723 4780 24768 4808
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 24581 4675 24639 4681
rect 24581 4641 24593 4675
rect 24627 4672 24639 4675
rect 24670 4672 24676 4684
rect 24627 4644 24676 4672
rect 24627 4641 24639 4644
rect 24581 4635 24639 4641
rect 24670 4632 24676 4644
rect 24728 4632 24734 4684
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 24578 4196 24584 4208
rect 24539 4168 24584 4196
rect 24578 4156 24584 4168
rect 24636 4156 24642 4208
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 2314 3040 2320 3052
rect 2275 3012 2320 3040
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 2590 2913 2596 2916
rect 2225 2907 2283 2913
rect 2225 2873 2237 2907
rect 2271 2904 2283 2907
rect 2584 2904 2596 2913
rect 2271 2876 2596 2904
rect 2271 2873 2283 2876
rect 2225 2867 2283 2873
rect 2584 2867 2596 2876
rect 2590 2864 2596 2867
rect 2648 2864 2654 2916
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3697 2839 3755 2845
rect 3697 2836 3709 2839
rect 2832 2808 3709 2836
rect 2832 2796 2838 2808
rect 3697 2805 3709 2808
rect 3743 2805 3755 2839
rect 3697 2799 3755 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2314 2632 2320 2644
rect 2275 2604 2320 2632
rect 2314 2592 2320 2604
rect 2372 2592 2378 2644
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 3424 27344 3476 27396
rect 7196 27344 7248 27396
rect 3516 26324 3568 26376
rect 9220 26324 9272 26376
rect 3424 26256 3476 26308
rect 8116 26256 8168 26308
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 4896 25440 4948 25492
rect 7656 25440 7708 25492
rect 8116 25440 8168 25492
rect 1952 25372 2004 25424
rect 2044 25304 2096 25356
rect 2320 25304 2372 25356
rect 4620 25304 4672 25356
rect 5172 25347 5224 25356
rect 5172 25313 5181 25347
rect 5181 25313 5215 25347
rect 5215 25313 5224 25347
rect 5172 25304 5224 25313
rect 5080 25236 5132 25288
rect 6276 25372 6328 25424
rect 7104 25304 7156 25356
rect 9772 25347 9824 25356
rect 9772 25313 9781 25347
rect 9781 25313 9815 25347
rect 9815 25313 9824 25347
rect 9772 25304 9824 25313
rect 10876 25279 10928 25288
rect 10876 25245 10885 25279
rect 10885 25245 10919 25279
rect 10919 25245 10928 25279
rect 10876 25236 10928 25245
rect 2780 25168 2832 25220
rect 3516 25168 3568 25220
rect 7196 25168 7248 25220
rect 2872 25100 2924 25152
rect 3884 25100 3936 25152
rect 5540 25100 5592 25152
rect 11612 25100 11664 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 4896 24939 4948 24948
rect 4896 24905 4905 24939
rect 4905 24905 4939 24939
rect 4939 24905 4948 24939
rect 4896 24896 4948 24905
rect 5172 24896 5224 24948
rect 11612 24896 11664 24948
rect 2320 24828 2372 24880
rect 3240 24828 3292 24880
rect 3884 24803 3936 24812
rect 3884 24769 3893 24803
rect 3893 24769 3927 24803
rect 3927 24769 3936 24803
rect 3884 24760 3936 24769
rect 3976 24803 4028 24812
rect 3976 24769 3985 24803
rect 3985 24769 4019 24803
rect 4019 24769 4028 24803
rect 3976 24760 4028 24769
rect 5448 24760 5500 24812
rect 6276 24803 6328 24812
rect 6276 24769 6285 24803
rect 6285 24769 6319 24803
rect 6319 24769 6328 24803
rect 6276 24760 6328 24769
rect 8852 24803 8904 24812
rect 8852 24769 8861 24803
rect 8861 24769 8895 24803
rect 8895 24769 8904 24803
rect 8852 24760 8904 24769
rect 1676 24692 1728 24744
rect 3792 24735 3844 24744
rect 3792 24701 3801 24735
rect 3801 24701 3835 24735
rect 3835 24701 3844 24735
rect 3792 24692 3844 24701
rect 6828 24735 6880 24744
rect 6828 24701 6837 24735
rect 6837 24701 6871 24735
rect 6871 24701 6880 24735
rect 6828 24692 6880 24701
rect 7932 24735 7984 24744
rect 7932 24701 7941 24735
rect 7941 24701 7975 24735
rect 7975 24701 7984 24735
rect 11336 24803 11388 24812
rect 11336 24769 11345 24803
rect 11345 24769 11379 24803
rect 11379 24769 11388 24803
rect 11336 24760 11388 24769
rect 12992 24828 13044 24880
rect 12900 24803 12952 24812
rect 12900 24769 12909 24803
rect 12909 24769 12943 24803
rect 12943 24769 12952 24803
rect 12900 24760 12952 24769
rect 7932 24692 7984 24701
rect 12440 24692 12492 24744
rect 6552 24667 6604 24676
rect 6552 24633 6561 24667
rect 6561 24633 6595 24667
rect 6595 24633 6604 24667
rect 6552 24624 6604 24633
rect 12256 24624 12308 24676
rect 1400 24556 1452 24608
rect 2044 24599 2096 24608
rect 2044 24565 2053 24599
rect 2053 24565 2087 24599
rect 2087 24565 2096 24599
rect 2044 24556 2096 24565
rect 3424 24599 3476 24608
rect 3424 24565 3433 24599
rect 3433 24565 3467 24599
rect 3467 24565 3476 24599
rect 3424 24556 3476 24565
rect 4620 24556 4672 24608
rect 5172 24599 5224 24608
rect 5172 24565 5181 24599
rect 5181 24565 5215 24599
rect 5215 24565 5224 24599
rect 5172 24556 5224 24565
rect 7012 24599 7064 24608
rect 7012 24565 7021 24599
rect 7021 24565 7055 24599
rect 7055 24565 7064 24599
rect 7012 24556 7064 24565
rect 8208 24556 8260 24608
rect 9220 24599 9272 24608
rect 9220 24565 9229 24599
rect 9229 24565 9263 24599
rect 9263 24565 9272 24599
rect 9220 24556 9272 24565
rect 9772 24599 9824 24608
rect 9772 24565 9781 24599
rect 9781 24565 9815 24599
rect 9815 24565 9824 24599
rect 9772 24556 9824 24565
rect 10692 24599 10744 24608
rect 10692 24565 10701 24599
rect 10701 24565 10735 24599
rect 10735 24565 10744 24599
rect 10692 24556 10744 24565
rect 11612 24556 11664 24608
rect 12808 24556 12860 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 3976 24352 4028 24404
rect 6552 24352 6604 24404
rect 8116 24395 8168 24404
rect 8116 24361 8125 24395
rect 8125 24361 8159 24395
rect 8159 24361 8168 24395
rect 8116 24352 8168 24361
rect 10692 24352 10744 24404
rect 12808 24352 12860 24404
rect 14188 24395 14240 24404
rect 14188 24361 14197 24395
rect 14197 24361 14231 24395
rect 14231 24361 14240 24395
rect 14188 24352 14240 24361
rect 16764 24395 16816 24404
rect 16764 24361 16773 24395
rect 16773 24361 16807 24395
rect 16807 24361 16816 24395
rect 16764 24352 16816 24361
rect 17868 24395 17920 24404
rect 17868 24361 17877 24395
rect 17877 24361 17911 24395
rect 17911 24361 17920 24395
rect 17868 24352 17920 24361
rect 19064 24395 19116 24404
rect 19064 24361 19073 24395
rect 19073 24361 19107 24395
rect 19107 24361 19116 24395
rect 19064 24352 19116 24361
rect 22468 24352 22520 24404
rect 1860 24327 1912 24336
rect 1860 24293 1869 24327
rect 1869 24293 1903 24327
rect 1903 24293 1912 24327
rect 1860 24284 1912 24293
rect 3792 24284 3844 24336
rect 1584 24259 1636 24268
rect 1584 24225 1593 24259
rect 1593 24225 1627 24259
rect 1627 24225 1636 24259
rect 1584 24216 1636 24225
rect 2964 24216 3016 24268
rect 3884 24216 3936 24268
rect 6000 24284 6052 24336
rect 5448 24259 5500 24268
rect 5448 24225 5482 24259
rect 5482 24225 5500 24259
rect 5448 24216 5500 24225
rect 7288 24216 7340 24268
rect 8024 24259 8076 24268
rect 8024 24225 8033 24259
rect 8033 24225 8067 24259
rect 8067 24225 8076 24259
rect 8024 24216 8076 24225
rect 11336 24216 11388 24268
rect 12716 24216 12768 24268
rect 16764 24216 16816 24268
rect 17684 24259 17736 24268
rect 17684 24225 17693 24259
rect 17693 24225 17727 24259
rect 17727 24225 17736 24259
rect 17684 24216 17736 24225
rect 18880 24259 18932 24268
rect 18880 24225 18889 24259
rect 18889 24225 18923 24259
rect 18923 24225 18932 24259
rect 18880 24216 18932 24225
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 8208 24191 8260 24200
rect 8208 24157 8217 24191
rect 8217 24157 8251 24191
rect 8251 24157 8260 24191
rect 10140 24191 10192 24200
rect 8208 24148 8260 24157
rect 10140 24157 10149 24191
rect 10149 24157 10183 24191
rect 10183 24157 10192 24191
rect 10140 24148 10192 24157
rect 12348 24080 12400 24132
rect 3056 24055 3108 24064
rect 3056 24021 3065 24055
rect 3065 24021 3099 24055
rect 3099 24021 3108 24055
rect 3056 24012 3108 24021
rect 4252 24055 4304 24064
rect 4252 24021 4261 24055
rect 4261 24021 4295 24055
rect 4295 24021 4304 24055
rect 4252 24012 4304 24021
rect 5080 24012 5132 24064
rect 7104 24055 7156 24064
rect 7104 24021 7113 24055
rect 7113 24021 7147 24055
rect 7147 24021 7156 24055
rect 7104 24012 7156 24021
rect 11520 24055 11572 24064
rect 11520 24021 11529 24055
rect 11529 24021 11563 24055
rect 11563 24021 11572 24055
rect 11520 24012 11572 24021
rect 12440 24055 12492 24064
rect 12440 24021 12449 24055
rect 12449 24021 12483 24055
rect 12483 24021 12492 24055
rect 13728 24055 13780 24064
rect 12440 24012 12492 24021
rect 13728 24021 13737 24055
rect 13737 24021 13771 24055
rect 13771 24021 13780 24055
rect 13728 24012 13780 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 2044 23715 2096 23724
rect 2044 23681 2053 23715
rect 2053 23681 2087 23715
rect 2087 23681 2096 23715
rect 2044 23672 2096 23681
rect 3424 23808 3476 23860
rect 7288 23851 7340 23860
rect 7288 23817 7297 23851
rect 7297 23817 7331 23851
rect 7331 23817 7340 23851
rect 7288 23808 7340 23817
rect 8116 23808 8168 23860
rect 12808 23808 12860 23860
rect 16488 23808 16540 23860
rect 17868 23808 17920 23860
rect 19248 23808 19300 23860
rect 20260 23808 20312 23860
rect 20444 23851 20496 23860
rect 20444 23817 20453 23851
rect 20453 23817 20487 23851
rect 20487 23817 20496 23851
rect 20444 23808 20496 23817
rect 21548 23851 21600 23860
rect 21548 23817 21557 23851
rect 21557 23817 21591 23851
rect 21591 23817 21600 23851
rect 21548 23808 21600 23817
rect 12716 23783 12768 23792
rect 12716 23749 12725 23783
rect 12725 23749 12759 23783
rect 12759 23749 12768 23783
rect 12716 23740 12768 23749
rect 10692 23715 10744 23724
rect 3792 23647 3844 23656
rect 3792 23613 3801 23647
rect 3801 23613 3835 23647
rect 3835 23613 3844 23647
rect 3792 23604 3844 23613
rect 10692 23681 10701 23715
rect 10701 23681 10735 23715
rect 10735 23681 10744 23715
rect 10692 23672 10744 23681
rect 10784 23715 10836 23724
rect 10784 23681 10793 23715
rect 10793 23681 10827 23715
rect 10827 23681 10836 23715
rect 10784 23672 10836 23681
rect 11520 23672 11572 23724
rect 5080 23604 5132 23656
rect 7012 23604 7064 23656
rect 10876 23604 10928 23656
rect 12624 23604 12676 23656
rect 18328 23672 18380 23724
rect 18880 23672 18932 23724
rect 13728 23604 13780 23656
rect 15476 23604 15528 23656
rect 16120 23604 16172 23656
rect 19156 23647 19208 23656
rect 2504 23536 2556 23588
rect 3884 23536 3936 23588
rect 4804 23536 4856 23588
rect 5356 23536 5408 23588
rect 5448 23536 5500 23588
rect 2228 23468 2280 23520
rect 2964 23468 3016 23520
rect 4160 23468 4212 23520
rect 6000 23468 6052 23520
rect 8208 23536 8260 23588
rect 16764 23536 16816 23588
rect 19156 23613 19165 23647
rect 19165 23613 19199 23647
rect 19199 23613 19208 23647
rect 19156 23604 19208 23613
rect 20260 23647 20312 23656
rect 20260 23613 20269 23647
rect 20269 23613 20303 23647
rect 20303 23613 20312 23647
rect 20260 23604 20312 23613
rect 21364 23647 21416 23656
rect 21364 23613 21373 23647
rect 21373 23613 21407 23647
rect 21407 23613 21416 23647
rect 21364 23604 21416 23613
rect 23480 23536 23532 23588
rect 24768 23536 24820 23588
rect 9680 23468 9732 23520
rect 11336 23511 11388 23520
rect 11336 23477 11345 23511
rect 11345 23477 11379 23511
rect 11379 23477 11388 23511
rect 11336 23468 11388 23477
rect 16580 23468 16632 23520
rect 17684 23511 17736 23520
rect 17684 23477 17693 23511
rect 17693 23477 17727 23511
rect 17727 23477 17736 23511
rect 17684 23468 17736 23477
rect 18604 23511 18656 23520
rect 18604 23477 18613 23511
rect 18613 23477 18647 23511
rect 18647 23477 18656 23511
rect 18604 23468 18656 23477
rect 20904 23468 20956 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 7012 23307 7064 23316
rect 7012 23273 7021 23307
rect 7021 23273 7055 23307
rect 7055 23273 7064 23307
rect 7012 23264 7064 23273
rect 8208 23264 8260 23316
rect 13820 23264 13872 23316
rect 16672 23307 16724 23316
rect 16672 23273 16681 23307
rect 16681 23273 16715 23307
rect 16715 23273 16724 23307
rect 16672 23264 16724 23273
rect 19984 23264 20036 23316
rect 1860 23239 1912 23248
rect 1860 23205 1869 23239
rect 1869 23205 1903 23239
rect 1903 23205 1912 23239
rect 1860 23196 1912 23205
rect 4160 23196 4212 23248
rect 1584 23171 1636 23180
rect 1584 23137 1593 23171
rect 1593 23137 1627 23171
rect 1627 23137 1636 23171
rect 1584 23128 1636 23137
rect 3424 23128 3476 23180
rect 3792 23171 3844 23180
rect 3792 23137 3801 23171
rect 3801 23137 3835 23171
rect 3835 23137 3844 23171
rect 3792 23128 3844 23137
rect 9588 23196 9640 23248
rect 10784 23196 10836 23248
rect 12992 23239 13044 23248
rect 12992 23205 13026 23239
rect 13026 23205 13044 23239
rect 12992 23196 13044 23205
rect 7380 23171 7432 23180
rect 7380 23137 7414 23171
rect 7414 23137 7432 23171
rect 7380 23128 7432 23137
rect 10140 23128 10192 23180
rect 15568 23171 15620 23180
rect 15568 23137 15602 23171
rect 15602 23137 15620 23171
rect 15568 23128 15620 23137
rect 19432 23171 19484 23180
rect 19432 23137 19441 23171
rect 19441 23137 19475 23171
rect 19475 23137 19484 23171
rect 19432 23128 19484 23137
rect 15292 23103 15344 23112
rect 15292 23069 15301 23103
rect 15301 23069 15335 23103
rect 15335 23069 15344 23103
rect 15292 23060 15344 23069
rect 2412 22967 2464 22976
rect 2412 22933 2421 22967
rect 2421 22933 2455 22967
rect 2455 22933 2464 22967
rect 2412 22924 2464 22933
rect 2872 22924 2924 22976
rect 3240 22924 3292 22976
rect 5264 22924 5316 22976
rect 10692 22924 10744 22976
rect 12624 22967 12676 22976
rect 12624 22933 12633 22967
rect 12633 22933 12667 22967
rect 12667 22933 12676 22967
rect 12624 22924 12676 22933
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1584 22720 1636 22772
rect 2596 22720 2648 22772
rect 4160 22763 4212 22772
rect 4160 22729 4169 22763
rect 4169 22729 4203 22763
rect 4203 22729 4212 22763
rect 4160 22720 4212 22729
rect 5172 22763 5224 22772
rect 5172 22729 5181 22763
rect 5181 22729 5215 22763
rect 5215 22729 5224 22763
rect 5172 22720 5224 22729
rect 9588 22763 9640 22772
rect 9588 22729 9597 22763
rect 9597 22729 9631 22763
rect 9631 22729 9640 22763
rect 9588 22720 9640 22729
rect 12992 22763 13044 22772
rect 12992 22729 13001 22763
rect 13001 22729 13035 22763
rect 13035 22729 13044 22763
rect 12992 22720 13044 22729
rect 2504 22584 2556 22636
rect 3240 22627 3292 22636
rect 3240 22593 3249 22627
rect 3249 22593 3283 22627
rect 3283 22593 3292 22627
rect 3240 22584 3292 22593
rect 4068 22584 4120 22636
rect 5448 22584 5500 22636
rect 7012 22584 7064 22636
rect 10692 22627 10744 22636
rect 10692 22593 10701 22627
rect 10701 22593 10735 22627
rect 10735 22593 10744 22627
rect 10692 22584 10744 22593
rect 12716 22584 12768 22636
rect 2412 22516 2464 22568
rect 5540 22559 5592 22568
rect 5540 22525 5549 22559
rect 5549 22525 5583 22559
rect 5583 22525 5592 22559
rect 5540 22516 5592 22525
rect 8024 22516 8076 22568
rect 10876 22516 10928 22568
rect 10968 22516 11020 22568
rect 12624 22516 12676 22568
rect 13636 22516 13688 22568
rect 15292 22516 15344 22568
rect 3148 22491 3200 22500
rect 3148 22457 3157 22491
rect 3157 22457 3191 22491
rect 3191 22457 3200 22491
rect 3148 22448 3200 22457
rect 6828 22448 6880 22500
rect 6000 22380 6052 22432
rect 7012 22380 7064 22432
rect 9864 22448 9916 22500
rect 7380 22380 7432 22432
rect 9956 22380 10008 22432
rect 13544 22423 13596 22432
rect 13544 22389 13553 22423
rect 13553 22389 13587 22423
rect 13587 22389 13596 22423
rect 13544 22380 13596 22389
rect 13820 22380 13872 22432
rect 15568 22380 15620 22432
rect 19432 22423 19484 22432
rect 19432 22389 19441 22423
rect 19441 22389 19475 22423
rect 19475 22389 19484 22423
rect 19432 22380 19484 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2596 22219 2648 22228
rect 2596 22185 2605 22219
rect 2605 22185 2639 22219
rect 2639 22185 2648 22219
rect 2596 22176 2648 22185
rect 3240 22176 3292 22228
rect 9864 22176 9916 22228
rect 15384 22176 15436 22228
rect 16304 22219 16356 22228
rect 16304 22185 16313 22219
rect 16313 22185 16347 22219
rect 16347 22185 16356 22219
rect 16304 22176 16356 22185
rect 3792 22151 3844 22160
rect 3792 22117 3801 22151
rect 3801 22117 3835 22151
rect 3835 22117 3844 22151
rect 3792 22108 3844 22117
rect 8208 22151 8260 22160
rect 8208 22117 8217 22151
rect 8217 22117 8251 22151
rect 8251 22117 8260 22151
rect 8208 22108 8260 22117
rect 10692 22108 10744 22160
rect 13636 22108 13688 22160
rect 2320 22040 2372 22092
rect 2780 22083 2832 22092
rect 2780 22049 2789 22083
rect 2789 22049 2823 22083
rect 2823 22049 2832 22083
rect 2780 22040 2832 22049
rect 4436 22083 4488 22092
rect 4436 22049 4445 22083
rect 4445 22049 4479 22083
rect 4479 22049 4488 22083
rect 4436 22040 4488 22049
rect 4528 22083 4580 22092
rect 4528 22049 4537 22083
rect 4537 22049 4571 22083
rect 4571 22049 4580 22083
rect 4528 22040 4580 22049
rect 5448 22040 5500 22092
rect 6184 22040 6236 22092
rect 8760 22040 8812 22092
rect 10140 22040 10192 22092
rect 10968 22040 11020 22092
rect 13176 22083 13228 22092
rect 13176 22049 13185 22083
rect 13185 22049 13219 22083
rect 13219 22049 13228 22083
rect 13176 22040 13228 22049
rect 15200 22108 15252 22160
rect 2412 21972 2464 22024
rect 5172 21972 5224 22024
rect 6736 22015 6788 22024
rect 6736 21981 6745 22015
rect 6745 21981 6779 22015
rect 6779 21981 6788 22015
rect 6736 21972 6788 21981
rect 7012 21972 7064 22024
rect 8024 21972 8076 22024
rect 12900 21972 12952 22024
rect 2320 21947 2372 21956
rect 2320 21913 2329 21947
rect 2329 21913 2363 21947
rect 2363 21913 2372 21947
rect 2320 21904 2372 21913
rect 2964 21947 3016 21956
rect 2964 21913 2973 21947
rect 2973 21913 3007 21947
rect 3007 21913 3016 21947
rect 2964 21904 3016 21913
rect 6920 21904 6972 21956
rect 12256 21904 12308 21956
rect 13728 21972 13780 22024
rect 3424 21879 3476 21888
rect 3424 21845 3433 21879
rect 3433 21845 3467 21879
rect 3467 21845 3476 21879
rect 3424 21836 3476 21845
rect 5172 21836 5224 21888
rect 6000 21879 6052 21888
rect 6000 21845 6009 21879
rect 6009 21845 6043 21879
rect 6043 21845 6052 21879
rect 6000 21836 6052 21845
rect 6276 21879 6328 21888
rect 6276 21845 6285 21879
rect 6285 21845 6319 21879
rect 6319 21845 6328 21879
rect 6276 21836 6328 21845
rect 7564 21879 7616 21888
rect 7564 21845 7573 21879
rect 7573 21845 7607 21879
rect 7607 21845 7616 21879
rect 7564 21836 7616 21845
rect 10140 21836 10192 21888
rect 12808 21879 12860 21888
rect 12808 21845 12817 21879
rect 12817 21845 12851 21879
rect 12851 21845 12860 21879
rect 12808 21836 12860 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 2780 21675 2832 21684
rect 2780 21641 2789 21675
rect 2789 21641 2823 21675
rect 2823 21641 2832 21675
rect 2780 21632 2832 21641
rect 3516 21632 3568 21684
rect 4160 21632 4212 21684
rect 4528 21632 4580 21684
rect 5264 21675 5316 21684
rect 5264 21641 5273 21675
rect 5273 21641 5307 21675
rect 5307 21641 5316 21675
rect 5264 21632 5316 21641
rect 8760 21632 8812 21684
rect 9496 21675 9548 21684
rect 9496 21641 9505 21675
rect 9505 21641 9539 21675
rect 9539 21641 9548 21675
rect 9496 21632 9548 21641
rect 10692 21632 10744 21684
rect 6736 21564 6788 21616
rect 8300 21564 8352 21616
rect 8852 21607 8904 21616
rect 8852 21573 8861 21607
rect 8861 21573 8895 21607
rect 8895 21573 8904 21607
rect 8852 21564 8904 21573
rect 1676 21539 1728 21548
rect 1676 21505 1685 21539
rect 1685 21505 1719 21539
rect 1719 21505 1728 21539
rect 1676 21496 1728 21505
rect 2320 21428 2372 21480
rect 7932 21539 7984 21548
rect 7932 21505 7941 21539
rect 7941 21505 7975 21539
rect 7975 21505 7984 21539
rect 7932 21496 7984 21505
rect 8208 21496 8260 21548
rect 9956 21539 10008 21548
rect 9956 21505 9965 21539
rect 9965 21505 9999 21539
rect 9999 21505 10008 21539
rect 9956 21496 10008 21505
rect 10140 21539 10192 21548
rect 10140 21505 10149 21539
rect 10149 21505 10183 21539
rect 10183 21505 10192 21539
rect 10140 21496 10192 21505
rect 11244 21539 11296 21548
rect 11244 21505 11253 21539
rect 11253 21505 11287 21539
rect 11287 21505 11296 21539
rect 11244 21496 11296 21505
rect 5264 21428 5316 21480
rect 3792 21360 3844 21412
rect 5172 21360 5224 21412
rect 7564 21428 7616 21480
rect 12348 21632 12400 21684
rect 13176 21675 13228 21684
rect 13176 21641 13185 21675
rect 13185 21641 13219 21675
rect 13219 21641 13228 21675
rect 13176 21632 13228 21641
rect 12256 21607 12308 21616
rect 12256 21573 12265 21607
rect 12265 21573 12299 21607
rect 12299 21573 12308 21607
rect 12256 21564 12308 21573
rect 13636 21496 13688 21548
rect 7012 21360 7064 21412
rect 10692 21360 10744 21412
rect 15200 21360 15252 21412
rect 23572 21360 23624 21412
rect 24216 21360 24268 21412
rect 24860 21360 24912 21412
rect 25964 21360 26016 21412
rect 5540 21335 5592 21344
rect 5540 21301 5549 21335
rect 5549 21301 5583 21335
rect 5583 21301 5592 21335
rect 5540 21292 5592 21301
rect 6184 21292 6236 21344
rect 13544 21292 13596 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 2412 21131 2464 21140
rect 2412 21097 2421 21131
rect 2421 21097 2455 21131
rect 2455 21097 2464 21131
rect 2412 21088 2464 21097
rect 3792 21088 3844 21140
rect 6736 21088 6788 21140
rect 8024 21088 8076 21140
rect 12900 21131 12952 21140
rect 12900 21097 12909 21131
rect 12909 21097 12943 21131
rect 12943 21097 12952 21131
rect 12900 21088 12952 21097
rect 13360 21131 13412 21140
rect 13360 21097 13369 21131
rect 13369 21097 13403 21131
rect 13403 21097 13412 21131
rect 13360 21088 13412 21097
rect 13636 21088 13688 21140
rect 13820 21088 13872 21140
rect 15292 21131 15344 21140
rect 15292 21097 15301 21131
rect 15301 21097 15335 21131
rect 15335 21097 15344 21131
rect 15292 21088 15344 21097
rect 1952 21020 2004 21072
rect 5264 21020 5316 21072
rect 10140 21020 10192 21072
rect 2688 20952 2740 21004
rect 3056 20952 3108 21004
rect 5448 20952 5500 21004
rect 6828 20952 6880 21004
rect 7012 20995 7064 21004
rect 7012 20961 7046 20995
rect 7046 20961 7064 20995
rect 7012 20952 7064 20961
rect 12440 20952 12492 21004
rect 13176 20952 13228 21004
rect 5172 20927 5224 20936
rect 5172 20893 5181 20927
rect 5181 20893 5215 20927
rect 5215 20893 5224 20927
rect 5172 20884 5224 20893
rect 6000 20927 6052 20936
rect 6000 20893 6009 20927
rect 6009 20893 6043 20927
rect 6043 20893 6052 20927
rect 6736 20927 6788 20936
rect 6000 20884 6052 20893
rect 3976 20816 4028 20868
rect 4436 20816 4488 20868
rect 4896 20816 4948 20868
rect 6736 20893 6745 20927
rect 6745 20893 6779 20927
rect 6779 20893 6788 20927
rect 6736 20884 6788 20893
rect 10048 20927 10100 20936
rect 10048 20893 10057 20927
rect 10057 20893 10091 20927
rect 10091 20893 10100 20927
rect 10048 20884 10100 20893
rect 12992 20884 13044 20936
rect 13544 20884 13596 20936
rect 12532 20859 12584 20868
rect 12532 20825 12541 20859
rect 12541 20825 12575 20859
rect 12575 20825 12584 20859
rect 12532 20816 12584 20825
rect 13820 20816 13872 20868
rect 3148 20748 3200 20800
rect 4528 20748 4580 20800
rect 8208 20748 8260 20800
rect 9312 20748 9364 20800
rect 11060 20748 11112 20800
rect 14096 20748 14148 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 4068 20544 4120 20596
rect 5172 20544 5224 20596
rect 5540 20544 5592 20596
rect 6000 20587 6052 20596
rect 6000 20553 6009 20587
rect 6009 20553 6043 20587
rect 6043 20553 6052 20587
rect 6000 20544 6052 20553
rect 7012 20544 7064 20596
rect 9036 20587 9088 20596
rect 9036 20553 9045 20587
rect 9045 20553 9079 20587
rect 9079 20553 9088 20587
rect 9036 20544 9088 20553
rect 10140 20544 10192 20596
rect 11888 20587 11940 20596
rect 11888 20553 11897 20587
rect 11897 20553 11931 20587
rect 11931 20553 11940 20587
rect 11888 20544 11940 20553
rect 12348 20544 12400 20596
rect 13360 20544 13412 20596
rect 15292 20544 15344 20596
rect 5264 20476 5316 20528
rect 6460 20476 6512 20528
rect 2320 20451 2372 20460
rect 2320 20417 2329 20451
rect 2329 20417 2363 20451
rect 2363 20417 2372 20451
rect 2320 20408 2372 20417
rect 1768 20383 1820 20392
rect 1768 20349 1777 20383
rect 1777 20349 1811 20383
rect 1811 20349 1820 20383
rect 1768 20340 1820 20349
rect 3792 20340 3844 20392
rect 6736 20340 6788 20392
rect 4068 20272 4120 20324
rect 9036 20340 9088 20392
rect 7104 20315 7156 20324
rect 7104 20281 7138 20315
rect 7138 20281 7156 20315
rect 7104 20272 7156 20281
rect 8208 20272 8260 20324
rect 9956 20408 10008 20460
rect 10968 20408 11020 20460
rect 11152 20408 11204 20460
rect 12348 20408 12400 20460
rect 13820 20451 13872 20460
rect 13820 20417 13829 20451
rect 13829 20417 13863 20451
rect 13863 20417 13872 20451
rect 13820 20408 13872 20417
rect 10876 20340 10928 20392
rect 12808 20340 12860 20392
rect 13360 20340 13412 20392
rect 10692 20272 10744 20324
rect 12716 20315 12768 20324
rect 12716 20281 12725 20315
rect 12725 20281 12759 20315
rect 12759 20281 12768 20315
rect 12716 20272 12768 20281
rect 14096 20315 14148 20324
rect 14096 20281 14130 20315
rect 14130 20281 14148 20315
rect 14096 20272 14148 20281
rect 14188 20272 14240 20324
rect 2688 20247 2740 20256
rect 2688 20213 2697 20247
rect 2697 20213 2731 20247
rect 2731 20213 2740 20247
rect 2688 20204 2740 20213
rect 3056 20247 3108 20256
rect 3056 20213 3065 20247
rect 3065 20213 3099 20247
rect 3099 20213 3108 20247
rect 3056 20204 3108 20213
rect 3516 20204 3568 20256
rect 9588 20247 9640 20256
rect 9588 20213 9597 20247
rect 9597 20213 9631 20247
rect 9631 20213 9640 20247
rect 9588 20204 9640 20213
rect 11336 20247 11388 20256
rect 11336 20213 11345 20247
rect 11345 20213 11379 20247
rect 11379 20213 11388 20247
rect 11336 20204 11388 20213
rect 13176 20204 13228 20256
rect 16304 20247 16356 20256
rect 16304 20213 16313 20247
rect 16313 20213 16347 20247
rect 16347 20213 16356 20247
rect 16304 20204 16356 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 7104 20000 7156 20052
rect 8760 20000 8812 20052
rect 9588 20000 9640 20052
rect 12992 20043 13044 20052
rect 12992 20009 13001 20043
rect 13001 20009 13035 20043
rect 13035 20009 13044 20043
rect 12992 20000 13044 20009
rect 16028 20000 16080 20052
rect 2228 19932 2280 19984
rect 5172 19932 5224 19984
rect 9036 19975 9088 19984
rect 9036 19941 9045 19975
rect 9045 19941 9079 19975
rect 9079 19941 9088 19975
rect 9036 19932 9088 19941
rect 9956 19975 10008 19984
rect 9956 19941 9965 19975
rect 9965 19941 9999 19975
rect 9999 19941 10008 19975
rect 9956 19932 10008 19941
rect 13728 19932 13780 19984
rect 14188 19975 14240 19984
rect 14188 19941 14197 19975
rect 14197 19941 14231 19975
rect 14231 19941 14240 19975
rect 14188 19932 14240 19941
rect 15660 19975 15712 19984
rect 15660 19941 15669 19975
rect 15669 19941 15703 19975
rect 15703 19941 15712 19975
rect 15660 19932 15712 19941
rect 3424 19864 3476 19916
rect 3976 19864 4028 19916
rect 4436 19864 4488 19916
rect 5448 19864 5500 19916
rect 2320 19839 2372 19848
rect 2320 19805 2329 19839
rect 2329 19805 2363 19839
rect 2363 19805 2372 19839
rect 2320 19796 2372 19805
rect 7012 19864 7064 19916
rect 8392 19907 8444 19916
rect 8392 19873 8401 19907
rect 8401 19873 8435 19907
rect 8435 19873 8444 19907
rect 8392 19864 8444 19873
rect 10048 19907 10100 19916
rect 10048 19873 10057 19907
rect 10057 19873 10091 19907
rect 10091 19873 10100 19907
rect 10048 19864 10100 19873
rect 11152 19864 11204 19916
rect 12808 19864 12860 19916
rect 13544 19907 13596 19916
rect 13544 19873 13553 19907
rect 13553 19873 13587 19907
rect 13587 19873 13596 19907
rect 13544 19864 13596 19873
rect 7932 19796 7984 19848
rect 8668 19839 8720 19848
rect 8668 19805 8677 19839
rect 8677 19805 8711 19839
rect 8711 19805 8720 19839
rect 8668 19796 8720 19805
rect 8024 19771 8076 19780
rect 8024 19737 8033 19771
rect 8033 19737 8067 19771
rect 8067 19737 8076 19771
rect 8024 19728 8076 19737
rect 2504 19660 2556 19712
rect 3056 19660 3108 19712
rect 3424 19703 3476 19712
rect 3424 19669 3433 19703
rect 3433 19669 3467 19703
rect 3467 19669 3476 19703
rect 3424 19660 3476 19669
rect 3976 19660 4028 19712
rect 6184 19660 6236 19712
rect 6920 19660 6972 19712
rect 7380 19703 7432 19712
rect 7380 19669 7389 19703
rect 7389 19669 7423 19703
rect 7423 19669 7432 19703
rect 7380 19660 7432 19669
rect 14096 19796 14148 19848
rect 14648 19796 14700 19848
rect 15292 19796 15344 19848
rect 16304 19796 16356 19848
rect 15292 19703 15344 19712
rect 15292 19669 15301 19703
rect 15301 19669 15335 19703
rect 15335 19669 15344 19703
rect 15292 19660 15344 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 4068 19499 4120 19508
rect 4068 19465 4077 19499
rect 4077 19465 4111 19499
rect 4111 19465 4120 19499
rect 4068 19456 4120 19465
rect 5172 19499 5224 19508
rect 5172 19465 5181 19499
rect 5181 19465 5215 19499
rect 5215 19465 5224 19499
rect 5172 19456 5224 19465
rect 5448 19499 5500 19508
rect 5448 19465 5457 19499
rect 5457 19465 5491 19499
rect 5491 19465 5500 19499
rect 5448 19456 5500 19465
rect 9312 19499 9364 19508
rect 9312 19465 9321 19499
rect 9321 19465 9355 19499
rect 9355 19465 9364 19499
rect 9312 19456 9364 19465
rect 9956 19456 10008 19508
rect 11612 19456 11664 19508
rect 11888 19456 11940 19508
rect 12808 19499 12860 19508
rect 12808 19465 12817 19499
rect 12817 19465 12851 19499
rect 12851 19465 12860 19499
rect 12808 19456 12860 19465
rect 13636 19456 13688 19508
rect 14648 19499 14700 19508
rect 14648 19465 14657 19499
rect 14657 19465 14691 19499
rect 14691 19465 14700 19499
rect 14648 19456 14700 19465
rect 15660 19456 15712 19508
rect 16304 19499 16356 19508
rect 16304 19465 16313 19499
rect 16313 19465 16347 19499
rect 16347 19465 16356 19499
rect 16304 19456 16356 19465
rect 2596 19363 2648 19372
rect 2596 19329 2605 19363
rect 2605 19329 2639 19363
rect 2639 19329 2648 19363
rect 2596 19320 2648 19329
rect 6092 19320 6144 19372
rect 7932 19363 7984 19372
rect 7932 19329 7941 19363
rect 7941 19329 7975 19363
rect 7975 19329 7984 19363
rect 7932 19320 7984 19329
rect 4528 19295 4580 19304
rect 4528 19261 4537 19295
rect 4537 19261 4571 19295
rect 4571 19261 4580 19295
rect 4528 19252 4580 19261
rect 1400 19184 1452 19236
rect 2964 19184 3016 19236
rect 8668 19252 8720 19304
rect 6276 19227 6328 19236
rect 2044 19159 2096 19168
rect 2044 19125 2053 19159
rect 2053 19125 2087 19159
rect 2087 19125 2096 19159
rect 2044 19116 2096 19125
rect 2504 19159 2556 19168
rect 2504 19125 2513 19159
rect 2513 19125 2547 19159
rect 2547 19125 2556 19159
rect 2504 19116 2556 19125
rect 3792 19116 3844 19168
rect 4160 19116 4212 19168
rect 6276 19193 6285 19227
rect 6285 19193 6319 19227
rect 6319 19193 6328 19227
rect 6276 19184 6328 19193
rect 6644 19159 6696 19168
rect 6644 19125 6653 19159
rect 6653 19125 6687 19159
rect 6687 19125 6696 19159
rect 6644 19116 6696 19125
rect 6828 19159 6880 19168
rect 6828 19125 6837 19159
rect 6837 19125 6871 19159
rect 6871 19125 6880 19159
rect 6828 19116 6880 19125
rect 8208 19116 8260 19168
rect 10140 19116 10192 19168
rect 11888 19295 11940 19304
rect 11888 19261 11897 19295
rect 11897 19261 11931 19295
rect 11931 19261 11940 19295
rect 11888 19252 11940 19261
rect 13360 19252 13412 19304
rect 15568 19252 15620 19304
rect 11152 19184 11204 19236
rect 11980 19184 12032 19236
rect 13912 19184 13964 19236
rect 15936 19159 15988 19168
rect 15936 19125 15945 19159
rect 15945 19125 15979 19159
rect 15979 19125 15988 19159
rect 15936 19116 15988 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1400 18955 1452 18964
rect 1400 18921 1409 18955
rect 1409 18921 1443 18955
rect 1443 18921 1452 18955
rect 1400 18912 1452 18921
rect 4436 18955 4488 18964
rect 4436 18921 4445 18955
rect 4445 18921 4479 18955
rect 4479 18921 4488 18955
rect 4436 18912 4488 18921
rect 4712 18912 4764 18964
rect 5540 18955 5592 18964
rect 5540 18921 5549 18955
rect 5549 18921 5583 18955
rect 5583 18921 5592 18955
rect 6092 18955 6144 18964
rect 5540 18912 5592 18921
rect 6092 18921 6101 18955
rect 6101 18921 6135 18955
rect 6135 18921 6144 18955
rect 6092 18912 6144 18921
rect 8760 18955 8812 18964
rect 8760 18921 8769 18955
rect 8769 18921 8803 18955
rect 8803 18921 8812 18955
rect 8760 18912 8812 18921
rect 13912 18955 13964 18964
rect 13912 18921 13921 18955
rect 13921 18921 13955 18955
rect 13955 18921 13964 18955
rect 13912 18912 13964 18921
rect 16028 18955 16080 18964
rect 16028 18921 16037 18955
rect 16037 18921 16071 18955
rect 16071 18921 16080 18955
rect 16028 18912 16080 18921
rect 4252 18844 4304 18896
rect 5264 18844 5316 18896
rect 6000 18844 6052 18896
rect 8668 18844 8720 18896
rect 12532 18844 12584 18896
rect 15568 18887 15620 18896
rect 15568 18853 15577 18887
rect 15577 18853 15611 18887
rect 15611 18853 15620 18887
rect 15568 18844 15620 18853
rect 2780 18819 2832 18828
rect 2780 18785 2789 18819
rect 2789 18785 2823 18819
rect 2823 18785 2832 18819
rect 2780 18776 2832 18785
rect 2872 18751 2924 18760
rect 2872 18717 2881 18751
rect 2881 18717 2915 18751
rect 2915 18717 2924 18751
rect 2872 18708 2924 18717
rect 2964 18751 3016 18760
rect 2964 18717 2973 18751
rect 2973 18717 3007 18751
rect 3007 18717 3016 18751
rect 2964 18708 3016 18717
rect 7656 18819 7708 18828
rect 7656 18785 7665 18819
rect 7665 18785 7699 18819
rect 7699 18785 7708 18819
rect 7656 18776 7708 18785
rect 7932 18776 7984 18828
rect 11336 18819 11388 18828
rect 4620 18751 4672 18760
rect 4620 18717 4629 18751
rect 4629 18717 4663 18751
rect 4663 18717 4672 18751
rect 4620 18708 4672 18717
rect 6368 18751 6420 18760
rect 6368 18717 6377 18751
rect 6377 18717 6411 18751
rect 6411 18717 6420 18751
rect 6368 18708 6420 18717
rect 8208 18708 8260 18760
rect 9864 18751 9916 18760
rect 9864 18717 9873 18751
rect 9873 18717 9907 18751
rect 9907 18717 9916 18751
rect 9864 18708 9916 18717
rect 4068 18683 4120 18692
rect 4068 18649 4077 18683
rect 4077 18649 4111 18683
rect 4111 18649 4120 18683
rect 4068 18640 4120 18649
rect 5632 18640 5684 18692
rect 7288 18683 7340 18692
rect 7288 18649 7297 18683
rect 7297 18649 7331 18683
rect 7331 18649 7340 18683
rect 7288 18640 7340 18649
rect 11336 18785 11345 18819
rect 11345 18785 11379 18819
rect 11379 18785 11388 18819
rect 11336 18776 11388 18785
rect 15292 18819 15344 18828
rect 15292 18785 15301 18819
rect 15301 18785 15335 18819
rect 15335 18785 15344 18819
rect 15292 18776 15344 18785
rect 11428 18751 11480 18760
rect 11428 18717 11437 18751
rect 11437 18717 11471 18751
rect 11471 18717 11480 18751
rect 11428 18708 11480 18717
rect 11980 18708 12032 18760
rect 2044 18572 2096 18624
rect 2596 18572 2648 18624
rect 2964 18572 3016 18624
rect 7196 18572 7248 18624
rect 9312 18615 9364 18624
rect 9312 18581 9321 18615
rect 9321 18581 9355 18615
rect 9355 18581 9364 18615
rect 9312 18572 9364 18581
rect 10876 18615 10928 18624
rect 10876 18581 10885 18615
rect 10885 18581 10919 18615
rect 10919 18581 10928 18615
rect 10876 18572 10928 18581
rect 12164 18572 12216 18624
rect 12532 18572 12584 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 6000 18368 6052 18420
rect 6552 18368 6604 18420
rect 10692 18411 10744 18420
rect 10692 18377 10701 18411
rect 10701 18377 10735 18411
rect 10735 18377 10744 18411
rect 10692 18368 10744 18377
rect 11336 18368 11388 18420
rect 11980 18368 12032 18420
rect 15292 18411 15344 18420
rect 15292 18377 15301 18411
rect 15301 18377 15335 18411
rect 15335 18377 15344 18411
rect 15292 18368 15344 18377
rect 15384 18368 15436 18420
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 6368 18232 6420 18284
rect 9312 18232 9364 18284
rect 9680 18275 9732 18284
rect 9680 18241 9689 18275
rect 9689 18241 9723 18275
rect 9723 18241 9732 18275
rect 9680 18232 9732 18241
rect 2044 18207 2096 18216
rect 2044 18173 2078 18207
rect 2078 18173 2096 18207
rect 2044 18164 2096 18173
rect 4344 18164 4396 18216
rect 5632 18164 5684 18216
rect 4620 18096 4672 18148
rect 5080 18096 5132 18148
rect 11060 18232 11112 18284
rect 16120 18232 16172 18284
rect 10876 18164 10928 18216
rect 11244 18164 11296 18216
rect 12164 18164 12216 18216
rect 12532 18164 12584 18216
rect 6644 18096 6696 18148
rect 7196 18139 7248 18148
rect 7196 18105 7205 18139
rect 7205 18105 7239 18139
rect 7239 18105 7248 18139
rect 7196 18096 7248 18105
rect 9404 18096 9456 18148
rect 13544 18096 13596 18148
rect 6736 18028 6788 18080
rect 8208 18028 8260 18080
rect 9220 18071 9272 18080
rect 9220 18037 9229 18071
rect 9229 18037 9263 18071
rect 9263 18037 9272 18071
rect 9220 18028 9272 18037
rect 10692 18028 10744 18080
rect 11520 18028 11572 18080
rect 15292 18164 15344 18216
rect 14372 18071 14424 18080
rect 14372 18037 14381 18071
rect 14381 18037 14415 18071
rect 14415 18037 14424 18071
rect 14372 18028 14424 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1768 17824 1820 17876
rect 2780 17824 2832 17876
rect 4712 17824 4764 17876
rect 5632 17867 5684 17876
rect 5632 17833 5641 17867
rect 5641 17833 5675 17867
rect 5675 17833 5684 17867
rect 5632 17824 5684 17833
rect 11428 17824 11480 17876
rect 13544 17867 13596 17876
rect 13544 17833 13553 17867
rect 13553 17833 13587 17867
rect 13587 17833 13596 17867
rect 13544 17824 13596 17833
rect 14372 17867 14424 17876
rect 14372 17833 14381 17867
rect 14381 17833 14415 17867
rect 14415 17833 14424 17867
rect 14372 17824 14424 17833
rect 3608 17756 3660 17808
rect 4436 17799 4488 17808
rect 4436 17765 4445 17799
rect 4445 17765 4479 17799
rect 4479 17765 4488 17799
rect 4436 17756 4488 17765
rect 2044 17688 2096 17740
rect 6276 17731 6328 17740
rect 4252 17620 4304 17672
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 6276 17697 6310 17731
rect 6310 17697 6328 17731
rect 6276 17688 6328 17697
rect 7380 17688 7432 17740
rect 8024 17688 8076 17740
rect 9956 17731 10008 17740
rect 9956 17697 9990 17731
rect 9990 17697 10008 17731
rect 9956 17688 10008 17697
rect 11060 17688 11112 17740
rect 13544 17688 13596 17740
rect 7932 17663 7984 17672
rect 2964 17552 3016 17604
rect 5632 17552 5684 17604
rect 7932 17629 7941 17663
rect 7941 17629 7975 17663
rect 7975 17629 7984 17663
rect 7932 17620 7984 17629
rect 8576 17663 8628 17672
rect 8576 17629 8585 17663
rect 8585 17629 8619 17663
rect 8619 17629 8628 17663
rect 8576 17620 8628 17629
rect 6368 17484 6420 17536
rect 7380 17527 7432 17536
rect 7380 17493 7389 17527
rect 7389 17493 7423 17527
rect 7423 17493 7432 17527
rect 7380 17484 7432 17493
rect 8300 17527 8352 17536
rect 8300 17493 8309 17527
rect 8309 17493 8343 17527
rect 8343 17493 8352 17527
rect 8300 17484 8352 17493
rect 9036 17527 9088 17536
rect 9036 17493 9045 17527
rect 9045 17493 9079 17527
rect 9079 17493 9088 17527
rect 9036 17484 9088 17493
rect 12164 17663 12216 17672
rect 11152 17484 11204 17536
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2872 17323 2924 17332
rect 2872 17289 2881 17323
rect 2881 17289 2915 17323
rect 2915 17289 2924 17323
rect 2872 17280 2924 17289
rect 4252 17280 4304 17332
rect 4436 17323 4488 17332
rect 4436 17289 4445 17323
rect 4445 17289 4479 17323
rect 4479 17289 4488 17323
rect 4436 17280 4488 17289
rect 5172 17323 5224 17332
rect 5172 17289 5181 17323
rect 5181 17289 5215 17323
rect 5215 17289 5224 17323
rect 5172 17280 5224 17289
rect 6276 17323 6328 17332
rect 6276 17289 6285 17323
rect 6285 17289 6319 17323
rect 6319 17289 6328 17323
rect 6276 17280 6328 17289
rect 6368 17280 6420 17332
rect 9404 17323 9456 17332
rect 2044 17187 2096 17196
rect 2044 17153 2053 17187
rect 2053 17153 2087 17187
rect 2087 17153 2096 17187
rect 2044 17144 2096 17153
rect 3332 17076 3384 17128
rect 3424 17076 3476 17128
rect 4620 17144 4672 17196
rect 6736 17212 6788 17264
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 11336 17280 11388 17332
rect 13544 17323 13596 17332
rect 13544 17289 13553 17323
rect 13553 17289 13587 17323
rect 13587 17289 13596 17323
rect 13544 17280 13596 17289
rect 9312 17187 9364 17196
rect 4712 17076 4764 17128
rect 5540 17119 5592 17128
rect 5540 17085 5549 17119
rect 5549 17085 5583 17119
rect 5583 17085 5592 17119
rect 5540 17076 5592 17085
rect 2320 17008 2372 17060
rect 9312 17153 9321 17187
rect 9321 17153 9355 17187
rect 9355 17153 9364 17187
rect 9312 17144 9364 17153
rect 9772 17144 9824 17196
rect 9036 17076 9088 17128
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 3240 16983 3292 16992
rect 3240 16949 3249 16983
rect 3249 16949 3283 16983
rect 3283 16949 3292 16983
rect 3240 16940 3292 16949
rect 7380 17008 7432 17060
rect 9956 17144 10008 17196
rect 10048 17008 10100 17060
rect 4712 16940 4764 16992
rect 6000 16940 6052 16992
rect 8208 16983 8260 16992
rect 8208 16949 8217 16983
rect 8217 16949 8251 16983
rect 8251 16949 8260 16983
rect 8208 16940 8260 16949
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 11244 17144 11296 17196
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 13452 17144 13504 17196
rect 14372 17187 14424 17196
rect 14372 17153 14381 17187
rect 14381 17153 14415 17187
rect 14415 17153 14424 17187
rect 14372 17144 14424 17153
rect 10692 16940 10744 16992
rect 12532 16983 12584 16992
rect 12532 16949 12541 16983
rect 12541 16949 12575 16983
rect 12575 16949 12584 16983
rect 12532 16940 12584 16949
rect 13176 16940 13228 16992
rect 14188 16983 14240 16992
rect 14188 16949 14197 16983
rect 14197 16949 14231 16983
rect 14231 16949 14240 16983
rect 14188 16940 14240 16949
rect 15752 16983 15804 16992
rect 15752 16949 15761 16983
rect 15761 16949 15795 16983
rect 15795 16949 15804 16983
rect 15752 16940 15804 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2504 16736 2556 16788
rect 3332 16779 3384 16788
rect 3332 16745 3341 16779
rect 3341 16745 3375 16779
rect 3375 16745 3384 16779
rect 3332 16736 3384 16745
rect 3700 16736 3752 16788
rect 4620 16779 4672 16788
rect 4620 16745 4629 16779
rect 4629 16745 4663 16779
rect 4663 16745 4672 16779
rect 4620 16736 4672 16745
rect 5080 16779 5132 16788
rect 5080 16745 5089 16779
rect 5089 16745 5123 16779
rect 5123 16745 5132 16779
rect 5080 16736 5132 16745
rect 5540 16736 5592 16788
rect 6644 16779 6696 16788
rect 6644 16745 6653 16779
rect 6653 16745 6687 16779
rect 6687 16745 6696 16779
rect 6644 16736 6696 16745
rect 6920 16736 6972 16788
rect 8024 16779 8076 16788
rect 8024 16745 8033 16779
rect 8033 16745 8067 16779
rect 8067 16745 8076 16779
rect 8024 16736 8076 16745
rect 8576 16736 8628 16788
rect 9772 16736 9824 16788
rect 2596 16668 2648 16720
rect 2688 16668 2740 16720
rect 2136 16600 2188 16652
rect 2412 16600 2464 16652
rect 3240 16600 3292 16652
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 6828 16600 6880 16652
rect 3424 16532 3476 16584
rect 5080 16532 5132 16584
rect 9036 16668 9088 16720
rect 8576 16600 8628 16652
rect 9220 16600 9272 16652
rect 9680 16668 9732 16720
rect 11428 16736 11480 16788
rect 13820 16736 13872 16788
rect 14832 16736 14884 16788
rect 10784 16668 10836 16720
rect 10968 16600 11020 16652
rect 11060 16600 11112 16652
rect 11612 16643 11664 16652
rect 11612 16609 11621 16643
rect 11621 16609 11655 16643
rect 11655 16609 11664 16643
rect 11612 16600 11664 16609
rect 7288 16575 7340 16584
rect 7288 16541 7297 16575
rect 7297 16541 7331 16575
rect 7331 16541 7340 16575
rect 8484 16575 8536 16584
rect 7288 16532 7340 16541
rect 6552 16464 6604 16516
rect 8484 16541 8493 16575
rect 8493 16541 8527 16575
rect 8527 16541 8536 16575
rect 8484 16532 8536 16541
rect 10692 16575 10744 16584
rect 10692 16541 10701 16575
rect 10701 16541 10735 16575
rect 10735 16541 10744 16575
rect 10692 16532 10744 16541
rect 11704 16532 11756 16584
rect 12164 16532 12216 16584
rect 13452 16668 13504 16720
rect 13636 16668 13688 16720
rect 12532 16575 12584 16584
rect 12532 16541 12541 16575
rect 12541 16541 12575 16575
rect 12575 16541 12584 16575
rect 12532 16532 12584 16541
rect 12624 16575 12676 16584
rect 12624 16541 12633 16575
rect 12633 16541 12667 16575
rect 12667 16541 12676 16575
rect 12624 16532 12676 16541
rect 14188 16575 14240 16584
rect 14188 16541 14197 16575
rect 14197 16541 14231 16575
rect 14231 16541 14240 16575
rect 14188 16532 14240 16541
rect 2044 16396 2096 16448
rect 4988 16439 5040 16448
rect 4988 16405 4997 16439
rect 4997 16405 5031 16439
rect 5031 16405 5040 16439
rect 4988 16396 5040 16405
rect 7748 16439 7800 16448
rect 7748 16405 7757 16439
rect 7757 16405 7791 16439
rect 7791 16405 7800 16439
rect 7748 16396 7800 16405
rect 9128 16439 9180 16448
rect 9128 16405 9137 16439
rect 9137 16405 9171 16439
rect 9171 16405 9180 16439
rect 9128 16396 9180 16405
rect 11060 16396 11112 16448
rect 12256 16396 12308 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 3424 16192 3476 16244
rect 6736 16192 6788 16244
rect 7748 16192 7800 16244
rect 10692 16192 10744 16244
rect 14188 16192 14240 16244
rect 13728 16167 13780 16176
rect 13728 16133 13737 16167
rect 13737 16133 13771 16167
rect 13771 16133 13780 16167
rect 13728 16124 13780 16133
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 5448 16056 5500 16108
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 9404 16099 9456 16108
rect 9404 16065 9413 16099
rect 9413 16065 9447 16099
rect 9447 16065 9456 16099
rect 9404 16056 9456 16065
rect 11152 16056 11204 16108
rect 13636 16056 13688 16108
rect 16764 16056 16816 16108
rect 2136 15988 2188 16040
rect 2688 15988 2740 16040
rect 3148 15988 3200 16040
rect 7196 16031 7248 16040
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 9220 15988 9272 16040
rect 11336 15988 11388 16040
rect 16304 15988 16356 16040
rect 5264 15920 5316 15972
rect 6920 15920 6972 15972
rect 14188 15963 14240 15972
rect 14188 15929 14222 15963
rect 14222 15929 14240 15963
rect 14188 15920 14240 15929
rect 14372 15920 14424 15972
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 1860 15895 1912 15904
rect 1860 15861 1869 15895
rect 1869 15861 1903 15895
rect 1903 15861 1912 15895
rect 1860 15852 1912 15861
rect 2688 15852 2740 15904
rect 3516 15852 3568 15904
rect 5080 15895 5132 15904
rect 5080 15861 5089 15895
rect 5089 15861 5123 15895
rect 5123 15861 5132 15895
rect 5080 15852 5132 15861
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 6552 15852 6604 15861
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 6828 15852 6880 15861
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 8852 15895 8904 15904
rect 8852 15861 8861 15895
rect 8861 15861 8895 15895
rect 8895 15861 8904 15895
rect 8852 15852 8904 15861
rect 9220 15895 9272 15904
rect 9220 15861 9229 15895
rect 9229 15861 9263 15895
rect 9263 15861 9272 15895
rect 9220 15852 9272 15861
rect 10968 15852 11020 15904
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2136 15648 2188 15700
rect 3148 15691 3200 15700
rect 3148 15657 3157 15691
rect 3157 15657 3191 15691
rect 3191 15657 3200 15691
rect 3148 15648 3200 15657
rect 3516 15691 3568 15700
rect 3516 15657 3525 15691
rect 3525 15657 3559 15691
rect 3559 15657 3568 15691
rect 3516 15648 3568 15657
rect 4528 15648 4580 15700
rect 5448 15648 5500 15700
rect 6000 15648 6052 15700
rect 6736 15648 6788 15700
rect 7380 15648 7432 15700
rect 8576 15691 8628 15700
rect 8576 15657 8585 15691
rect 8585 15657 8619 15691
rect 8619 15657 8628 15691
rect 8576 15648 8628 15657
rect 9404 15648 9456 15700
rect 10048 15648 10100 15700
rect 10784 15691 10836 15700
rect 10784 15657 10793 15691
rect 10793 15657 10827 15691
rect 10827 15657 10836 15691
rect 10784 15648 10836 15657
rect 11336 15691 11388 15700
rect 11336 15657 11345 15691
rect 11345 15657 11379 15691
rect 11379 15657 11388 15691
rect 11336 15648 11388 15657
rect 12532 15648 12584 15700
rect 13084 15648 13136 15700
rect 14372 15648 14424 15700
rect 1860 15580 1912 15632
rect 12624 15580 12676 15632
rect 15476 15580 15528 15632
rect 2228 15512 2280 15564
rect 4068 15555 4120 15564
rect 4068 15521 4077 15555
rect 4077 15521 4111 15555
rect 4111 15521 4120 15555
rect 4068 15512 4120 15521
rect 4252 15512 4304 15564
rect 5540 15555 5592 15564
rect 5540 15521 5574 15555
rect 5574 15521 5592 15555
rect 5540 15512 5592 15521
rect 7748 15555 7800 15564
rect 7748 15521 7757 15555
rect 7757 15521 7791 15555
rect 7791 15521 7800 15555
rect 7748 15512 7800 15521
rect 9680 15512 9732 15564
rect 10876 15512 10928 15564
rect 11704 15555 11756 15564
rect 11704 15521 11713 15555
rect 11713 15521 11747 15555
rect 11747 15521 11756 15555
rect 11704 15512 11756 15521
rect 13268 15555 13320 15564
rect 13268 15521 13277 15555
rect 13277 15521 13311 15555
rect 13311 15521 13320 15555
rect 13268 15512 13320 15521
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 2320 15444 2372 15496
rect 2596 15444 2648 15496
rect 3516 15444 3568 15496
rect 5264 15487 5316 15496
rect 5264 15453 5273 15487
rect 5273 15453 5307 15487
rect 5307 15453 5316 15487
rect 5264 15444 5316 15453
rect 7932 15487 7984 15496
rect 7932 15453 7941 15487
rect 7941 15453 7975 15487
rect 7975 15453 7984 15487
rect 7932 15444 7984 15453
rect 9404 15444 9456 15496
rect 10508 15444 10560 15496
rect 11796 15487 11848 15496
rect 11796 15453 11805 15487
rect 11805 15453 11839 15487
rect 11839 15453 11848 15487
rect 11796 15444 11848 15453
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 11888 15444 11940 15453
rect 13360 15444 13412 15496
rect 14188 15376 14240 15428
rect 3424 15308 3476 15360
rect 8116 15308 8168 15360
rect 9220 15351 9272 15360
rect 9220 15317 9229 15351
rect 9229 15317 9263 15351
rect 9263 15317 9272 15351
rect 9220 15308 9272 15317
rect 9772 15308 9824 15360
rect 11060 15308 11112 15360
rect 12256 15308 12308 15360
rect 12900 15351 12952 15360
rect 12900 15317 12909 15351
rect 12909 15317 12943 15351
rect 12943 15317 12952 15351
rect 12900 15308 12952 15317
rect 14280 15351 14332 15360
rect 14280 15317 14289 15351
rect 14289 15317 14323 15351
rect 14323 15317 14332 15351
rect 14280 15308 14332 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 5540 15104 5592 15156
rect 6736 15104 6788 15156
rect 7196 15104 7248 15156
rect 8208 15104 8260 15156
rect 9496 15104 9548 15156
rect 10508 15147 10560 15156
rect 10508 15113 10517 15147
rect 10517 15113 10551 15147
rect 10551 15113 10560 15147
rect 10508 15104 10560 15113
rect 10692 15104 10744 15156
rect 11888 15104 11940 15156
rect 13084 15147 13136 15156
rect 13084 15113 13093 15147
rect 13093 15113 13127 15147
rect 13127 15113 13136 15147
rect 13084 15104 13136 15113
rect 14188 15104 14240 15156
rect 15292 15104 15344 15156
rect 21824 15147 21876 15156
rect 21824 15113 21833 15147
rect 21833 15113 21867 15147
rect 21867 15113 21876 15147
rect 21824 15104 21876 15113
rect 7380 15011 7432 15020
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7380 14968 7432 14977
rect 8116 14968 8168 15020
rect 1492 14943 1544 14952
rect 1492 14909 1501 14943
rect 1501 14909 1535 14943
rect 1535 14909 1544 14943
rect 1492 14900 1544 14909
rect 4068 14900 4120 14952
rect 5264 14900 5316 14952
rect 1952 14832 2004 14884
rect 4988 14832 5040 14884
rect 6276 14832 6328 14884
rect 6736 14832 6788 14884
rect 7748 14832 7800 14884
rect 9128 14943 9180 14952
rect 9128 14909 9137 14943
rect 9137 14909 9171 14943
rect 9171 14909 9180 14943
rect 9128 14900 9180 14909
rect 9404 14875 9456 14884
rect 9404 14841 9438 14875
rect 9438 14841 9456 14875
rect 9404 14832 9456 14841
rect 11796 14832 11848 14884
rect 12348 14832 12400 14884
rect 12624 14832 12676 14884
rect 14280 14900 14332 14952
rect 20996 14900 21048 14952
rect 14372 14832 14424 14884
rect 2044 14764 2096 14816
rect 3056 14764 3108 14816
rect 3424 14807 3476 14816
rect 3424 14773 3433 14807
rect 3433 14773 3467 14807
rect 3467 14773 3476 14807
rect 3424 14764 3476 14773
rect 7472 14764 7524 14816
rect 12072 14764 12124 14816
rect 12532 14807 12584 14816
rect 12532 14773 12541 14807
rect 12541 14773 12575 14807
rect 12575 14773 12584 14807
rect 12532 14764 12584 14773
rect 12808 14764 12860 14816
rect 13268 14764 13320 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1860 14560 1912 14612
rect 3516 14603 3568 14612
rect 3516 14569 3525 14603
rect 3525 14569 3559 14603
rect 3559 14569 3568 14603
rect 3516 14560 3568 14569
rect 4252 14560 4304 14612
rect 7748 14560 7800 14612
rect 8208 14560 8260 14612
rect 8852 14560 8904 14612
rect 10048 14560 10100 14612
rect 11704 14560 11756 14612
rect 12348 14560 12400 14612
rect 12624 14603 12676 14612
rect 12624 14569 12633 14603
rect 12633 14569 12667 14603
rect 12667 14569 12676 14603
rect 12624 14560 12676 14569
rect 13820 14560 13872 14612
rect 14280 14560 14332 14612
rect 14372 14560 14424 14612
rect 2780 14424 2832 14476
rect 3976 14424 4028 14476
rect 5264 14492 5316 14544
rect 6736 14492 6788 14544
rect 8116 14492 8168 14544
rect 9588 14492 9640 14544
rect 10692 14492 10744 14544
rect 12072 14492 12124 14544
rect 6000 14424 6052 14476
rect 9128 14424 9180 14476
rect 10968 14424 11020 14476
rect 12256 14424 12308 14476
rect 12624 14424 12676 14476
rect 13360 14424 13412 14476
rect 1860 14399 1912 14408
rect 1860 14365 1869 14399
rect 1869 14365 1903 14399
rect 1903 14365 1912 14399
rect 1860 14356 1912 14365
rect 1952 14356 2004 14408
rect 3516 14356 3568 14408
rect 8576 14399 8628 14408
rect 8576 14365 8585 14399
rect 8585 14365 8619 14399
rect 8619 14365 8628 14399
rect 8576 14356 8628 14365
rect 4436 14288 4488 14340
rect 6276 14288 6328 14340
rect 6920 14288 6972 14340
rect 2596 14220 2648 14272
rect 3608 14220 3660 14272
rect 4988 14263 5040 14272
rect 4988 14229 4997 14263
rect 4997 14229 5031 14263
rect 5031 14229 5040 14263
rect 4988 14220 5040 14229
rect 7196 14263 7248 14272
rect 7196 14229 7205 14263
rect 7205 14229 7239 14263
rect 7239 14229 7248 14263
rect 7196 14220 7248 14229
rect 7472 14220 7524 14272
rect 9404 14220 9456 14272
rect 9588 14220 9640 14272
rect 11612 14263 11664 14272
rect 11612 14229 11621 14263
rect 11621 14229 11655 14263
rect 11655 14229 11664 14263
rect 11612 14220 11664 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 3516 14016 3568 14068
rect 3976 14059 4028 14068
rect 3976 14025 3985 14059
rect 3985 14025 4019 14059
rect 4019 14025 4028 14059
rect 3976 14016 4028 14025
rect 6828 14059 6880 14068
rect 6828 14025 6837 14059
rect 6837 14025 6871 14059
rect 6871 14025 6880 14059
rect 6828 14016 6880 14025
rect 8576 14016 8628 14068
rect 8760 14016 8812 14068
rect 10692 14016 10744 14068
rect 11336 14059 11388 14068
rect 11336 14025 11345 14059
rect 11345 14025 11379 14059
rect 11379 14025 11388 14059
rect 11336 14016 11388 14025
rect 11612 14016 11664 14068
rect 12072 13948 12124 14000
rect 4896 13880 4948 13932
rect 5448 13880 5500 13932
rect 6000 13880 6052 13932
rect 7196 13880 7248 13932
rect 13360 14016 13412 14068
rect 16396 13923 16448 13932
rect 1492 13812 1544 13864
rect 1768 13812 1820 13864
rect 3056 13812 3108 13864
rect 4160 13787 4212 13796
rect 4160 13753 4169 13787
rect 4169 13753 4203 13787
rect 4203 13753 4212 13787
rect 4160 13744 4212 13753
rect 6920 13812 6972 13864
rect 8392 13855 8444 13864
rect 8392 13821 8401 13855
rect 8401 13821 8435 13855
rect 8435 13821 8444 13855
rect 8392 13812 8444 13821
rect 16396 13889 16405 13923
rect 16405 13889 16439 13923
rect 16439 13889 16448 13923
rect 16396 13880 16448 13889
rect 20996 13923 21048 13932
rect 20996 13889 21005 13923
rect 21005 13889 21039 13923
rect 21039 13889 21048 13923
rect 20996 13880 21048 13889
rect 16120 13855 16172 13864
rect 6460 13744 6512 13796
rect 10876 13787 10928 13796
rect 10876 13753 10885 13787
rect 10885 13753 10919 13787
rect 10919 13753 10928 13787
rect 10876 13744 10928 13753
rect 16120 13821 16129 13855
rect 16129 13821 16163 13855
rect 16163 13821 16172 13855
rect 16120 13812 16172 13821
rect 20720 13855 20772 13864
rect 20720 13821 20729 13855
rect 20729 13821 20763 13855
rect 20763 13821 20772 13855
rect 20720 13812 20772 13821
rect 2320 13676 2372 13728
rect 6000 13676 6052 13728
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 12624 13676 12676 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2780 13515 2832 13524
rect 2780 13481 2789 13515
rect 2789 13481 2823 13515
rect 2823 13481 2832 13515
rect 2780 13472 2832 13481
rect 3056 13515 3108 13524
rect 3056 13481 3065 13515
rect 3065 13481 3099 13515
rect 3099 13481 3108 13515
rect 3056 13472 3108 13481
rect 3884 13472 3936 13524
rect 4068 13472 4120 13524
rect 6368 13472 6420 13524
rect 4712 13404 4764 13456
rect 6092 13404 6144 13456
rect 1676 13336 1728 13388
rect 3608 13379 3660 13388
rect 3608 13345 3617 13379
rect 3617 13345 3651 13379
rect 3651 13345 3660 13379
rect 3608 13336 3660 13345
rect 2136 13311 2188 13320
rect 2136 13277 2145 13311
rect 2145 13277 2179 13311
rect 2179 13277 2188 13311
rect 2136 13268 2188 13277
rect 2320 13311 2372 13320
rect 2320 13277 2329 13311
rect 2329 13277 2363 13311
rect 2363 13277 2372 13311
rect 2320 13268 2372 13277
rect 5172 13268 5224 13320
rect 6000 13268 6052 13320
rect 7196 13472 7248 13524
rect 8208 13472 8260 13524
rect 10140 13515 10192 13524
rect 10140 13481 10149 13515
rect 10149 13481 10183 13515
rect 10183 13481 10192 13515
rect 10140 13472 10192 13481
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12900 13515 12952 13524
rect 12440 13472 12492 13481
rect 12900 13481 12909 13515
rect 12909 13481 12943 13515
rect 12943 13481 12952 13515
rect 12900 13472 12952 13481
rect 6920 13447 6972 13456
rect 6920 13413 6929 13447
rect 6929 13413 6963 13447
rect 6963 13413 6972 13447
rect 6920 13404 6972 13413
rect 8116 13404 8168 13456
rect 9588 13404 9640 13456
rect 10048 13379 10100 13388
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 7932 13268 7984 13320
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 12624 13404 12676 13456
rect 17592 13404 17644 13456
rect 11888 13336 11940 13388
rect 12164 13336 12216 13388
rect 17408 13379 17460 13388
rect 17408 13345 17417 13379
rect 17417 13345 17451 13379
rect 17451 13345 17460 13379
rect 17408 13336 17460 13345
rect 8024 13243 8076 13252
rect 8024 13209 8033 13243
rect 8033 13209 8067 13243
rect 8067 13209 8076 13243
rect 8024 13200 8076 13209
rect 2688 13132 2740 13184
rect 13728 13268 13780 13320
rect 10876 13200 10928 13252
rect 12624 13200 12676 13252
rect 9220 13132 9272 13184
rect 10968 13132 11020 13184
rect 11428 13175 11480 13184
rect 11428 13141 11437 13175
rect 11437 13141 11471 13175
rect 11471 13141 11480 13175
rect 11428 13132 11480 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1676 12971 1728 12980
rect 1676 12937 1685 12971
rect 1685 12937 1719 12971
rect 1719 12937 1728 12971
rect 1676 12928 1728 12937
rect 2136 12971 2188 12980
rect 2136 12937 2145 12971
rect 2145 12937 2179 12971
rect 2179 12937 2188 12971
rect 2136 12928 2188 12937
rect 1768 12860 1820 12912
rect 3884 12928 3936 12980
rect 4804 12971 4856 12980
rect 4804 12937 4813 12971
rect 4813 12937 4847 12971
rect 4847 12937 4856 12971
rect 4804 12928 4856 12937
rect 6368 12928 6420 12980
rect 7932 12971 7984 12980
rect 7932 12937 7941 12971
rect 7941 12937 7975 12971
rect 7975 12937 7984 12971
rect 7932 12928 7984 12937
rect 9680 12928 9732 12980
rect 10140 12928 10192 12980
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 12440 12971 12492 12980
rect 12440 12937 12449 12971
rect 12449 12937 12483 12971
rect 12483 12937 12492 12971
rect 12440 12928 12492 12937
rect 12900 12928 12952 12980
rect 16212 12928 16264 12980
rect 4712 12903 4764 12912
rect 4712 12869 4721 12903
rect 4721 12869 4755 12903
rect 4755 12869 4764 12903
rect 4712 12860 4764 12869
rect 10416 12903 10468 12912
rect 10416 12869 10425 12903
rect 10425 12869 10459 12903
rect 10459 12869 10468 12903
rect 10416 12860 10468 12869
rect 5264 12835 5316 12844
rect 5264 12801 5273 12835
rect 5273 12801 5307 12835
rect 5307 12801 5316 12835
rect 5264 12792 5316 12801
rect 2412 12724 2464 12776
rect 5172 12767 5224 12776
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 5172 12724 5224 12733
rect 4712 12656 4764 12708
rect 7840 12792 7892 12844
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 10968 12835 11020 12844
rect 10968 12801 10977 12835
rect 10977 12801 11011 12835
rect 11011 12801 11020 12835
rect 10968 12792 11020 12801
rect 13084 12792 13136 12844
rect 13728 12860 13780 12912
rect 16764 12860 16816 12912
rect 17408 12860 17460 12912
rect 16948 12835 17000 12844
rect 8300 12767 8352 12776
rect 8300 12733 8309 12767
rect 8309 12733 8343 12767
rect 8343 12733 8352 12767
rect 8300 12724 8352 12733
rect 12164 12767 12216 12776
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 12532 12724 12584 12776
rect 14004 12767 14056 12776
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 18328 12835 18380 12844
rect 18328 12801 18337 12835
rect 18337 12801 18371 12835
rect 18371 12801 18380 12835
rect 18328 12792 18380 12801
rect 14004 12724 14056 12733
rect 16672 12767 16724 12776
rect 16672 12733 16681 12767
rect 16681 12733 16715 12767
rect 16715 12733 16724 12767
rect 16672 12724 16724 12733
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 5540 12656 5592 12708
rect 6000 12656 6052 12708
rect 9220 12656 9272 12708
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 7840 12588 7892 12640
rect 10784 12631 10836 12640
rect 10784 12597 10793 12631
rect 10793 12597 10827 12631
rect 10827 12597 10836 12631
rect 10784 12588 10836 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2412 12384 2464 12436
rect 7472 12427 7524 12436
rect 6552 12359 6604 12368
rect 6552 12325 6561 12359
rect 6561 12325 6595 12359
rect 6595 12325 6604 12359
rect 6552 12316 6604 12325
rect 1952 12248 2004 12300
rect 3884 12248 3936 12300
rect 4712 12248 4764 12300
rect 6000 12248 6052 12300
rect 6920 12316 6972 12368
rect 7472 12393 7481 12427
rect 7481 12393 7515 12427
rect 7515 12393 7524 12427
rect 7472 12384 7524 12393
rect 9220 12427 9272 12436
rect 9220 12393 9229 12427
rect 9229 12393 9263 12427
rect 9263 12393 9272 12427
rect 9220 12384 9272 12393
rect 10784 12384 10836 12436
rect 12532 12384 12584 12436
rect 13084 12427 13136 12436
rect 13084 12393 13093 12427
rect 13093 12393 13127 12427
rect 13127 12393 13136 12427
rect 13084 12384 13136 12393
rect 13268 12427 13320 12436
rect 13268 12393 13277 12427
rect 13277 12393 13311 12427
rect 13311 12393 13320 12427
rect 13268 12384 13320 12393
rect 8484 12316 8536 12368
rect 10968 12316 11020 12368
rect 1676 12180 1728 12232
rect 2412 12223 2464 12232
rect 2412 12189 2421 12223
rect 2421 12189 2455 12223
rect 2455 12189 2464 12223
rect 2412 12180 2464 12189
rect 6552 12180 6604 12232
rect 9036 12248 9088 12300
rect 11428 12248 11480 12300
rect 14372 12248 14424 12300
rect 7840 12223 7892 12232
rect 1768 12155 1820 12164
rect 1768 12121 1777 12155
rect 1777 12121 1811 12155
rect 1811 12121 1820 12155
rect 1768 12112 1820 12121
rect 6276 12112 6328 12164
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 9128 12180 9180 12232
rect 10784 12223 10836 12232
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 11888 12180 11940 12232
rect 12440 12180 12492 12232
rect 13820 12223 13872 12232
rect 13820 12189 13829 12223
rect 13829 12189 13863 12223
rect 13863 12189 13872 12223
rect 13820 12180 13872 12189
rect 3148 12087 3200 12096
rect 3148 12053 3157 12087
rect 3157 12053 3191 12087
rect 3191 12053 3200 12087
rect 3148 12044 3200 12053
rect 5448 12087 5500 12096
rect 5448 12053 5457 12087
rect 5457 12053 5491 12087
rect 5491 12053 5500 12087
rect 5448 12044 5500 12053
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 6920 12087 6972 12096
rect 6920 12053 6929 12087
rect 6929 12053 6963 12087
rect 6963 12053 6972 12087
rect 6920 12044 6972 12053
rect 10140 12044 10192 12096
rect 12164 12087 12216 12096
rect 12164 12053 12173 12087
rect 12173 12053 12207 12087
rect 12207 12053 12216 12087
rect 12164 12044 12216 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2412 11840 2464 11892
rect 3240 11840 3292 11892
rect 5356 11883 5408 11892
rect 2228 11747 2280 11756
rect 2228 11713 2237 11747
rect 2237 11713 2271 11747
rect 2271 11713 2280 11747
rect 2228 11704 2280 11713
rect 5356 11849 5365 11883
rect 5365 11849 5399 11883
rect 5399 11849 5408 11883
rect 5356 11840 5408 11849
rect 6276 11883 6328 11892
rect 6276 11849 6285 11883
rect 6285 11849 6319 11883
rect 6319 11849 6328 11883
rect 6276 11840 6328 11849
rect 7840 11840 7892 11892
rect 10968 11840 11020 11892
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 14372 11883 14424 11892
rect 14372 11849 14381 11883
rect 14381 11849 14415 11883
rect 14415 11849 14424 11883
rect 14372 11840 14424 11849
rect 2320 11636 2372 11688
rect 3148 11636 3200 11688
rect 3884 11679 3936 11688
rect 3884 11645 3893 11679
rect 3893 11645 3927 11679
rect 3927 11645 3936 11679
rect 3884 11636 3936 11645
rect 6920 11636 6972 11688
rect 7840 11636 7892 11688
rect 9128 11636 9180 11688
rect 9588 11679 9640 11688
rect 9588 11645 9622 11679
rect 9622 11645 9640 11679
rect 4988 11568 5040 11620
rect 9588 11636 9640 11645
rect 12348 11636 12400 11688
rect 12532 11636 12584 11688
rect 9680 11568 9732 11620
rect 1676 11543 1728 11552
rect 1676 11509 1685 11543
rect 1685 11509 1719 11543
rect 1719 11509 1728 11543
rect 1676 11500 1728 11509
rect 2136 11543 2188 11552
rect 2136 11509 2145 11543
rect 2145 11509 2179 11543
rect 2179 11509 2188 11543
rect 3056 11543 3108 11552
rect 2136 11500 2188 11509
rect 3056 11509 3065 11543
rect 3065 11509 3099 11543
rect 3099 11509 3108 11543
rect 3056 11500 3108 11509
rect 3608 11500 3660 11552
rect 6552 11543 6604 11552
rect 6552 11509 6561 11543
rect 6561 11509 6595 11543
rect 6595 11509 6604 11543
rect 6552 11500 6604 11509
rect 9036 11500 9088 11552
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2136 11296 2188 11348
rect 4712 11339 4764 11348
rect 4712 11305 4721 11339
rect 4721 11305 4755 11339
rect 4755 11305 4764 11339
rect 4712 11296 4764 11305
rect 6276 11296 6328 11348
rect 6920 11296 6972 11348
rect 7472 11296 7524 11348
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 8944 11339 8996 11348
rect 8944 11305 8953 11339
rect 8953 11305 8987 11339
rect 8987 11305 8996 11339
rect 8944 11296 8996 11305
rect 10784 11296 10836 11348
rect 12348 11296 12400 11348
rect 12532 11339 12584 11348
rect 12532 11305 12541 11339
rect 12541 11305 12575 11339
rect 12575 11305 12584 11339
rect 12532 11296 12584 11305
rect 14096 11339 14148 11348
rect 14096 11305 14105 11339
rect 14105 11305 14139 11339
rect 14139 11305 14148 11339
rect 14096 11296 14148 11305
rect 1676 11228 1728 11280
rect 5448 11228 5500 11280
rect 1860 11160 1912 11212
rect 2504 11160 2556 11212
rect 4528 11160 4580 11212
rect 4988 11203 5040 11212
rect 4988 11169 4997 11203
rect 4997 11169 5031 11203
rect 5031 11169 5040 11203
rect 4988 11160 5040 11169
rect 5540 11160 5592 11212
rect 8484 11160 8536 11212
rect 8760 11160 8812 11212
rect 10968 11160 11020 11212
rect 13728 11228 13780 11280
rect 12808 11160 12860 11212
rect 18512 11203 18564 11212
rect 18512 11169 18521 11203
rect 18521 11169 18555 11203
rect 18555 11169 18564 11203
rect 18512 11160 18564 11169
rect 18788 11203 18840 11212
rect 18788 11169 18797 11203
rect 18797 11169 18831 11203
rect 18831 11169 18840 11203
rect 18788 11160 18840 11169
rect 1768 11092 1820 11144
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 7288 11092 7340 11144
rect 8208 11092 8260 11144
rect 10692 11135 10744 11144
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 2136 11024 2188 11076
rect 3056 11024 3108 11076
rect 7472 11067 7524 11076
rect 7472 11033 7481 11067
rect 7481 11033 7515 11067
rect 7515 11033 7524 11067
rect 7472 11024 7524 11033
rect 8300 11024 8352 11076
rect 8576 11024 8628 11076
rect 10232 11067 10284 11076
rect 10232 11033 10241 11067
rect 10241 11033 10275 11067
rect 10275 11033 10284 11067
rect 10232 11024 10284 11033
rect 2228 10956 2280 11008
rect 2412 10956 2464 11008
rect 10876 10956 10928 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 3240 10795 3292 10804
rect 3240 10761 3249 10795
rect 3249 10761 3283 10795
rect 3283 10761 3292 10795
rect 3240 10752 3292 10761
rect 4160 10795 4212 10804
rect 4160 10761 4169 10795
rect 4169 10761 4203 10795
rect 4203 10761 4212 10795
rect 4160 10752 4212 10761
rect 5448 10795 5500 10804
rect 5448 10761 5457 10795
rect 5457 10761 5491 10795
rect 5491 10761 5500 10795
rect 5448 10752 5500 10761
rect 5540 10752 5592 10804
rect 9036 10795 9088 10804
rect 9036 10761 9045 10795
rect 9045 10761 9079 10795
rect 9079 10761 9088 10795
rect 9036 10752 9088 10761
rect 9772 10752 9824 10804
rect 10048 10752 10100 10804
rect 10692 10752 10744 10804
rect 12440 10795 12492 10804
rect 12440 10761 12449 10795
rect 12449 10761 12483 10795
rect 12483 10761 12492 10795
rect 12440 10752 12492 10761
rect 13728 10752 13780 10804
rect 18512 10795 18564 10804
rect 18512 10761 18521 10795
rect 18521 10761 18555 10795
rect 18555 10761 18564 10795
rect 18512 10752 18564 10761
rect 7564 10616 7616 10668
rect 10876 10616 10928 10668
rect 12532 10616 12584 10668
rect 21364 10616 21416 10668
rect 2412 10548 2464 10600
rect 4160 10548 4212 10600
rect 20168 10591 20220 10600
rect 20168 10557 20177 10591
rect 20177 10557 20211 10591
rect 20211 10557 20220 10591
rect 20168 10548 20220 10557
rect 2136 10523 2188 10532
rect 2136 10489 2170 10523
rect 2170 10489 2188 10523
rect 2136 10480 2188 10489
rect 4528 10480 4580 10532
rect 7288 10480 7340 10532
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 4620 10412 4672 10464
rect 8208 10480 8260 10532
rect 12164 10523 12216 10532
rect 12164 10489 12173 10523
rect 12173 10489 12207 10523
rect 12207 10489 12216 10523
rect 12164 10480 12216 10489
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 11060 10412 11112 10464
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 12716 10412 12768 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 2320 10208 2372 10260
rect 2688 10208 2740 10260
rect 4620 10208 4672 10260
rect 5632 10251 5684 10260
rect 5632 10217 5641 10251
rect 5641 10217 5675 10251
rect 5675 10217 5684 10251
rect 5632 10208 5684 10217
rect 6000 10251 6052 10260
rect 6000 10217 6009 10251
rect 6009 10217 6043 10251
rect 6043 10217 6052 10251
rect 6000 10208 6052 10217
rect 6828 10208 6880 10260
rect 7288 10251 7340 10260
rect 7288 10217 7297 10251
rect 7297 10217 7331 10251
rect 7331 10217 7340 10251
rect 7288 10208 7340 10217
rect 7748 10251 7800 10260
rect 7748 10217 7757 10251
rect 7757 10217 7791 10251
rect 7791 10217 7800 10251
rect 7748 10208 7800 10217
rect 8760 10208 8812 10260
rect 10048 10251 10100 10260
rect 10048 10217 10057 10251
rect 10057 10217 10091 10251
rect 10091 10217 10100 10251
rect 10048 10208 10100 10217
rect 12716 10208 12768 10260
rect 12808 10251 12860 10260
rect 12808 10217 12817 10251
rect 12817 10217 12851 10251
rect 12851 10217 12860 10251
rect 12808 10208 12860 10217
rect 10232 10140 10284 10192
rect 10876 10140 10928 10192
rect 1584 10072 1636 10124
rect 2504 10072 2556 10124
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 4436 10115 4488 10124
rect 4436 10081 4445 10115
rect 4445 10081 4479 10115
rect 4479 10081 4488 10115
rect 4436 10072 4488 10081
rect 7656 10115 7708 10124
rect 7656 10081 7665 10115
rect 7665 10081 7699 10115
rect 7699 10081 7708 10115
rect 7656 10072 7708 10081
rect 18880 10115 18932 10124
rect 18880 10081 18889 10115
rect 18889 10081 18923 10115
rect 18923 10081 18932 10115
rect 18880 10072 18932 10081
rect 19156 10115 19208 10124
rect 19156 10081 19165 10115
rect 19165 10081 19199 10115
rect 19199 10081 19208 10115
rect 19156 10072 19208 10081
rect 2228 10004 2280 10056
rect 4160 10004 4212 10056
rect 4712 10047 4764 10056
rect 4068 9979 4120 9988
rect 4068 9945 4077 9979
rect 4077 9945 4111 9979
rect 4111 9945 4120 9979
rect 4068 9936 4120 9945
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 7932 10004 7984 10056
rect 10140 10047 10192 10056
rect 3884 9911 3936 9920
rect 3884 9877 3893 9911
rect 3893 9877 3927 9911
rect 3927 9877 3936 9911
rect 3884 9868 3936 9877
rect 6828 9911 6880 9920
rect 6828 9877 6837 9911
rect 6837 9877 6871 9911
rect 6871 9877 6880 9911
rect 6828 9868 6880 9877
rect 7564 9868 7616 9920
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 10784 9868 10836 9920
rect 11520 9911 11572 9920
rect 11520 9877 11529 9911
rect 11529 9877 11563 9911
rect 11563 9877 11572 9911
rect 11520 9868 11572 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 4436 9664 4488 9716
rect 6000 9707 6052 9716
rect 6000 9673 6009 9707
rect 6009 9673 6043 9707
rect 6043 9673 6052 9707
rect 6000 9664 6052 9673
rect 6644 9639 6696 9648
rect 6644 9605 6653 9639
rect 6653 9605 6687 9639
rect 6687 9605 6696 9639
rect 7656 9664 7708 9716
rect 10232 9707 10284 9716
rect 10232 9673 10241 9707
rect 10241 9673 10275 9707
rect 10275 9673 10284 9707
rect 10232 9664 10284 9673
rect 18880 9707 18932 9716
rect 18880 9673 18889 9707
rect 18889 9673 18923 9707
rect 18923 9673 18932 9707
rect 18880 9664 18932 9673
rect 9680 9639 9732 9648
rect 6644 9596 6696 9605
rect 9680 9605 9689 9639
rect 9689 9605 9723 9639
rect 9723 9605 9732 9639
rect 9680 9596 9732 9605
rect 10968 9528 11020 9580
rect 20628 9528 20680 9580
rect 2596 9460 2648 9512
rect 4160 9460 4212 9512
rect 5448 9460 5500 9512
rect 6920 9460 6972 9512
rect 7564 9460 7616 9512
rect 7932 9503 7984 9512
rect 7932 9469 7966 9503
rect 7966 9469 7984 9503
rect 7932 9460 7984 9469
rect 19340 9503 19392 9512
rect 19340 9469 19349 9503
rect 19349 9469 19383 9503
rect 19383 9469 19392 9503
rect 19340 9460 19392 9469
rect 2228 9392 2280 9444
rect 3884 9392 3936 9444
rect 5080 9392 5132 9444
rect 7748 9392 7800 9444
rect 2136 9324 2188 9376
rect 5448 9367 5500 9376
rect 5448 9333 5457 9367
rect 5457 9333 5491 9367
rect 5491 9333 5500 9367
rect 5448 9324 5500 9333
rect 8300 9324 8352 9376
rect 10140 9324 10192 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2688 9163 2740 9172
rect 2688 9129 2697 9163
rect 2697 9129 2731 9163
rect 2731 9129 2740 9163
rect 2688 9120 2740 9129
rect 2872 9120 2924 9172
rect 2044 9052 2096 9104
rect 2504 9052 2556 9104
rect 4160 9120 4212 9172
rect 6276 9120 6328 9172
rect 7932 9120 7984 9172
rect 8944 9120 8996 9172
rect 11888 9163 11940 9172
rect 11888 9129 11897 9163
rect 11897 9129 11931 9163
rect 11931 9129 11940 9163
rect 11888 9120 11940 9129
rect 4712 9095 4764 9104
rect 4712 9061 4746 9095
rect 4746 9061 4764 9095
rect 4712 9052 4764 9061
rect 5448 9052 5500 9104
rect 3516 8984 3568 9036
rect 4160 8984 4212 9036
rect 4528 8984 4580 9036
rect 7472 8984 7524 9036
rect 10140 8984 10192 9036
rect 10600 8984 10652 9036
rect 10784 9027 10836 9036
rect 10784 8993 10807 9027
rect 10807 8993 10836 9027
rect 10784 8984 10836 8993
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 2688 8848 2740 8900
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 5540 8780 5592 8832
rect 6736 8823 6788 8832
rect 6736 8789 6745 8823
rect 6745 8789 6779 8823
rect 6779 8789 6788 8823
rect 6736 8780 6788 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1952 8576 2004 8628
rect 2688 8619 2740 8628
rect 2688 8585 2697 8619
rect 2697 8585 2731 8619
rect 2731 8585 2740 8619
rect 2688 8576 2740 8585
rect 2964 8619 3016 8628
rect 2964 8585 2973 8619
rect 2973 8585 3007 8619
rect 3007 8585 3016 8619
rect 2964 8576 3016 8585
rect 4068 8576 4120 8628
rect 4712 8576 4764 8628
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 6736 8576 6788 8628
rect 8300 8619 8352 8628
rect 6828 8551 6880 8560
rect 6828 8517 6837 8551
rect 6837 8517 6871 8551
rect 6871 8517 6880 8551
rect 6828 8508 6880 8517
rect 1584 8440 1636 8492
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 2872 8440 2924 8492
rect 3884 8440 3936 8492
rect 5540 8440 5592 8492
rect 8300 8585 8309 8619
rect 8309 8585 8343 8619
rect 8343 8585 8352 8619
rect 10600 8619 10652 8628
rect 8300 8576 8352 8585
rect 8484 8508 8536 8560
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 10600 8585 10609 8619
rect 10609 8585 10643 8619
rect 10643 8585 10652 8619
rect 10600 8576 10652 8585
rect 10140 8508 10192 8560
rect 8944 8483 8996 8492
rect 8944 8449 8953 8483
rect 8953 8449 8987 8483
rect 8987 8449 8996 8483
rect 8944 8440 8996 8449
rect 2780 8372 2832 8424
rect 2964 8372 3016 8424
rect 4896 8372 4948 8424
rect 4804 8304 4856 8356
rect 6736 8304 6788 8356
rect 1952 8279 2004 8288
rect 1952 8245 1961 8279
rect 1961 8245 1995 8279
rect 1995 8245 2004 8279
rect 1952 8236 2004 8245
rect 8116 8236 8168 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1952 8032 2004 8084
rect 2780 8075 2832 8084
rect 2780 8041 2789 8075
rect 2789 8041 2823 8075
rect 2823 8041 2832 8075
rect 2780 8032 2832 8041
rect 2872 8032 2924 8084
rect 3884 8032 3936 8084
rect 4436 8032 4488 8084
rect 4528 8032 4580 8084
rect 4804 8032 4856 8084
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 7472 8032 7524 8084
rect 8116 8075 8168 8084
rect 8116 8041 8125 8075
rect 8125 8041 8159 8075
rect 8159 8041 8168 8075
rect 8116 8032 8168 8041
rect 8944 8032 8996 8084
rect 2044 8007 2096 8016
rect 2044 7973 2053 8007
rect 2053 7973 2087 8007
rect 2087 7973 2096 8007
rect 2044 7964 2096 7973
rect 6000 7964 6052 8016
rect 5540 7828 5592 7880
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2136 7488 2188 7540
rect 2320 7488 2372 7540
rect 2504 7488 2556 7540
rect 3516 7531 3568 7540
rect 3516 7497 3525 7531
rect 3525 7497 3559 7531
rect 3559 7497 3568 7531
rect 3516 7488 3568 7497
rect 4528 7531 4580 7540
rect 4528 7497 4537 7531
rect 4537 7497 4571 7531
rect 4571 7497 4580 7531
rect 4528 7488 4580 7497
rect 5540 7488 5592 7540
rect 6920 7488 6972 7540
rect 8576 7531 8628 7540
rect 8576 7497 8585 7531
rect 8585 7497 8619 7531
rect 8619 7497 8628 7531
rect 8576 7488 8628 7497
rect 23572 7488 23624 7540
rect 6000 7352 6052 7404
rect 6736 7352 6788 7404
rect 8576 7284 8628 7336
rect 22284 7327 22336 7336
rect 22284 7293 22293 7327
rect 22293 7293 22327 7327
rect 22327 7293 22336 7327
rect 22284 7284 22336 7293
rect 2228 7148 2280 7200
rect 2688 7148 2740 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 22744 6851 22796 6860
rect 22744 6817 22753 6851
rect 22753 6817 22787 6851
rect 22787 6817 22796 6851
rect 22744 6808 22796 6817
rect 23388 6672 23440 6724
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 22744 6443 22796 6452
rect 22744 6409 22753 6443
rect 22753 6409 22787 6443
rect 22787 6409 22796 6443
rect 22744 6400 22796 6409
rect 23848 6443 23900 6452
rect 23848 6409 23857 6443
rect 23857 6409 23891 6443
rect 23891 6409 23900 6443
rect 23848 6400 23900 6409
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 24860 5856 24912 5908
rect 24032 5763 24084 5772
rect 24032 5729 24041 5763
rect 24041 5729 24075 5763
rect 24075 5729 24084 5763
rect 24032 5720 24084 5729
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 24032 5355 24084 5364
rect 24032 5321 24041 5355
rect 24041 5321 24075 5355
rect 24075 5321 24084 5355
rect 24032 5312 24084 5321
rect 24768 5355 24820 5364
rect 24768 5321 24777 5355
rect 24777 5321 24811 5355
rect 24811 5321 24820 5355
rect 24768 5312 24820 5321
rect 24584 5151 24636 5160
rect 24584 5117 24593 5151
rect 24593 5117 24627 5151
rect 24627 5117 24636 5151
rect 24584 5108 24636 5117
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 24768 4811 24820 4820
rect 24768 4777 24777 4811
rect 24777 4777 24811 4811
rect 24811 4777 24820 4811
rect 24768 4768 24820 4777
rect 24676 4632 24728 4684
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 24584 4199 24636 4208
rect 24584 4165 24593 4199
rect 24593 4165 24627 4199
rect 24627 4165 24636 4199
rect 24584 4156 24636 4165
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 2596 2907 2648 2916
rect 2596 2873 2630 2907
rect 2630 2873 2648 2907
rect 2596 2864 2648 2873
rect 2780 2796 2832 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2320 2635 2372 2644
rect 2320 2601 2329 2635
rect 2329 2601 2363 2635
rect 2363 2601 2372 2635
rect 2320 2592 2372 2601
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 3146 27520 3202 28000
rect 3422 27704 3478 27713
rect 3422 27639 3478 27648
rect 308 17105 336 27520
rect 860 22137 888 27520
rect 1412 26874 1440 27520
rect 1964 26874 1992 27520
rect 2516 26874 2544 27520
rect 1412 26846 1532 26874
rect 1400 24608 1452 24614
rect 1400 24550 1452 24556
rect 846 22128 902 22137
rect 846 22063 902 22072
rect 1412 21049 1440 24550
rect 1398 21040 1454 21049
rect 1398 20975 1454 20984
rect 1400 19236 1452 19242
rect 1400 19178 1452 19184
rect 1412 18970 1440 19178
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1504 17785 1532 26846
rect 1872 26846 1992 26874
rect 2148 26846 2544 26874
rect 1676 24744 1728 24750
rect 1872 24698 1900 26846
rect 1952 25424 2004 25430
rect 1952 25366 2004 25372
rect 1676 24686 1728 24692
rect 1582 24304 1638 24313
rect 1582 24239 1584 24248
rect 1636 24239 1638 24248
rect 1584 24210 1636 24216
rect 1596 23866 1624 24210
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1584 23180 1636 23186
rect 1584 23122 1636 23128
rect 1596 22778 1624 23122
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1688 21554 1716 24686
rect 1780 24670 1900 24698
rect 1780 21729 1808 24670
rect 1858 24576 1914 24585
rect 1858 24511 1914 24520
rect 1872 24342 1900 24511
rect 1860 24336 1912 24342
rect 1860 24278 1912 24284
rect 1858 23624 1914 23633
rect 1858 23559 1914 23568
rect 1872 23254 1900 23559
rect 1860 23248 1912 23254
rect 1860 23190 1912 23196
rect 1766 21720 1822 21729
rect 1766 21655 1822 21664
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1766 21312 1822 21321
rect 1766 21247 1822 21256
rect 1780 20398 1808 21247
rect 1964 21078 1992 25366
rect 2044 25356 2096 25362
rect 2044 25298 2096 25304
rect 2056 24614 2084 25298
rect 2044 24608 2096 24614
rect 2044 24550 2096 24556
rect 2056 24177 2084 24550
rect 2042 24168 2098 24177
rect 2042 24103 2098 24112
rect 2042 23760 2098 23769
rect 2042 23695 2044 23704
rect 2096 23695 2098 23704
rect 2044 23666 2096 23672
rect 1952 21072 2004 21078
rect 1952 21014 2004 21020
rect 1768 20392 1820 20398
rect 1768 20334 1820 20340
rect 2148 19394 2176 26846
rect 2320 25356 2372 25362
rect 2320 25298 2372 25304
rect 2332 24886 2360 25298
rect 2780 25220 2832 25226
rect 2780 25162 2832 25168
rect 2320 24880 2372 24886
rect 2320 24822 2372 24828
rect 2228 23520 2280 23526
rect 2228 23462 2280 23468
rect 2240 19990 2268 23462
rect 2332 22098 2360 24822
rect 2504 23588 2556 23594
rect 2504 23530 2556 23536
rect 2412 22976 2464 22982
rect 2410 22944 2412 22953
rect 2464 22944 2466 22953
rect 2410 22879 2466 22888
rect 2424 22574 2452 22879
rect 2516 22642 2544 23530
rect 2792 22817 2820 25162
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2884 23497 2912 25094
rect 2964 24268 3016 24274
rect 2964 24210 3016 24216
rect 2976 23526 3004 24210
rect 3056 24064 3108 24070
rect 3056 24006 3108 24012
rect 2964 23520 3016 23526
rect 2870 23488 2926 23497
rect 2964 23462 3016 23468
rect 2870 23423 2926 23432
rect 2872 22976 2924 22982
rect 2872 22918 2924 22924
rect 2778 22808 2834 22817
rect 2596 22772 2648 22778
rect 2778 22743 2834 22752
rect 2596 22714 2648 22720
rect 2504 22636 2556 22642
rect 2504 22578 2556 22584
rect 2412 22568 2464 22574
rect 2412 22510 2464 22516
rect 2608 22234 2636 22714
rect 2596 22228 2648 22234
rect 2596 22170 2648 22176
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2780 22092 2832 22098
rect 2780 22034 2832 22040
rect 2412 22024 2464 22030
rect 2318 21992 2374 22001
rect 2412 21966 2464 21972
rect 2318 21927 2320 21936
rect 2372 21927 2374 21936
rect 2320 21898 2372 21904
rect 2332 21486 2360 21898
rect 2320 21480 2372 21486
rect 2320 21422 2372 21428
rect 2424 21185 2452 21966
rect 2792 21690 2820 22034
rect 2780 21684 2832 21690
rect 2780 21626 2832 21632
rect 2410 21176 2466 21185
rect 2410 21111 2412 21120
rect 2464 21111 2466 21120
rect 2412 21082 2464 21088
rect 2688 21004 2740 21010
rect 2688 20946 2740 20952
rect 2318 20496 2374 20505
rect 2318 20431 2320 20440
rect 2372 20431 2374 20440
rect 2320 20402 2372 20408
rect 2700 20262 2728 20946
rect 2778 20904 2834 20913
rect 2778 20839 2834 20848
rect 2792 20369 2820 20839
rect 2778 20360 2834 20369
rect 2778 20295 2834 20304
rect 2688 20256 2740 20262
rect 2686 20224 2688 20233
rect 2740 20224 2742 20233
rect 2686 20159 2742 20168
rect 2228 19984 2280 19990
rect 2884 19961 2912 22918
rect 2962 22264 3018 22273
rect 2962 22199 3018 22208
rect 2976 21962 3004 22199
rect 2964 21956 3016 21962
rect 2964 21898 3016 21904
rect 3068 21593 3096 24006
rect 3160 23066 3188 27520
rect 3436 27402 3464 27639
rect 3698 27520 3754 28000
rect 4250 27520 4306 28000
rect 4802 27520 4858 28000
rect 5354 27520 5410 28000
rect 5998 27520 6054 28000
rect 6550 27520 6606 28000
rect 7102 27520 7158 28000
rect 7654 27520 7710 28000
rect 8206 27520 8262 28000
rect 8850 27520 8906 28000
rect 9402 27520 9458 28000
rect 9954 27520 10010 28000
rect 10506 27520 10562 28000
rect 11058 27520 11114 28000
rect 11702 27520 11758 28000
rect 12254 27520 12310 28000
rect 12806 27520 12862 28000
rect 13358 27520 13414 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15106 27520 15162 28000
rect 15658 27520 15714 28000
rect 16210 27520 16266 28000
rect 16762 27520 16818 28000
rect 17406 27520 17462 28000
rect 17958 27520 18014 28000
rect 18510 27520 18566 28000
rect 19062 27520 19118 28000
rect 19614 27520 19670 28000
rect 20258 27520 20314 28000
rect 20810 27520 20866 28000
rect 21362 27520 21418 28000
rect 21914 27520 21970 28000
rect 22466 27520 22522 28000
rect 23110 27520 23166 28000
rect 23662 27520 23718 28000
rect 24214 27520 24270 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 3424 27396 3476 27402
rect 3424 27338 3476 27344
rect 3514 27160 3570 27169
rect 3514 27095 3570 27104
rect 3422 26480 3478 26489
rect 3422 26415 3478 26424
rect 3436 26314 3464 26415
rect 3528 26382 3556 27095
rect 3516 26376 3568 26382
rect 3516 26318 3568 26324
rect 3424 26308 3476 26314
rect 3424 26250 3476 26256
rect 3238 25936 3294 25945
rect 3238 25871 3294 25880
rect 3252 24886 3280 25871
rect 3514 25256 3570 25265
rect 3514 25191 3516 25200
rect 3568 25191 3570 25200
rect 3516 25162 3568 25168
rect 3240 24880 3292 24886
rect 3240 24822 3292 24828
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3436 23866 3464 24550
rect 3424 23860 3476 23866
rect 3424 23802 3476 23808
rect 3424 23180 3476 23186
rect 3424 23122 3476 23128
rect 3160 23038 3372 23066
rect 3240 22976 3292 22982
rect 3240 22918 3292 22924
rect 3252 22642 3280 22918
rect 3240 22636 3292 22642
rect 3240 22578 3292 22584
rect 3146 22536 3202 22545
rect 3146 22471 3148 22480
rect 3200 22471 3202 22480
rect 3148 22442 3200 22448
rect 3252 22234 3280 22578
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3054 21584 3110 21593
rect 3054 21519 3110 21528
rect 3056 21004 3108 21010
rect 3056 20946 3108 20952
rect 3068 20262 3096 20946
rect 3148 20800 3200 20806
rect 3148 20742 3200 20748
rect 3056 20256 3108 20262
rect 3056 20198 3108 20204
rect 2228 19926 2280 19932
rect 2870 19952 2926 19961
rect 2870 19887 2926 19896
rect 2320 19848 2372 19854
rect 2318 19816 2320 19825
rect 2372 19816 2374 19825
rect 2318 19751 2374 19760
rect 2504 19712 2556 19718
rect 2504 19654 2556 19660
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 1688 19366 2176 19394
rect 1490 17776 1546 17785
rect 1490 17711 1546 17720
rect 1688 17513 1716 19366
rect 2516 19174 2544 19654
rect 2596 19372 2648 19378
rect 2596 19314 2648 19320
rect 2044 19168 2096 19174
rect 2044 19110 2096 19116
rect 2504 19168 2556 19174
rect 2504 19110 2556 19116
rect 2056 19009 2084 19110
rect 2042 19000 2098 19009
rect 2042 18935 2098 18944
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 2056 18222 2084 18566
rect 1768 18216 1820 18222
rect 1766 18184 1768 18193
rect 2044 18216 2096 18222
rect 1820 18184 1822 18193
rect 2044 18158 2096 18164
rect 1766 18119 1822 18128
rect 1780 17882 1808 18119
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 2410 17776 2466 17785
rect 2044 17740 2096 17746
rect 2410 17711 2466 17720
rect 2044 17682 2096 17688
rect 1674 17504 1730 17513
rect 1674 17439 1730 17448
rect 294 17096 350 17105
rect 294 17031 350 17040
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 16697 1624 16934
rect 1582 16688 1638 16697
rect 1582 16623 1638 16632
rect 1490 16008 1546 16017
rect 1490 15943 1546 15952
rect 1504 15910 1532 15943
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1492 14952 1544 14958
rect 1492 14894 1544 14900
rect 1504 13870 1532 14894
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1688 13512 1716 17439
rect 2056 17202 2084 17682
rect 2134 17640 2190 17649
rect 2134 17575 2190 17584
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2148 16658 2176 17575
rect 2318 17096 2374 17105
rect 2318 17031 2320 17040
rect 2372 17031 2374 17040
rect 2320 17002 2372 17008
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 2056 16114 2084 16390
rect 2148 16130 2176 16594
rect 2044 16108 2096 16114
rect 2148 16102 2268 16130
rect 2044 16050 2096 16056
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1872 15638 1900 15846
rect 1860 15632 1912 15638
rect 1860 15574 1912 15580
rect 1872 14618 1900 15574
rect 1952 14884 2004 14890
rect 1952 14826 2004 14832
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1964 14414 1992 14826
rect 2056 14822 2084 16050
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 2148 15706 2176 15982
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2240 15570 2268 16102
rect 2228 15564 2280 15570
rect 2228 15506 2280 15512
rect 2332 15502 2360 17002
rect 2424 16658 2452 17711
rect 2516 16794 2544 19110
rect 2608 18630 2636 19314
rect 2964 19236 3016 19242
rect 2964 19178 3016 19184
rect 2976 19145 3004 19178
rect 2962 19136 3018 19145
rect 2962 19071 3018 19080
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 2792 17882 2820 18770
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2884 17338 2912 18702
rect 2976 18630 3004 18702
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2976 17610 3004 18566
rect 2964 17604 3016 17610
rect 2964 17546 3016 17552
rect 3068 17377 3096 19654
rect 3160 18601 3188 20742
rect 3344 19145 3372 23038
rect 3436 21894 3464 23122
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3436 21457 3464 21830
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 3528 21593 3556 21626
rect 3514 21584 3570 21593
rect 3514 21519 3570 21528
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 3712 21162 3740 27520
rect 4264 26874 4292 27520
rect 4264 26846 4384 26874
rect 3790 25256 3846 25265
rect 3790 25191 3846 25200
rect 3804 24750 3832 25191
rect 3884 25152 3936 25158
rect 3884 25094 3936 25100
rect 3896 24818 3924 25094
rect 3884 24812 3936 24818
rect 3884 24754 3936 24760
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 3792 24744 3844 24750
rect 3792 24686 3844 24692
rect 3988 24410 4016 24754
rect 3976 24404 4028 24410
rect 3976 24346 4028 24352
rect 3792 24336 3844 24342
rect 3792 24278 3844 24284
rect 3804 23662 3832 24278
rect 3884 24268 3936 24274
rect 3884 24210 3936 24216
rect 3792 23656 3844 23662
rect 3792 23598 3844 23604
rect 3804 23186 3832 23598
rect 3896 23594 3924 24210
rect 3884 23588 3936 23594
rect 3884 23530 3936 23536
rect 3988 23474 4016 24346
rect 4252 24064 4304 24070
rect 4250 24032 4252 24041
rect 4304 24032 4306 24041
rect 4250 23967 4306 23976
rect 4172 23526 4200 23557
rect 4160 23520 4212 23526
rect 3988 23468 4160 23474
rect 3988 23462 4212 23468
rect 3988 23446 4200 23462
rect 4172 23254 4200 23446
rect 4160 23248 4212 23254
rect 4160 23190 4212 23196
rect 3792 23180 3844 23186
rect 3792 23122 3844 23128
rect 3804 22166 3832 23122
rect 4172 22778 4200 23190
rect 4160 22772 4212 22778
rect 4160 22714 4212 22720
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 3792 22160 3844 22166
rect 3792 22102 3844 22108
rect 3804 21418 3832 22102
rect 4080 21706 4108 22578
rect 4080 21690 4200 21706
rect 4080 21684 4212 21690
rect 4080 21678 4160 21684
rect 3792 21412 3844 21418
rect 3792 21354 3844 21360
rect 3620 21134 3740 21162
rect 3804 21146 3832 21354
rect 3792 21140 3844 21146
rect 3516 20256 3568 20262
rect 3516 20198 3568 20204
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3436 19718 3464 19858
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 3330 19136 3386 19145
rect 3330 19071 3386 19080
rect 3146 18592 3202 18601
rect 3146 18527 3202 18536
rect 3436 17785 3464 19654
rect 3528 18329 3556 20198
rect 3514 18320 3570 18329
rect 3514 18255 3570 18264
rect 3620 17814 3648 21134
rect 3792 21082 3844 21088
rect 3698 21040 3754 21049
rect 3698 20975 3754 20984
rect 3608 17808 3660 17814
rect 3422 17776 3478 17785
rect 3608 17750 3660 17756
rect 3422 17711 3478 17720
rect 3054 17368 3110 17377
rect 2872 17332 2924 17338
rect 3054 17303 3110 17312
rect 2872 17274 2924 17280
rect 3330 17232 3386 17241
rect 3330 17167 3386 17176
rect 3344 17134 3372 17167
rect 3332 17128 3384 17134
rect 2870 17096 2926 17105
rect 3332 17070 3384 17076
rect 3424 17128 3476 17134
rect 3620 17105 3648 17750
rect 3424 17070 3476 17076
rect 3606 17096 3662 17105
rect 2870 17031 2926 17040
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1768 13864 1820 13870
rect 1872 13841 1900 14350
rect 1768 13806 1820 13812
rect 1858 13832 1914 13841
rect 1596 13484 1716 13512
rect 1596 10130 1624 13484
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1688 13161 1716 13330
rect 1674 13152 1730 13161
rect 1674 13087 1730 13096
rect 1688 12986 1716 13087
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1780 12918 1808 13806
rect 1858 13767 1914 13776
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 13326 2360 13670
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2148 13025 2176 13262
rect 2134 13016 2190 13025
rect 2134 12951 2136 12960
rect 2188 12951 2190 12960
rect 2136 12922 2188 12928
rect 1768 12912 1820 12918
rect 1768 12854 1820 12860
rect 2332 12866 2360 13262
rect 2424 13002 2452 16594
rect 2608 15858 2636 16662
rect 2700 16046 2728 16662
rect 2688 16040 2740 16046
rect 2688 15982 2740 15988
rect 2688 15904 2740 15910
rect 2608 15852 2688 15858
rect 2740 15852 2820 15858
rect 2608 15830 2820 15852
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2608 14278 2636 15438
rect 2792 14929 2820 15830
rect 2778 14920 2834 14929
rect 2778 14855 2834 14864
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2424 12974 2544 13002
rect 2332 12838 2452 12866
rect 2424 12782 2452 12838
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2424 12442 2452 12718
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 1952 12300 2004 12306
rect 1952 12242 2004 12248
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1766 12200 1822 12209
rect 1688 11558 1716 12174
rect 1766 12135 1768 12144
rect 1820 12135 1822 12144
rect 1768 12106 1820 12112
rect 1676 11552 1728 11558
rect 1676 11494 1728 11500
rect 1688 11286 1716 11494
rect 1676 11280 1728 11286
rect 1676 11222 1728 11228
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10470 1808 11086
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1780 10305 1808 10406
rect 1766 10296 1822 10305
rect 1872 10266 1900 11154
rect 1766 10231 1822 10240
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1596 8498 1624 8774
rect 1964 8634 1992 12242
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2424 11898 2452 12174
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2148 11354 2176 11494
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2240 11098 2268 11698
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2148 11082 2268 11098
rect 2136 11076 2268 11082
rect 2188 11070 2268 11076
rect 2136 11018 2188 11024
rect 2148 10538 2176 11018
rect 2228 11008 2280 11014
rect 2228 10950 2280 10956
rect 2136 10532 2188 10538
rect 2136 10474 2188 10480
rect 2148 9382 2176 10474
rect 2240 10062 2268 10950
rect 2332 10266 2360 11630
rect 2516 11218 2544 12974
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2424 11014 2452 11086
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2502 10840 2558 10849
rect 2502 10775 2558 10784
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 2424 10010 2452 10542
rect 2516 10130 2544 10775
rect 2608 10305 2636 14214
rect 2792 13530 2820 14418
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2700 12889 2728 13126
rect 2686 12880 2742 12889
rect 2686 12815 2742 12824
rect 2594 10296 2650 10305
rect 2884 10282 2912 17031
rect 3240 16992 3292 16998
rect 3146 16960 3202 16969
rect 3240 16934 3292 16940
rect 3146 16895 3202 16904
rect 3160 16046 3188 16895
rect 3252 16658 3280 16934
rect 3344 16794 3372 17070
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3436 16590 3464 17070
rect 3606 17031 3662 17040
rect 3712 16794 3740 20975
rect 3804 20398 3832 21082
rect 3976 20868 4028 20874
rect 3976 20810 4028 20816
rect 3792 20392 3844 20398
rect 3792 20334 3844 20340
rect 3988 19922 4016 20810
rect 4080 20602 4108 21678
rect 4160 21626 4212 21632
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 4080 20330 4108 20538
rect 4068 20324 4120 20330
rect 4068 20266 4120 20272
rect 4066 20224 4122 20233
rect 4066 20159 4122 20168
rect 3976 19916 4028 19922
rect 3976 19858 4028 19864
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3988 19258 4016 19654
rect 4080 19514 4108 20159
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 4356 19417 4384 26846
rect 4620 25356 4672 25362
rect 4620 25298 4672 25304
rect 4632 24614 4660 25298
rect 4620 24608 4672 24614
rect 4620 24550 4672 24556
rect 4526 23080 4582 23089
rect 4526 23015 4582 23024
rect 4540 22098 4568 23015
rect 4436 22092 4488 22098
rect 4436 22034 4488 22040
rect 4528 22092 4580 22098
rect 4528 22034 4580 22040
rect 4448 20874 4476 22034
rect 4540 21690 4568 22034
rect 4528 21684 4580 21690
rect 4528 21626 4580 21632
rect 4436 20868 4488 20874
rect 4436 20810 4488 20816
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4436 19916 4488 19922
rect 4436 19858 4488 19864
rect 4342 19408 4398 19417
rect 4342 19343 4398 19352
rect 3988 19230 4292 19258
rect 3792 19168 3844 19174
rect 4160 19168 4212 19174
rect 3844 19116 4160 19122
rect 3792 19110 4212 19116
rect 3804 19094 4200 19110
rect 4066 18728 4122 18737
rect 4066 18663 4068 18672
rect 4120 18663 4122 18672
rect 4068 18634 4120 18640
rect 3790 17096 3846 17105
rect 3790 17031 3846 17040
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 3436 16250 3464 16526
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 3160 15706 3188 15982
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3528 15706 3556 15846
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3528 15502 3556 15642
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3424 15360 3476 15366
rect 3424 15302 3476 15308
rect 3436 14822 3464 15302
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3068 13870 3096 14758
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3330 13832 3386 13841
rect 3068 13530 3096 13806
rect 3330 13767 3386 13776
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3160 11694 3188 12038
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 3068 11082 3096 11494
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 3252 10810 3280 11834
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 2700 10266 2912 10282
rect 2594 10231 2650 10240
rect 2688 10260 2912 10266
rect 2740 10254 2912 10260
rect 2688 10202 2740 10208
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2240 9450 2268 9998
rect 2424 9982 2544 10010
rect 2516 9466 2544 9982
rect 2596 9512 2648 9518
rect 2516 9460 2596 9466
rect 2516 9454 2648 9460
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 2516 9438 2636 9454
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1964 8090 1992 8230
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 2056 8022 2084 9046
rect 2148 8498 2176 9318
rect 2240 8974 2268 9386
rect 2516 9110 2544 9438
rect 2700 9178 2728 10066
rect 2884 9178 2912 10254
rect 2962 10024 3018 10033
rect 2962 9959 3018 9968
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2686 9072 2742 9081
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2044 8016 2096 8022
rect 2044 7958 2096 7964
rect 2056 3913 2084 7958
rect 2148 7546 2176 8434
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2240 7206 2268 8910
rect 2516 7546 2544 9046
rect 2686 9007 2742 9016
rect 2700 8906 2728 9007
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2700 8634 2728 8842
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2884 8498 2912 9114
rect 2976 8634 3004 9959
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2792 8090 2820 8366
rect 2884 8090 2912 8434
rect 2976 8430 3004 8570
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2042 3904 2098 3913
rect 2042 3839 2098 3848
rect 2332 3058 2360 7482
rect 2688 7200 2740 7206
rect 2740 7148 2820 7154
rect 2688 7142 2820 7148
rect 2700 7126 2820 7142
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2332 2650 2360 2994
rect 2594 2952 2650 2961
rect 2594 2887 2596 2896
rect 2648 2887 2650 2896
rect 2596 2858 2648 2864
rect 2792 2854 2820 7126
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 3344 377 3372 13767
rect 3436 9081 3464 14758
rect 3528 14618 3556 15438
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3528 14414 3556 14554
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3528 14074 3556 14350
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3620 13394 3648 14214
rect 3608 13388 3660 13394
rect 3608 13330 3660 13336
rect 3620 11558 3648 13330
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3698 11520 3754 11529
rect 3514 11248 3570 11257
rect 3514 11183 3570 11192
rect 3528 10577 3556 11183
rect 3514 10568 3570 10577
rect 3514 10503 3570 10512
rect 3422 9072 3478 9081
rect 3422 9007 3478 9016
rect 3516 9036 3568 9042
rect 3620 9024 3648 11494
rect 3698 11455 3754 11464
rect 3568 8996 3648 9024
rect 3516 8978 3568 8984
rect 3528 7546 3556 8978
rect 3712 8265 3740 11455
rect 3698 8256 3754 8265
rect 3698 8191 3754 8200
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3804 2689 3832 17031
rect 4066 16144 4122 16153
rect 4066 16079 4122 16088
rect 3974 15600 4030 15609
rect 4080 15570 4108 16079
rect 3974 15535 4030 15544
rect 4068 15564 4120 15570
rect 3988 14482 4016 15535
rect 4068 15506 4120 15512
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3988 14074 4016 14418
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4080 13530 4108 14894
rect 4172 13802 4200 19094
rect 4264 18902 4292 19230
rect 4448 19122 4476 19858
rect 4540 19310 4568 20742
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4632 19122 4660 24550
rect 4816 23594 4844 27520
rect 4896 25492 4948 25498
rect 4896 25434 4948 25440
rect 4908 24954 4936 25434
rect 5172 25356 5224 25362
rect 5172 25298 5224 25304
rect 5080 25288 5132 25294
rect 5080 25230 5132 25236
rect 4896 24948 4948 24954
rect 4896 24890 4948 24896
rect 5092 24070 5120 25230
rect 5184 24954 5212 25298
rect 5172 24948 5224 24954
rect 5172 24890 5224 24896
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 5184 24313 5212 24550
rect 5368 24449 5396 27520
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5552 24834 5580 25094
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6012 24857 6040 27520
rect 6564 26874 6592 27520
rect 7116 26874 7144 27520
rect 7196 27396 7248 27402
rect 7196 27338 7248 27344
rect 6472 26846 6592 26874
rect 7024 26846 7144 26874
rect 6276 25424 6328 25430
rect 6276 25366 6328 25372
rect 5460 24818 5580 24834
rect 5448 24812 5580 24818
rect 5500 24806 5580 24812
rect 5998 24848 6054 24857
rect 6288 24818 6316 25366
rect 5998 24783 6054 24792
rect 6276 24812 6328 24818
rect 5448 24754 5500 24760
rect 6276 24754 6328 24760
rect 5354 24440 5410 24449
rect 5354 24375 5410 24384
rect 5170 24304 5226 24313
rect 5460 24274 5488 24754
rect 6000 24336 6052 24342
rect 6000 24278 6052 24284
rect 5170 24239 5226 24248
rect 5448 24268 5500 24274
rect 5448 24210 5500 24216
rect 5080 24064 5132 24070
rect 5080 24006 5132 24012
rect 5092 23662 5120 24006
rect 5080 23656 5132 23662
rect 5080 23598 5132 23604
rect 5460 23594 5488 24210
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 4804 23588 4856 23594
rect 4804 23530 4856 23536
rect 5356 23588 5408 23594
rect 5356 23530 5408 23536
rect 5448 23588 5500 23594
rect 5448 23530 5500 23536
rect 5264 22976 5316 22982
rect 5170 22944 5226 22953
rect 5264 22918 5316 22924
rect 5170 22879 5226 22888
rect 5184 22778 5212 22879
rect 5172 22772 5224 22778
rect 5172 22714 5224 22720
rect 4986 22128 5042 22137
rect 4986 22063 5042 22072
rect 4896 20868 4948 20874
rect 4896 20810 4948 20816
rect 4356 19094 4476 19122
rect 4540 19094 4660 19122
rect 4252 18896 4304 18902
rect 4252 18838 4304 18844
rect 4356 18222 4384 19094
rect 4434 19000 4490 19009
rect 4434 18935 4436 18944
rect 4488 18935 4490 18944
rect 4436 18906 4488 18912
rect 4344 18216 4396 18222
rect 4342 18184 4344 18193
rect 4396 18184 4398 18193
rect 4342 18119 4398 18128
rect 4540 18034 4568 19094
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4632 18154 4660 18702
rect 4620 18148 4672 18154
rect 4620 18090 4672 18096
rect 4356 18006 4568 18034
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4264 17513 4292 17614
rect 4250 17504 4306 17513
rect 4250 17439 4306 17448
rect 4264 17338 4292 17439
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4264 14618 4292 15506
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 3896 12986 3924 13466
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3896 12306 3924 12922
rect 3974 12744 4030 12753
rect 3974 12679 4030 12688
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3882 11792 3938 11801
rect 3882 11727 3938 11736
rect 3896 11694 3924 11727
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9450 3924 9862
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3896 8498 3924 9386
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3896 8090 3924 8434
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3988 3369 4016 12679
rect 4066 12472 4122 12481
rect 4066 12407 4122 12416
rect 4080 10962 4108 12407
rect 4080 10934 4200 10962
rect 4172 10810 4200 10934
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4172 10606 4200 10746
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4160 10056 4212 10062
rect 4066 10024 4122 10033
rect 4160 9998 4212 10004
rect 4066 9959 4068 9968
rect 4120 9959 4122 9968
rect 4068 9930 4120 9936
rect 4172 9874 4200 9998
rect 4080 9846 4200 9874
rect 4080 8634 4108 9846
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4172 9178 4200 9454
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4172 9042 4200 9114
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3974 3360 4030 3369
rect 3974 3295 4030 3304
rect 3790 2680 3846 2689
rect 3790 2615 3846 2624
rect 4356 2145 4384 18006
rect 4526 17912 4582 17921
rect 4724 17882 4752 18906
rect 4802 17912 4858 17921
rect 4526 17847 4582 17856
rect 4712 17876 4764 17882
rect 4436 17808 4488 17814
rect 4436 17750 4488 17756
rect 4448 17338 4476 17750
rect 4436 17332 4488 17338
rect 4436 17274 4488 17280
rect 4434 15872 4490 15881
rect 4434 15807 4490 15816
rect 4448 14346 4476 15807
rect 4540 15706 4568 17847
rect 4802 17847 4858 17856
rect 4712 17818 4764 17824
rect 4712 17672 4764 17678
rect 4816 17649 4844 17847
rect 4712 17614 4764 17620
rect 4802 17640 4858 17649
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4632 16794 4660 17138
rect 4724 17134 4752 17614
rect 4802 17575 4858 17584
rect 4712 17128 4764 17134
rect 4908 17105 4936 20810
rect 5000 18136 5028 22063
rect 5172 22024 5224 22030
rect 5276 22012 5304 22918
rect 5224 21984 5304 22012
rect 5172 21966 5224 21972
rect 5172 21888 5224 21894
rect 5172 21830 5224 21836
rect 5184 21418 5212 21830
rect 5276 21690 5304 21984
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 5276 21486 5304 21626
rect 5264 21480 5316 21486
rect 5264 21422 5316 21428
rect 5172 21412 5224 21418
rect 5172 21354 5224 21360
rect 5184 21321 5212 21354
rect 5170 21312 5226 21321
rect 5170 21247 5226 21256
rect 5264 21072 5316 21078
rect 5264 21014 5316 21020
rect 5172 20936 5224 20942
rect 5172 20878 5224 20884
rect 5184 20602 5212 20878
rect 5172 20596 5224 20602
rect 5172 20538 5224 20544
rect 5184 19990 5212 20538
rect 5276 20534 5304 21014
rect 5264 20528 5316 20534
rect 5264 20470 5316 20476
rect 5172 19984 5224 19990
rect 5172 19926 5224 19932
rect 5184 19514 5212 19926
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5264 18896 5316 18902
rect 5264 18838 5316 18844
rect 5080 18148 5132 18154
rect 5000 18108 5080 18136
rect 4712 17070 4764 17076
rect 4894 17096 4950 17105
rect 4724 16998 4752 17070
rect 4894 17031 4950 17040
rect 4712 16992 4764 16998
rect 5000 16946 5028 18108
rect 5080 18090 5132 18096
rect 5170 17640 5226 17649
rect 5170 17575 5226 17584
rect 5184 17338 5212 17575
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 4712 16934 4764 16940
rect 4816 16918 5028 16946
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4436 14340 4488 14346
rect 4436 14282 4488 14288
rect 4816 14090 4844 16918
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5092 16697 5120 16730
rect 5078 16688 5134 16697
rect 5078 16623 5134 16632
rect 5080 16584 5132 16590
rect 5080 16526 5132 16532
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 5000 14890 5028 16390
rect 5092 15910 5120 16526
rect 5276 15978 5304 18838
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 5092 15473 5120 15846
rect 5276 15502 5304 15914
rect 5264 15496 5316 15502
rect 5078 15464 5134 15473
rect 5264 15438 5316 15444
rect 5078 15399 5134 15408
rect 5276 14958 5304 15438
rect 5368 15065 5396 23530
rect 6012 23526 6040 24278
rect 6000 23520 6052 23526
rect 6000 23462 6052 23468
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5538 22672 5594 22681
rect 5448 22636 5500 22642
rect 5538 22607 5594 22616
rect 5448 22578 5500 22584
rect 5460 22098 5488 22578
rect 5552 22574 5580 22607
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 6012 22438 6040 23462
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 5448 22092 5500 22098
rect 5448 22034 5500 22040
rect 6012 21894 6040 22374
rect 6184 22092 6236 22098
rect 6184 22034 6236 22040
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5446 21720 5502 21729
rect 5622 21712 5918 21732
rect 5502 21678 5580 21706
rect 5446 21655 5502 21664
rect 5552 21434 5580 21678
rect 5552 21406 5672 21434
rect 5540 21344 5592 21350
rect 5644 21321 5672 21406
rect 5540 21286 5592 21292
rect 5630 21312 5686 21321
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5460 20584 5488 20946
rect 5552 20913 5580 21286
rect 5630 21247 5686 21256
rect 6012 20942 6040 21830
rect 6196 21350 6224 22034
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6196 21049 6224 21286
rect 6288 21185 6316 21830
rect 6274 21176 6330 21185
rect 6274 21111 6330 21120
rect 6182 21040 6238 21049
rect 6182 20975 6238 20984
rect 6000 20936 6052 20942
rect 5538 20904 5594 20913
rect 6000 20878 6052 20884
rect 5538 20839 5594 20848
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5998 20632 6054 20641
rect 5540 20596 5592 20602
rect 5460 20556 5540 20584
rect 5998 20567 6000 20576
rect 5540 20538 5592 20544
rect 6052 20567 6054 20576
rect 6000 20538 6052 20544
rect 6472 20534 6500 26846
rect 7024 24834 7052 26846
rect 7104 25356 7156 25362
rect 7104 25298 7156 25304
rect 6932 24806 7052 24834
rect 6828 24744 6880 24750
rect 6828 24686 6880 24692
rect 6552 24676 6604 24682
rect 6552 24618 6604 24624
rect 6564 24410 6592 24618
rect 6840 24585 6868 24686
rect 6826 24576 6882 24585
rect 6826 24511 6882 24520
rect 6552 24404 6604 24410
rect 6552 24346 6604 24352
rect 6932 23089 6960 24806
rect 7010 24712 7066 24721
rect 7010 24647 7066 24656
rect 7024 24614 7052 24647
rect 7012 24608 7064 24614
rect 7012 24550 7064 24556
rect 7116 24070 7144 25298
rect 7208 25226 7236 27338
rect 7668 25498 7696 27520
rect 8116 26308 8168 26314
rect 8116 26250 8168 26256
rect 8128 25498 8156 26250
rect 7656 25492 7708 25498
rect 7656 25434 7708 25440
rect 8116 25492 8168 25498
rect 8116 25434 8168 25440
rect 7196 25220 7248 25226
rect 7196 25162 7248 25168
rect 7932 24744 7984 24750
rect 8220 24698 8248 27520
rect 8864 24970 8892 27520
rect 9220 26376 9272 26382
rect 9220 26318 9272 26324
rect 7932 24686 7984 24692
rect 7288 24268 7340 24274
rect 7288 24210 7340 24216
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 7116 23769 7144 24006
rect 7300 23866 7328 24210
rect 7288 23860 7340 23866
rect 7288 23802 7340 23808
rect 7102 23760 7158 23769
rect 7102 23695 7158 23704
rect 7012 23656 7064 23662
rect 7944 23633 7972 24686
rect 8128 24670 8248 24698
rect 8772 24942 8892 24970
rect 8128 24410 8156 24670
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 8116 24404 8168 24410
rect 8116 24346 8168 24352
rect 8024 24268 8076 24274
rect 8024 24210 8076 24216
rect 7012 23598 7064 23604
rect 7930 23624 7986 23633
rect 7024 23322 7052 23598
rect 8036 23610 8064 24210
rect 8128 23866 8156 24346
rect 8220 24206 8248 24550
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 8116 23860 8168 23866
rect 8116 23802 8168 23808
rect 8114 23624 8170 23633
rect 8036 23582 8114 23610
rect 7930 23559 7986 23568
rect 8220 23594 8248 24142
rect 8114 23559 8170 23568
rect 8208 23588 8260 23594
rect 8208 23530 8260 23536
rect 7930 23488 7986 23497
rect 7930 23423 7986 23432
rect 7012 23316 7064 23322
rect 7012 23258 7064 23264
rect 6918 23080 6974 23089
rect 6918 23015 6974 23024
rect 7024 22642 7052 23258
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 6828 22500 6880 22506
rect 6828 22442 6880 22448
rect 6840 22386 6868 22442
rect 7024 22438 7052 22578
rect 7392 22438 7420 23122
rect 7012 22432 7064 22438
rect 6840 22358 6960 22386
rect 7012 22374 7064 22380
rect 7380 22432 7432 22438
rect 7380 22374 7432 22380
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 6748 21622 6776 21966
rect 6932 21962 6960 22358
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 6920 21956 6972 21962
rect 6920 21898 6972 21904
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 6550 21312 6606 21321
rect 6550 21247 6606 21256
rect 6460 20528 6512 20534
rect 6460 20470 6512 20476
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5460 19514 5488 19858
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5538 19408 5594 19417
rect 6196 19394 6224 19654
rect 6104 19378 6224 19394
rect 5538 19343 5594 19352
rect 6092 19372 6224 19378
rect 5552 18970 5580 19343
rect 6144 19366 6224 19372
rect 6092 19314 6144 19320
rect 5998 19136 6054 19145
rect 5998 19071 6054 19080
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 6012 18902 6040 19071
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 6000 18896 6052 18902
rect 6000 18838 6052 18844
rect 5552 18698 5672 18714
rect 5552 18692 5684 18698
rect 5552 18686 5632 18692
rect 5552 17134 5580 18686
rect 5632 18634 5684 18640
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6012 18426 6040 18838
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 5632 18216 5684 18222
rect 5632 18158 5684 18164
rect 5644 17882 5672 18158
rect 5632 17876 5684 17882
rect 5632 17818 5684 17824
rect 5644 17610 5672 17818
rect 5632 17604 5684 17610
rect 5632 17546 5684 17552
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5552 16794 5580 17070
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5460 16114 5488 16594
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5460 15706 5488 16050
rect 6012 15706 6040 16934
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5552 15162 5580 15506
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5354 15056 5410 15065
rect 5354 14991 5410 15000
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 5276 14550 5304 14894
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 4816 14062 4936 14090
rect 4802 13968 4858 13977
rect 4908 13938 4936 14062
rect 4802 13903 4858 13912
rect 4896 13932 4948 13938
rect 4712 13456 4764 13462
rect 4712 13398 4764 13404
rect 4724 12918 4752 13398
rect 4816 12986 4844 13903
rect 4896 13874 4948 13880
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4712 12912 4764 12918
rect 4764 12860 4844 12866
rect 4712 12854 4844 12860
rect 4724 12838 4844 12854
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4724 12306 4752 12650
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4724 11354 4752 12242
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4540 10538 4568 11154
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4632 10266 4660 10406
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4448 9722 4476 10066
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4448 8090 4476 9658
rect 4724 9110 4752 9998
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4540 8090 4568 8978
rect 4724 8634 4752 9046
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4816 8362 4844 12838
rect 5000 11626 5028 14214
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6012 13938 6040 14418
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5184 12782 5212 13262
rect 5460 12889 5488 13874
rect 6012 13734 6040 13874
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13326 6040 13670
rect 6104 13462 6132 18906
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5262 12880 5318 12889
rect 5262 12815 5264 12824
rect 5316 12815 5318 12824
rect 5446 12880 5502 12889
rect 5446 12815 5502 12824
rect 5264 12786 5316 12792
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 6012 12714 6040 13262
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5552 12594 5580 12650
rect 5368 12566 5580 12594
rect 5368 11898 5396 12566
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6012 12102 6040 12242
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 5000 11218 5028 11562
rect 5460 11286 5488 12038
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11801 6040 12038
rect 5998 11792 6054 11801
rect 5998 11727 6054 11736
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 5460 10810 5488 11222
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5552 10810 5580 11154
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5552 9738 5580 10746
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5644 10169 5672 10202
rect 5630 10160 5686 10169
rect 5630 10095 5686 10104
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5460 9710 5580 9738
rect 6012 9722 6040 10202
rect 6000 9716 6052 9722
rect 5460 9518 5488 9710
rect 6000 9658 6052 9664
rect 5448 9512 5500 9518
rect 4894 9480 4950 9489
rect 4894 9415 4950 9424
rect 5078 9480 5134 9489
rect 5448 9454 5500 9460
rect 5078 9415 5080 9424
rect 4908 8634 4936 9415
rect 5132 9415 5134 9424
rect 5080 9386 5132 9392
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5460 9110 5488 9318
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4908 8430 4936 8570
rect 5552 8498 5580 8774
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4816 8090 4844 8298
rect 5552 8090 5580 8434
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 4540 7546 4568 8026
rect 6000 8016 6052 8022
rect 6000 7958 6052 7964
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5552 7546 5580 7822
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 6012 7410 6040 7958
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 4618 4040 4674 4049
rect 4618 3975 4674 3984
rect 4342 2136 4398 2145
rect 4342 2071 4398 2080
rect 4632 480 4660 3975
rect 6196 3505 6224 19366
rect 6274 19272 6330 19281
rect 6274 19207 6276 19216
rect 6328 19207 6330 19216
rect 6276 19178 6328 19184
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6380 18290 6408 18702
rect 6564 18578 6592 21247
rect 6748 21146 6776 21558
rect 7024 21418 7052 21966
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 7576 21486 7604 21830
rect 7944 21554 7972 23423
rect 8220 23322 8248 23530
rect 8208 23316 8260 23322
rect 8208 23258 8260 23264
rect 8024 22568 8076 22574
rect 8024 22510 8076 22516
rect 8036 22030 8064 22510
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 7932 21548 7984 21554
rect 7932 21490 7984 21496
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 7024 21010 7052 21354
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6748 20398 6776 20878
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6840 20074 6868 20946
rect 7024 20602 7052 20946
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 7104 20324 7156 20330
rect 7104 20266 7156 20272
rect 6840 20046 6960 20074
rect 7116 20058 7144 20266
rect 6932 19718 6960 20046
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7012 19916 7064 19922
rect 7012 19858 7064 19864
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6828 19168 6880 19174
rect 7024 19145 7052 19858
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 6828 19110 6880 19116
rect 7010 19136 7066 19145
rect 6656 18873 6684 19110
rect 6642 18864 6698 18873
rect 6642 18799 6698 18808
rect 6472 18550 6684 18578
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6380 17762 6408 18226
rect 6288 17746 6408 17762
rect 6276 17740 6408 17746
rect 6328 17734 6408 17740
rect 6276 17682 6328 17688
rect 6288 17338 6316 17682
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6380 17338 6408 17478
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6276 14884 6328 14890
rect 6276 14826 6328 14832
rect 6288 14346 6316 14826
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 6472 13802 6500 18550
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6564 16674 6592 18362
rect 6656 18154 6684 18550
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6642 17504 6698 17513
rect 6642 17439 6698 17448
rect 6656 16794 6684 17439
rect 6748 17270 6776 18022
rect 6736 17264 6788 17270
rect 6736 17206 6788 17212
rect 6840 16810 6868 19110
rect 7010 19071 7066 19080
rect 6918 18864 6974 18873
rect 7024 18850 7052 19071
rect 6974 18822 7052 18850
rect 6918 18799 6974 18808
rect 7286 18728 7342 18737
rect 7286 18663 7288 18672
rect 7340 18663 7342 18672
rect 7288 18634 7340 18640
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7208 18154 7236 18566
rect 7196 18148 7248 18154
rect 7196 18090 7248 18096
rect 7392 17746 7420 19654
rect 7576 19258 7604 21422
rect 8036 21146 8064 21966
rect 8220 21706 8248 22102
rect 8772 22098 8800 24942
rect 8850 24848 8906 24857
rect 8850 24783 8852 24792
rect 8904 24783 8906 24792
rect 8852 24754 8904 24760
rect 9232 24614 9260 26318
rect 9220 24608 9272 24614
rect 9220 24550 9272 24556
rect 9416 23497 9444 27520
rect 9772 25356 9824 25362
rect 9772 25298 9824 25304
rect 9784 24614 9812 25298
rect 9772 24608 9824 24614
rect 9772 24550 9824 24556
rect 9784 24449 9812 24550
rect 9770 24440 9826 24449
rect 9770 24375 9826 24384
rect 9968 24177 9996 27520
rect 10520 26874 10548 27520
rect 10152 26846 10548 26874
rect 10152 24290 10180 26846
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10876 25288 10928 25294
rect 10876 25230 10928 25236
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10704 24410 10732 24550
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 10060 24262 10180 24290
rect 9954 24168 10010 24177
rect 9954 24103 10010 24112
rect 9680 23520 9732 23526
rect 9402 23488 9458 23497
rect 9680 23462 9732 23468
rect 9402 23423 9458 23432
rect 9588 23248 9640 23254
rect 9588 23190 9640 23196
rect 9600 22778 9628 23190
rect 9588 22772 9640 22778
rect 9588 22714 9640 22720
rect 8760 22092 8812 22098
rect 8760 22034 8812 22040
rect 8220 21678 8340 21706
rect 8772 21690 8800 22034
rect 9494 21992 9550 22001
rect 9494 21927 9550 21936
rect 9508 21690 9536 21927
rect 8312 21622 8340 21678
rect 8760 21684 8812 21690
rect 8760 21626 8812 21632
rect 9496 21684 9548 21690
rect 9496 21626 9548 21632
rect 8300 21616 8352 21622
rect 8300 21558 8352 21564
rect 8852 21616 8904 21622
rect 8852 21558 8904 21564
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 8220 20806 8248 21490
rect 8864 21049 8892 21558
rect 8850 21040 8906 21049
rect 8850 20975 8906 20984
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 8220 20330 8248 20742
rect 9034 20632 9090 20641
rect 9034 20567 9036 20576
rect 9088 20567 9090 20576
rect 9036 20538 9088 20544
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 8208 20324 8260 20330
rect 8208 20266 8260 20272
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8390 19952 8446 19961
rect 8390 19887 8392 19896
rect 8444 19887 8446 19896
rect 8392 19858 8444 19864
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 8022 19816 8078 19825
rect 7944 19378 7972 19790
rect 8022 19751 8024 19760
rect 8076 19751 8078 19760
rect 8024 19722 8076 19728
rect 8404 19394 8432 19858
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 8220 19366 8432 19394
rect 7484 19230 7604 19258
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 17066 7420 17478
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7392 16946 7420 17002
rect 7300 16918 7420 16946
rect 6748 16794 6960 16810
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6748 16788 6972 16794
rect 6748 16782 6920 16788
rect 6564 16646 6684 16674
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 6564 15910 6592 16458
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6564 14385 6592 15846
rect 6550 14376 6606 14385
rect 6550 14311 6606 14320
rect 6460 13796 6512 13802
rect 6460 13738 6512 13744
rect 6472 13705 6500 13738
rect 6458 13696 6514 13705
rect 6458 13631 6514 13640
rect 6368 13524 6420 13530
rect 6656 13512 6684 16646
rect 6748 16250 6776 16782
rect 6920 16730 6972 16736
rect 7194 16688 7250 16697
rect 6828 16652 6880 16658
rect 7194 16623 7250 16632
rect 6828 16594 6880 16600
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6840 16130 6868 16594
rect 6840 16102 6960 16130
rect 6932 15978 6960 16102
rect 7208 16046 7236 16623
rect 7300 16590 7328 16918
rect 7484 16697 7512 19230
rect 8220 19174 8248 19366
rect 8680 19310 8708 19790
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8680 18902 8708 19246
rect 8772 18970 8800 19994
rect 9048 19990 9076 20334
rect 9036 19984 9088 19990
rect 9036 19926 9088 19932
rect 9324 19514 9352 20742
rect 9692 20505 9720 23462
rect 9864 22500 9916 22506
rect 9864 22442 9916 22448
rect 9876 22234 9904 22442
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9864 22228 9916 22234
rect 9864 22170 9916 22176
rect 9678 20496 9734 20505
rect 9678 20431 9734 20440
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9600 20058 9628 20198
rect 9588 20052 9640 20058
rect 9588 19994 9640 20000
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 8850 19136 8906 19145
rect 8850 19071 8906 19080
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 7656 18828 7708 18834
rect 7656 18770 7708 18776
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 7668 17513 7696 18770
rect 7944 17678 7972 18770
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8220 18086 8248 18702
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 7932 17672 7984 17678
rect 7930 17640 7932 17649
rect 7984 17640 7986 17649
rect 7930 17575 7986 17584
rect 7654 17504 7710 17513
rect 7654 17439 7710 17448
rect 8036 16794 8064 17682
rect 8220 16998 8248 18022
rect 8482 17776 8538 17785
rect 8482 17711 8538 17720
rect 8300 17536 8352 17542
rect 8298 17504 8300 17513
rect 8352 17504 8354 17513
rect 8298 17439 8354 17448
rect 8208 16992 8260 16998
rect 8206 16960 8208 16969
rect 8260 16960 8262 16969
rect 8206 16895 8262 16904
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 7470 16688 7526 16697
rect 7470 16623 7526 16632
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6748 15162 6776 15642
rect 6840 15473 6868 15846
rect 6826 15464 6882 15473
rect 6826 15399 6882 15408
rect 6932 15314 6960 15914
rect 6840 15286 6960 15314
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6734 14920 6790 14929
rect 6734 14855 6736 14864
rect 6788 14855 6790 14864
rect 6736 14826 6788 14832
rect 6748 14550 6776 14826
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 6840 14074 6868 15286
rect 7208 15162 7236 15982
rect 7392 15706 7420 16050
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7378 15056 7434 15065
rect 7378 14991 7380 15000
rect 7432 14991 7434 15000
rect 7380 14962 7432 14968
rect 7484 14822 7512 16623
rect 8496 16590 8524 17711
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8588 16794 8616 17614
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8576 16652 8628 16658
rect 8864 16640 8892 19071
rect 9876 18850 9904 22170
rect 9968 21554 9996 22374
rect 10060 21593 10088 24262
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 10152 23186 10180 24142
rect 10704 23730 10732 24346
rect 10692 23724 10744 23730
rect 10692 23666 10744 23672
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 10690 23624 10746 23633
rect 10690 23559 10746 23568
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23180 10192 23186
rect 10140 23122 10192 23128
rect 10152 22098 10180 23122
rect 10704 23066 10732 23559
rect 10796 23254 10824 23666
rect 10888 23662 10916 25230
rect 10876 23656 10928 23662
rect 10876 23598 10928 23604
rect 10874 23488 10930 23497
rect 10874 23423 10930 23432
rect 10784 23248 10836 23254
rect 10784 23190 10836 23196
rect 10704 23038 10824 23066
rect 10692 22976 10744 22982
rect 10692 22918 10744 22924
rect 10704 22642 10732 22918
rect 10692 22636 10744 22642
rect 10692 22578 10744 22584
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10704 22166 10732 22578
rect 10692 22160 10744 22166
rect 10692 22102 10744 22108
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 10046 21584 10102 21593
rect 9956 21548 10008 21554
rect 10152 21554 10180 21830
rect 10704 21690 10732 22102
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10046 21519 10102 21528
rect 10140 21548 10192 21554
rect 9956 21490 10008 21496
rect 10140 21490 10192 21496
rect 10152 21078 10180 21490
rect 10692 21412 10744 21418
rect 10692 21354 10744 21360
rect 10704 21321 10732 21354
rect 10690 21312 10746 21321
rect 10289 21244 10585 21264
rect 10690 21247 10746 21256
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10140 21072 10192 21078
rect 10140 21014 10192 21020
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9968 19990 9996 20402
rect 9956 19984 10008 19990
rect 9956 19926 10008 19932
rect 9968 19514 9996 19926
rect 10060 19922 10088 20878
rect 10152 20602 10180 21014
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 10140 19168 10192 19174
rect 10138 19136 10140 19145
rect 10192 19136 10194 19145
rect 10138 19071 10194 19080
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 9784 18822 9904 18850
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9324 18290 9352 18566
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9404 18148 9456 18154
rect 9404 18090 9456 18096
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9036 17536 9088 17542
rect 9036 17478 9088 17484
rect 9048 17134 9076 17478
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 9048 16726 9076 17070
rect 9036 16720 9088 16726
rect 9036 16662 9088 16668
rect 9232 16658 9260 18022
rect 9416 17338 9444 18090
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9324 17105 9352 17138
rect 9310 17096 9366 17105
rect 9310 17031 9366 17040
rect 9692 16726 9720 18226
rect 9784 17202 9812 18822
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9784 16794 9812 16934
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 8576 16594 8628 16600
rect 8772 16612 8892 16640
rect 9220 16652 9272 16658
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7760 16250 7788 16390
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 8300 15904 8352 15910
rect 8220 15864 8300 15892
rect 7930 15600 7986 15609
rect 7748 15564 7800 15570
rect 7930 15535 7986 15544
rect 7748 15506 7800 15512
rect 7760 14890 7788 15506
rect 7944 15502 7972 15535
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8128 15026 8156 15302
rect 8220 15162 8248 15864
rect 8300 15846 8352 15852
rect 8588 15706 8616 16594
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 7748 14884 7800 14890
rect 7748 14826 7800 14832
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6932 13870 6960 14282
rect 7484 14278 7512 14758
rect 7760 14618 7788 14826
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7208 13938 7236 14214
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 6920 13864 6972 13870
rect 7484 13841 7512 14214
rect 6920 13806 6972 13812
rect 7470 13832 7526 13841
rect 6420 13484 6684 13512
rect 6368 13466 6420 13472
rect 6380 12986 6408 13466
rect 6656 13433 6684 13484
rect 6932 13462 6960 13806
rect 7470 13767 7526 13776
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7208 13530 7236 13670
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 8128 13462 8156 14486
rect 8220 13530 8248 14554
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8588 14249 8616 14350
rect 8574 14240 8630 14249
rect 8574 14175 8630 14184
rect 8588 14074 8616 14175
rect 8772 14074 8800 16612
rect 9220 16594 9272 16600
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8864 14618 8892 15846
rect 9140 15450 9168 16390
rect 9876 16153 9904 18702
rect 10704 18426 10732 20266
rect 10796 20210 10824 23038
rect 10888 22574 10916 23423
rect 10876 22568 10928 22574
rect 10876 22510 10928 22516
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10980 22098 11008 22510
rect 10968 22092 11020 22098
rect 10968 22034 11020 22040
rect 11072 20890 11100 27520
rect 11612 25152 11664 25158
rect 11612 25094 11664 25100
rect 11624 24954 11652 25094
rect 11612 24948 11664 24954
rect 11612 24890 11664 24896
rect 11336 24812 11388 24818
rect 11336 24754 11388 24760
rect 11348 24274 11376 24754
rect 11624 24614 11652 24890
rect 11612 24608 11664 24614
rect 11612 24550 11664 24556
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11348 23526 11376 24210
rect 11520 24064 11572 24070
rect 11520 24006 11572 24012
rect 11532 23730 11560 24006
rect 11520 23724 11572 23730
rect 11520 23666 11572 23672
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 11624 23304 11652 24550
rect 11716 23497 11744 27520
rect 12268 24682 12296 27520
rect 12820 25514 12848 27520
rect 12820 25486 12940 25514
rect 12912 24818 12940 25486
rect 12992 24880 13044 24886
rect 12992 24822 13044 24828
rect 13082 24848 13138 24857
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 12440 24744 12492 24750
rect 12440 24686 12492 24692
rect 12256 24676 12308 24682
rect 12256 24618 12308 24624
rect 12348 24132 12400 24138
rect 12348 24074 12400 24080
rect 11702 23488 11758 23497
rect 11702 23423 11758 23432
rect 11624 23276 11744 23304
rect 11244 21548 11296 21554
rect 11244 21490 11296 21496
rect 11256 21457 11284 21490
rect 11242 21448 11298 21457
rect 11242 21383 11298 21392
rect 10980 20862 11100 20890
rect 10980 20618 11008 20862
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10888 20590 11008 20618
rect 10888 20398 10916 20590
rect 11072 20482 11100 20742
rect 10980 20466 11100 20482
rect 10968 20460 11100 20466
rect 11020 20454 11100 20460
rect 11152 20460 11204 20466
rect 10968 20402 11020 20408
rect 11152 20402 11204 20408
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 10796 20182 11008 20210
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10704 18086 10732 18362
rect 10888 18222 10916 18566
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9968 17202 9996 17682
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 9862 16144 9918 16153
rect 9404 16108 9456 16114
rect 9862 16079 9918 16088
rect 9404 16050 9456 16056
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9232 15910 9260 15982
rect 9220 15904 9272 15910
rect 9272 15864 9352 15892
rect 9220 15846 9272 15852
rect 9140 15422 9260 15450
rect 9232 15366 9260 15422
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9128 14952 9180 14958
rect 8942 14920 8998 14929
rect 9232 14929 9260 15302
rect 9128 14894 9180 14900
rect 9218 14920 9274 14929
rect 8942 14855 8998 14864
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 6920 13456 6972 13462
rect 6642 13424 6698 13433
rect 6920 13398 6972 13404
rect 8116 13456 8168 13462
rect 8116 13398 8168 13404
rect 6642 13359 6698 13368
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 8022 13288 8078 13297
rect 7944 12986 7972 13262
rect 8022 13223 8024 13232
rect 8076 13223 8078 13232
rect 8024 13194 8076 13200
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7470 12880 7526 12889
rect 7470 12815 7526 12824
rect 7840 12844 7892 12850
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6552 12368 6604 12374
rect 6550 12336 6552 12345
rect 6604 12336 6606 12345
rect 6550 12271 6606 12280
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6288 11898 6316 12106
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6564 11558 6592 12174
rect 6552 11552 6604 11558
rect 6550 11520 6552 11529
rect 6604 11520 6606 11529
rect 6550 11455 6606 11464
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6288 10062 6316 11290
rect 6840 10266 6868 12582
rect 7484 12442 7512 12815
rect 7840 12786 7892 12792
rect 7852 12646 7880 12786
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 6920 12368 6972 12374
rect 6972 12328 7052 12356
rect 6920 12310 6972 12316
rect 6920 12096 6972 12102
rect 7024 12073 7052 12328
rect 6920 12038 6972 12044
rect 7010 12064 7066 12073
rect 6932 11694 6960 12038
rect 7010 11999 7066 12008
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6932 11354 6960 11630
rect 7484 11354 7512 12378
rect 7852 12238 7880 12582
rect 8312 12345 8340 12718
rect 8298 12336 8354 12345
rect 8298 12271 8354 12280
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7852 11898 7880 12174
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7852 11694 7880 11834
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 7300 10538 7328 11086
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7484 10713 7512 11018
rect 7470 10704 7526 10713
rect 7470 10639 7526 10648
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7288 10532 7340 10538
rect 7288 10474 7340 10480
rect 7300 10266 7328 10474
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6288 9178 6316 9998
rect 7576 9926 7604 10610
rect 8220 10538 8248 11086
rect 8312 11082 8340 12271
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8220 10418 8248 10474
rect 8220 10390 8340 10418
rect 7746 10296 7802 10305
rect 7746 10231 7748 10240
rect 7800 10231 7802 10240
rect 7748 10202 7800 10208
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 6828 9920 6880 9926
rect 6826 9888 6828 9897
rect 7564 9920 7616 9926
rect 6880 9888 6882 9897
rect 7564 9862 7616 9868
rect 6826 9823 6882 9832
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6656 9081 6684 9590
rect 7576 9518 7604 9862
rect 7668 9722 7696 10066
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 6642 9072 6698 9081
rect 6642 9007 6698 9016
rect 6932 8974 6960 9454
rect 7760 9450 7788 10202
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7944 9518 7972 9998
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7944 9178 7972 9454
rect 8312 9382 8340 10390
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6748 8634 6776 8774
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6840 8401 6868 8502
rect 6826 8392 6882 8401
rect 6736 8356 6788 8362
rect 6826 8327 6882 8336
rect 6736 8298 6788 8304
rect 6748 7410 6776 8298
rect 6932 7546 6960 8910
rect 7484 8498 7512 8978
rect 8298 8936 8354 8945
rect 8298 8871 8354 8880
rect 8312 8634 8340 8871
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7484 8090 7512 8434
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8128 8090 8156 8230
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 8404 4049 8432 13806
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8496 12374 8524 13262
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8496 11354 8524 12310
rect 8772 12073 8800 14010
rect 8758 12064 8814 12073
rect 8758 11999 8814 12008
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8772 11218 8800 11999
rect 8956 11354 8984 14855
rect 9140 14482 9168 14894
rect 9218 14855 9274 14864
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9232 12714 9260 13126
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9232 12442 9260 12650
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 9048 11558 9076 12242
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9140 11694 9168 12174
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8496 9897 8524 11154
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8482 9888 8538 9897
rect 8482 9823 8538 9832
rect 8496 8566 8524 9823
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8588 7546 8616 11018
rect 8772 10266 8800 11154
rect 9048 10810 9076 11494
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8956 8498 8984 9114
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8956 8090 8984 8434
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8588 7342 8616 7482
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8390 4040 8446 4049
rect 8390 3975 8446 3984
rect 6182 3496 6238 3505
rect 6182 3431 6238 3440
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 9324 1465 9352 15864
rect 9416 15706 9444 16050
rect 10060 15706 10088 17002
rect 10692 16992 10744 16998
rect 10690 16960 10692 16969
rect 10744 16960 10746 16969
rect 10289 16892 10585 16912
rect 10690 16895 10746 16904
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16590 10732 16895
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10704 16250 10732 16526
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10796 15706 10824 16662
rect 10980 16658 11008 20182
rect 11164 19922 11192 20402
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11348 20097 11376 20198
rect 11334 20088 11390 20097
rect 11334 20023 11390 20032
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 11164 18329 11192 19178
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11348 18426 11376 18770
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11336 18420 11388 18426
rect 11336 18362 11388 18368
rect 11150 18320 11206 18329
rect 11060 18284 11112 18290
rect 11150 18255 11206 18264
rect 11060 18226 11112 18232
rect 11072 17746 11100 18226
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 11152 17536 11204 17542
rect 11072 17484 11152 17490
rect 11072 17478 11204 17484
rect 11072 17462 11192 17478
rect 11072 16658 11100 17462
rect 11150 17232 11206 17241
rect 11256 17202 11284 18158
rect 11348 17338 11376 18362
rect 11440 17882 11468 18702
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11150 17167 11206 17176
rect 11244 17196 11296 17202
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10980 15910 11008 16594
rect 11072 16454 11100 16594
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11164 16114 11192 17167
rect 11244 17138 11296 17144
rect 11440 16794 11468 17818
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 11348 15706 11376 15982
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 9416 15502 9444 15642
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9496 15156 9548 15162
rect 9692 15144 9720 15506
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9548 15116 9720 15144
rect 9496 15098 9548 15104
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 9416 14278 9444 14826
rect 9784 14634 9812 15302
rect 9600 14606 9812 14634
rect 10060 14618 10088 15642
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10520 15162 10548 15438
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10048 14612 10100 14618
rect 9600 14550 9628 14606
rect 10048 14554 10100 14560
rect 10704 14550 10732 15098
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 10692 14544 10744 14550
rect 10692 14486 10744 14492
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9588 14272 9640 14278
rect 9640 14220 9720 14226
rect 9588 14214 9720 14220
rect 9600 14198 9720 14214
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9600 11694 9628 13398
rect 9692 12986 9720 14198
rect 10704 14074 10732 14486
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10888 13802 10916 15506
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11072 14498 11100 15302
rect 11334 14920 11390 14929
rect 11334 14855 11390 14864
rect 10980 14482 11100 14498
rect 10968 14476 11100 14482
rect 11020 14470 11100 14476
rect 10968 14418 11020 14424
rect 11348 14074 11376 14855
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 10876 13796 10928 13802
rect 10876 13738 10928 13744
rect 10138 13696 10194 13705
rect 10138 13631 10194 13640
rect 10152 13530 10180 13631
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 9770 13424 9826 13433
rect 9770 13359 9826 13368
rect 10048 13388 10100 13394
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 9654 9720 11562
rect 9784 10810 9812 13359
rect 10048 13330 10100 13336
rect 10060 12322 10088 13330
rect 10152 12986 10180 13466
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10416 12912 10468 12918
rect 10414 12880 10416 12889
rect 10468 12880 10470 12889
rect 10888 12850 10916 13194
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 10980 12850 11008 13126
rect 10414 12815 10470 12824
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10784 12640 10836 12646
rect 10784 12582 10836 12588
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10796 12442 10824 12582
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10980 12374 11008 12786
rect 10968 12368 11020 12374
rect 10060 12294 10180 12322
rect 10968 12310 11020 12316
rect 10152 12102 10180 12294
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10152 11393 10180 12038
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10138 11384 10194 11393
rect 10289 11376 10585 11396
rect 10796 11354 10824 12174
rect 10980 11898 11008 12310
rect 11440 12306 11468 13126
rect 11532 12753 11560 18022
rect 11624 16658 11652 19450
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11716 16590 11744 23276
rect 12256 21956 12308 21962
rect 12256 21898 12308 21904
rect 12268 21622 12296 21898
rect 12360 21690 12388 24074
rect 12452 24070 12480 24686
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12820 24410 12848 24550
rect 12808 24404 12860 24410
rect 12808 24346 12860 24352
rect 12716 24268 12768 24274
rect 12716 24210 12768 24216
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12452 23633 12480 24006
rect 12728 23798 12756 24210
rect 12820 23866 12848 24346
rect 12808 23860 12860 23866
rect 12808 23802 12860 23808
rect 12716 23792 12768 23798
rect 12716 23734 12768 23740
rect 12624 23656 12676 23662
rect 12438 23624 12494 23633
rect 12624 23598 12676 23604
rect 12438 23559 12494 23568
rect 12636 22982 12664 23598
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12636 22574 12664 22918
rect 12728 22642 12756 23734
rect 13004 23497 13032 24822
rect 13082 24783 13138 24792
rect 12990 23488 13046 23497
rect 12990 23423 13046 23432
rect 13004 23254 13032 23423
rect 12992 23248 13044 23254
rect 12992 23190 13044 23196
rect 13004 22778 13032 23190
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12624 22568 12676 22574
rect 12624 22510 12676 22516
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 12440 21004 12492 21010
rect 12440 20946 12492 20952
rect 12452 20618 12480 20946
rect 12532 20868 12584 20874
rect 12532 20810 12584 20816
rect 12360 20602 12480 20618
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 12348 20596 12480 20602
rect 12400 20590 12480 20596
rect 12348 20538 12400 20544
rect 11900 19514 11928 20538
rect 12544 20482 12572 20810
rect 12360 20466 12572 20482
rect 12348 20460 12572 20466
rect 12400 20454 12572 20460
rect 12348 20402 12400 20408
rect 12820 20398 12848 21830
rect 12912 21146 12940 21966
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12716 20324 12768 20330
rect 12716 20266 12768 20272
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 11886 19408 11942 19417
rect 11886 19343 11942 19352
rect 11900 19310 11928 19343
rect 11888 19304 11940 19310
rect 12728 19281 12756 20266
rect 13004 20058 13032 20878
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12820 19514 12848 19858
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 11888 19246 11940 19252
rect 12714 19272 12770 19281
rect 11980 19236 12032 19242
rect 12714 19207 12770 19216
rect 11980 19178 12032 19184
rect 11992 18766 12020 19178
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11992 18426 12020 18702
rect 12544 18630 12572 18838
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 12176 18222 12204 18566
rect 12544 18222 12572 18566
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12532 18216 12584 18222
rect 12584 18176 12664 18204
rect 12532 18158 12584 18164
rect 12176 17678 12204 18158
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12544 16590 12572 16934
rect 12636 16590 12664 18176
rect 12990 17232 13046 17241
rect 12990 17167 12992 17176
rect 13044 17167 13046 17176
rect 12992 17138 13044 17144
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12176 15910 12204 16526
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11716 14618 11744 15506
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11808 14890 11836 15438
rect 11900 15162 11928 15438
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11796 14884 11848 14890
rect 11796 14826 11848 14832
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 12084 14550 12112 14758
rect 12072 14544 12124 14550
rect 12072 14486 12124 14492
rect 11612 14272 11664 14278
rect 11610 14240 11612 14249
rect 11664 14240 11666 14249
rect 11610 14175 11666 14184
rect 11624 14074 11652 14175
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 12084 14006 12112 14486
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 12176 13394 12204 15846
rect 12268 15366 12296 16390
rect 12544 15706 12572 16526
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12636 15638 12664 16526
rect 13096 15706 13124 24783
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 13188 21690 13216 22034
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 13372 21146 13400 27520
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13740 23746 13768 24006
rect 13740 23718 13860 23746
rect 13740 23662 13768 23718
rect 13728 23656 13780 23662
rect 13728 23598 13780 23604
rect 13832 23322 13860 23718
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 13544 22432 13596 22438
rect 13544 22374 13596 22380
rect 13556 21350 13584 22374
rect 13648 22166 13676 22510
rect 13820 22432 13872 22438
rect 13820 22374 13872 22380
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 13648 21554 13676 22102
rect 13728 22024 13780 22030
rect 13832 21978 13860 22374
rect 13780 21972 13860 21978
rect 13728 21966 13860 21972
rect 13740 21950 13860 21966
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13174 21040 13230 21049
rect 13174 20975 13176 20984
rect 13228 20975 13230 20984
rect 13176 20946 13228 20952
rect 13188 20262 13216 20946
rect 13372 20602 13400 21082
rect 13556 20942 13584 21286
rect 13648 21146 13676 21490
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13820 21140 13872 21146
rect 13820 21082 13872 21088
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13832 20874 13860 21082
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13832 20466 13860 20810
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 13360 20392 13412 20398
rect 13924 20346 13952 27520
rect 14186 25256 14242 25265
rect 14186 25191 14242 25200
rect 14200 24410 14228 25191
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 13360 20334 13412 20340
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13188 16998 13216 20198
rect 13372 19310 13400 20334
rect 13740 20318 13952 20346
rect 14108 20330 14136 20742
rect 14096 20324 14148 20330
rect 13740 19990 13768 20318
rect 14096 20266 14148 20272
rect 14188 20324 14240 20330
rect 14188 20266 14240 20272
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13556 18306 13584 19858
rect 13740 19530 13768 19926
rect 14108 19854 14136 20266
rect 14200 19990 14228 20266
rect 14188 19984 14240 19990
rect 14188 19926 14240 19932
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 13648 19514 13768 19530
rect 13636 19508 13768 19514
rect 13688 19502 13768 19508
rect 13636 19450 13688 19456
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 13924 18970 13952 19178
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13556 18278 13676 18306
rect 13544 18148 13596 18154
rect 13544 18090 13596 18096
rect 13556 17898 13584 18090
rect 13464 17882 13584 17898
rect 13464 17876 13596 17882
rect 13464 17870 13544 17876
rect 13464 17202 13492 17870
rect 13544 17818 13596 17824
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13556 17338 13584 17682
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13176 16992 13228 16998
rect 13176 16934 13228 16940
rect 13188 15994 13216 16934
rect 13464 16726 13492 17138
rect 13648 16726 13676 18278
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14384 17882 14412 18022
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14384 17202 14412 17818
rect 14568 17241 14596 27520
rect 15120 25242 15148 27520
rect 14844 25214 15148 25242
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14660 19514 14688 19790
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14554 17232 14610 17241
rect 14372 17196 14424 17202
rect 14554 17167 14610 17176
rect 14372 17138 14424 17144
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13452 16720 13504 16726
rect 13636 16720 13688 16726
rect 13452 16662 13504 16668
rect 13634 16688 13636 16697
rect 13688 16688 13690 16697
rect 13634 16623 13690 16632
rect 13648 16114 13676 16623
rect 13832 16572 13860 16730
rect 14200 16590 14228 16934
rect 13740 16544 13860 16572
rect 14188 16584 14240 16590
rect 13740 16182 13768 16544
rect 14188 16526 14240 16532
rect 14200 16250 14228 16526
rect 14188 16244 14240 16250
rect 14188 16186 14240 16192
rect 13728 16176 13780 16182
rect 13728 16118 13780 16124
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13188 15966 13308 15994
rect 14384 15978 14412 17138
rect 14844 16794 14872 25214
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15672 24857 15700 27520
rect 15658 24848 15714 24857
rect 15658 24783 15714 24792
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15476 23656 15528 23662
rect 15476 23598 15528 23604
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15304 22574 15332 23054
rect 15382 22672 15438 22681
rect 15382 22607 15438 22616
rect 15292 22568 15344 22574
rect 15212 22516 15292 22522
rect 15212 22510 15344 22516
rect 15212 22494 15332 22510
rect 15212 22166 15240 22494
rect 15304 22445 15332 22494
rect 15396 22234 15424 22607
rect 15384 22228 15436 22234
rect 15384 22170 15436 22176
rect 15200 22160 15252 22166
rect 15200 22102 15252 22108
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15200 21412 15252 21418
rect 15200 21354 15252 21360
rect 15212 20890 15240 21354
rect 15290 21312 15346 21321
rect 15290 21247 15346 21256
rect 15304 21146 15332 21247
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 15212 20862 15332 20890
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15304 20602 15332 20862
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15304 19854 15332 20538
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19417 15332 19654
rect 15290 19408 15346 19417
rect 15290 19343 15346 19352
rect 15290 18864 15346 18873
rect 15346 18822 15424 18850
rect 15290 18799 15292 18808
rect 15344 18799 15346 18808
rect 15292 18770 15344 18776
rect 15290 18728 15346 18737
rect 15290 18663 15346 18672
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15304 18426 15332 18663
rect 15396 18426 15424 18822
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15304 18222 15332 18362
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12268 14482 12296 15302
rect 12348 14884 12400 14890
rect 12624 14884 12676 14890
rect 12400 14844 12480 14872
rect 12348 14826 12400 14832
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12360 13410 12388 14554
rect 12452 13530 12480 14844
rect 12624 14826 12676 14832
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 12164 13388 12216 13394
rect 12360 13382 12480 13410
rect 12164 13330 12216 13336
rect 11900 12986 11928 13330
rect 12452 12986 12480 13382
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12544 12782 12572 14758
rect 12636 14618 12664 14826
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12636 14482 12664 14554
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12636 13734 12664 14418
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12636 13462 12664 13670
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12636 13258 12664 13398
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12820 13138 12848 14758
rect 12912 13530 12940 15302
rect 13096 15162 13124 15642
rect 13280 15570 13308 15966
rect 14188 15972 14240 15978
rect 14188 15914 14240 15920
rect 14372 15972 14424 15978
rect 14372 15914 14424 15920
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13280 14822 13308 15506
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13372 14482 13400 15438
rect 14200 15434 14228 15914
rect 14384 15706 14412 15914
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14188 15428 14240 15434
rect 14188 15370 14240 15376
rect 14200 15162 14228 15370
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14292 14958 14320 15302
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14292 14618 14320 14894
rect 14384 14890 14412 15642
rect 15488 15638 15516 23598
rect 15934 23352 15990 23361
rect 15934 23287 15990 23296
rect 15568 23180 15620 23186
rect 15568 23122 15620 23128
rect 15580 22438 15608 23122
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15658 20088 15714 20097
rect 15658 20023 15714 20032
rect 15672 19990 15700 20023
rect 15660 19984 15712 19990
rect 15660 19926 15712 19932
rect 15672 19514 15700 19926
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15580 18902 15608 19246
rect 15948 19174 15976 23287
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 16040 18970 16068 19994
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 16132 18290 16160 23598
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 15752 16992 15804 16998
rect 15750 16960 15752 16969
rect 15804 16960 15806 16969
rect 15750 16895 15806 16904
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15304 15473 15332 15506
rect 15290 15464 15346 15473
rect 15290 15399 15346 15408
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 15162 15332 15399
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14384 14618 14412 14826
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13372 14074 13400 14418
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12636 13110 12848 13138
rect 12164 12776 12216 12782
rect 11518 12744 11574 12753
rect 11518 12679 11574 12688
rect 12162 12744 12164 12753
rect 12532 12776 12584 12782
rect 12216 12744 12218 12753
rect 12532 12718 12584 12724
rect 12162 12679 12218 12688
rect 12544 12442 12572 12718
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 11900 11898 11928 12174
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12176 11898 12204 12038
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12360 11354 12388 11630
rect 10138 11319 10194 11328
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 10874 11248 10930 11257
rect 10874 11183 10930 11192
rect 10968 11212 11020 11218
rect 10692 11144 10744 11150
rect 10230 11112 10286 11121
rect 10692 11086 10744 11092
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10230 11047 10232 11056
rect 10284 11047 10286 11056
rect 10232 11018 10284 11024
rect 10704 10810 10732 11086
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 9956 10464 10008 10470
rect 9954 10432 9956 10441
rect 10008 10432 10010 10441
rect 9954 10367 10010 10376
rect 10060 10266 10088 10746
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 10232 10192 10284 10198
rect 10232 10134 10284 10140
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 10152 9382 10180 9998
rect 10244 9722 10272 10134
rect 10796 9926 10824 11086
rect 10888 11014 10916 11183
rect 10968 11154 11020 11160
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10888 10674 10916 10950
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10888 10198 10916 10610
rect 10980 10418 11008 11154
rect 12452 10810 12480 12174
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12544 11354 12572 11630
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12544 10674 12572 11290
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12162 10568 12218 10577
rect 12162 10503 12164 10512
rect 12216 10503 12218 10512
rect 12164 10474 12216 10480
rect 11060 10464 11112 10470
rect 10980 10412 11060 10418
rect 10980 10406 11112 10412
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 10980 10390 11100 10406
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10152 9042 10180 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10796 9042 10824 9862
rect 10980 9586 11008 10390
rect 11532 9926 11560 10406
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11886 9480 11942 9489
rect 11886 9415 11942 9424
rect 11900 9178 11928 9415
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10152 8566 10180 8978
rect 10612 8634 10640 8978
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 9310 1456 9366 1465
rect 9310 1391 9366 1400
rect 12636 1329 12664 13110
rect 12912 12986 12940 13466
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13740 13002 13768 13262
rect 13832 13002 13860 14554
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 16118 13968 16174 13977
rect 16118 13903 16174 13912
rect 16132 13870 16160 13903
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 13740 12974 13860 13002
rect 16224 12986 16252 27520
rect 16776 24562 16804 27520
rect 16500 24534 16804 24562
rect 16500 23866 16528 24534
rect 16762 24440 16818 24449
rect 16762 24375 16764 24384
rect 16816 24375 16818 24384
rect 16764 24346 16816 24352
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16488 23860 16540 23866
rect 16488 23802 16540 23808
rect 16408 23582 16620 23610
rect 16776 23594 16804 24210
rect 16302 22536 16358 22545
rect 16302 22471 16358 22480
rect 16316 22234 16344 22471
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16316 19961 16344 20198
rect 16302 19952 16358 19961
rect 16302 19887 16358 19896
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16316 19514 16344 19790
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16304 16040 16356 16046
rect 16302 16008 16304 16017
rect 16356 16008 16358 16017
rect 16302 15943 16358 15952
rect 16408 13938 16436 23582
rect 16592 23526 16620 23582
rect 16764 23588 16816 23594
rect 16764 23530 16816 23536
rect 16580 23520 16632 23526
rect 16580 23462 16632 23468
rect 16670 23488 16726 23497
rect 16670 23423 16726 23432
rect 16684 23322 16712 23423
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16776 16114 16804 23530
rect 17420 23361 17448 27520
rect 17866 24848 17922 24857
rect 17866 24783 17922 24792
rect 17880 24410 17908 24783
rect 17868 24404 17920 24410
rect 17868 24346 17920 24352
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 17590 23624 17646 23633
rect 17590 23559 17646 23568
rect 17406 23352 17462 23361
rect 17406 23287 17462 23296
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 17604 13462 17632 23559
rect 17696 23526 17724 24210
rect 17972 23882 18000 27520
rect 18524 24449 18552 27520
rect 19076 24857 19104 27520
rect 19628 25786 19656 27520
rect 19352 25758 19656 25786
rect 19062 24848 19118 24857
rect 19062 24783 19118 24792
rect 19062 24712 19118 24721
rect 19062 24647 19118 24656
rect 18510 24440 18566 24449
rect 19076 24410 19104 24647
rect 18510 24375 18566 24384
rect 19064 24404 19116 24410
rect 19064 24346 19116 24352
rect 18880 24268 18932 24274
rect 18880 24210 18932 24216
rect 17880 23866 18000 23882
rect 17868 23860 18000 23866
rect 17920 23854 18000 23860
rect 17868 23802 17920 23808
rect 18892 23730 18920 24210
rect 19352 24120 19380 25758
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19982 24848 20038 24857
rect 19982 24783 20038 24792
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19260 24092 19380 24120
rect 19260 23866 19288 24092
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 18328 23724 18380 23730
rect 18328 23666 18380 23672
rect 18880 23724 18932 23730
rect 18880 23666 18932 23672
rect 17684 23520 17736 23526
rect 17684 23462 17736 23468
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 16212 12980 16264 12986
rect 13740 12918 13768 12974
rect 16212 12922 16264 12928
rect 17420 12918 17448 13330
rect 13728 12912 13780 12918
rect 16764 12912 16816 12918
rect 13728 12854 13780 12860
rect 16762 12880 16764 12889
rect 17408 12912 17460 12918
rect 16816 12880 16818 12889
rect 13084 12844 13136 12850
rect 16762 12815 16818 12824
rect 16946 12880 17002 12889
rect 17408 12854 17460 12860
rect 18340 12850 18368 23666
rect 19156 23656 19208 23662
rect 19154 23624 19156 23633
rect 19208 23624 19210 23633
rect 19154 23559 19210 23568
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18616 12889 18644 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19996 23322 20024 24783
rect 20272 23866 20300 27520
rect 20824 24721 20852 27520
rect 21376 24857 21404 27520
rect 21362 24848 21418 24857
rect 21362 24783 21418 24792
rect 20810 24712 20866 24721
rect 20810 24647 20866 24656
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20442 24032 20498 24041
rect 20442 23967 20498 23976
rect 20456 23866 20484 23967
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20260 23656 20312 23662
rect 20260 23598 20312 23604
rect 19984 23316 20036 23322
rect 19984 23258 20036 23264
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 19444 22438 19472 23122
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 18602 12880 18658 12889
rect 16946 12815 16948 12824
rect 13084 12786 13136 12792
rect 17000 12815 17002 12824
rect 18328 12844 18380 12850
rect 16948 12786 17000 12792
rect 18602 12815 18658 12824
rect 18328 12786 18380 12792
rect 13096 12442 13124 12786
rect 14004 12776 14056 12782
rect 13266 12744 13322 12753
rect 14004 12718 14056 12724
rect 16672 12776 16724 12782
rect 18052 12776 18104 12782
rect 16672 12718 16724 12724
rect 18050 12744 18052 12753
rect 18104 12744 18106 12753
rect 13266 12679 13322 12688
rect 13280 12442 13308 12679
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13820 12232 13872 12238
rect 14016 12209 14044 12718
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 13820 12174 13872 12180
rect 14002 12200 14058 12209
rect 13832 11558 13860 12174
rect 14002 12135 14058 12144
rect 14384 11898 14412 12242
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 13820 11552 13872 11558
rect 13740 11512 13820 11540
rect 13740 11286 13768 11512
rect 13820 11494 13872 11500
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 13728 11280 13780 11286
rect 14108 11257 14136 11290
rect 13728 11222 13780 11228
rect 14094 11248 14150 11257
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12714 10976 12770 10985
rect 12714 10911 12770 10920
rect 12728 10470 12756 10911
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 10266 12756 10406
rect 12820 10266 12848 11154
rect 13740 10810 13768 11222
rect 14094 11183 14150 11192
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 16684 10169 16712 12718
rect 18050 12679 18106 12688
rect 19444 11257 19472 22374
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 18786 11248 18842 11257
rect 18512 11212 18564 11218
rect 18786 11183 18788 11192
rect 18512 11154 18564 11160
rect 18840 11183 18842 11192
rect 19430 11248 19486 11257
rect 19430 11183 19486 11192
rect 18788 11154 18840 11160
rect 18524 11121 18552 11154
rect 18510 11112 18566 11121
rect 18510 11047 18566 11056
rect 18524 10810 18552 11047
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 20166 10704 20222 10713
rect 20166 10639 20222 10648
rect 20180 10606 20208 10639
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 20272 10169 20300 23598
rect 20916 23526 20944 24210
rect 21928 24041 21956 27520
rect 22480 24410 22508 27520
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 21914 24032 21970 24041
rect 21914 23967 21970 23976
rect 23124 23905 23152 27520
rect 21546 23896 21602 23905
rect 21546 23831 21548 23840
rect 21600 23831 21602 23840
rect 23110 23896 23166 23905
rect 23110 23831 23166 23840
rect 21548 23802 21600 23808
rect 21364 23656 21416 23662
rect 21364 23598 21416 23604
rect 20904 23520 20956 23526
rect 20904 23462 20956 23468
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20732 13297 20760 13806
rect 20718 13288 20774 13297
rect 20718 13223 20774 13232
rect 16670 10160 16726 10169
rect 19154 10160 19210 10169
rect 16670 10095 16726 10104
rect 18880 10124 18932 10130
rect 19154 10095 19156 10104
rect 18880 10066 18932 10072
rect 19208 10095 19210 10104
rect 20258 10160 20314 10169
rect 20258 10095 20314 10104
rect 19156 10066 19208 10072
rect 18892 10033 18920 10066
rect 18878 10024 18934 10033
rect 18878 9959 18934 9968
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 18892 9722 18920 9959
rect 18880 9716 18932 9722
rect 18880 9658 18932 9664
rect 20916 9602 20944 23462
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 21008 13938 21036 14894
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 21376 10674 21404 23598
rect 23480 23588 23532 23594
rect 23480 23530 23532 23536
rect 21822 15192 21878 15201
rect 21822 15127 21824 15136
rect 21876 15127 21878 15136
rect 21824 15098 21876 15104
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 20640 9586 20944 9602
rect 20628 9580 20944 9586
rect 20680 9574 20944 9580
rect 20628 9522 20680 9528
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 19352 8401 19380 9454
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19338 8392 19394 8401
rect 19338 8327 19394 8336
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 22284 7336 22336 7342
rect 22282 7304 22284 7313
rect 22336 7304 22338 7313
rect 22282 7239 22338 7248
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 22742 6896 22798 6905
rect 22742 6831 22744 6840
rect 22796 6831 22798 6840
rect 22744 6802 22796 6808
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 22756 6458 22784 6802
rect 23492 6746 23520 23530
rect 23572 21412 23624 21418
rect 23572 21354 23624 21360
rect 23584 7546 23612 21354
rect 23676 15201 23704 27520
rect 24228 21418 24256 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24780 23594 24808 27520
rect 25332 27418 25360 27520
rect 24964 27390 25360 27418
rect 24768 23588 24820 23594
rect 24768 23530 24820 23536
rect 24766 23488 24822 23497
rect 24766 23423 24822 23432
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24216 21412 24268 21418
rect 24216 21354 24268 21360
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 23662 15192 23718 15201
rect 24289 15184 24585 15204
rect 23662 15127 23718 15136
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23846 6896 23902 6905
rect 23846 6831 23902 6840
rect 23400 6730 23520 6746
rect 23388 6724 23520 6730
rect 23440 6718 23520 6724
rect 23388 6666 23440 6672
rect 23860 6458 23888 6831
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 22744 6452 22796 6458
rect 22744 6394 22796 6400
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 23664 6248 23716 6254
rect 23662 6216 23664 6225
rect 23716 6216 23718 6225
rect 23662 6151 23718 6160
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 24030 5808 24086 5817
rect 24030 5743 24032 5752
rect 24084 5743 24086 5752
rect 24032 5714 24084 5720
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 24044 5370 24072 5714
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24780 5370 24808 23423
rect 24860 21412 24912 21418
rect 24860 21354 24912 21360
rect 24872 5914 24900 21354
rect 24964 6905 24992 27390
rect 25976 21418 26004 27520
rect 26528 23497 26556 27520
rect 27080 26194 27108 27520
rect 26712 26166 27108 26194
rect 26514 23488 26570 23497
rect 26514 23423 26570 23432
rect 25964 21412 26016 21418
rect 25964 21354 26016 21360
rect 26712 21298 26740 26166
rect 26252 21270 26740 21298
rect 24950 6896 25006 6905
rect 24950 6831 25006 6840
rect 24860 5908 24912 5914
rect 24860 5850 24912 5856
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24582 5264 24638 5273
rect 24582 5199 24638 5208
rect 24596 5166 24624 5199
rect 24584 5160 24636 5166
rect 24584 5102 24636 5108
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 26252 4865 26280 21270
rect 27632 17649 27660 27520
rect 27618 17640 27674 17649
rect 27618 17575 27674 17584
rect 24766 4856 24822 4865
rect 24766 4791 24768 4800
rect 24820 4791 24822 4800
rect 26238 4856 26294 4865
rect 26238 4791 26294 4800
rect 24768 4762 24820 4768
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24584 4208 24636 4214
rect 24582 4176 24584 4185
rect 24636 4176 24638 4185
rect 24688 4162 24716 4626
rect 24638 4134 24716 4162
rect 24582 4111 24638 4120
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 23202 3496 23258 3505
rect 23202 3431 23258 3440
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 13910 2952 13966 2961
rect 13910 2887 13966 2896
rect 12622 1320 12678 1329
rect 12622 1255 12678 1264
rect 13924 480 13952 2887
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 23216 480 23244 3431
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 3330 368 3386 377
rect 3330 303 3386 312
rect 4618 0 4674 480
rect 13910 0 13966 480
rect 23202 0 23258 480
<< via2 >>
rect 3422 27648 3478 27704
rect 846 22072 902 22128
rect 1398 20984 1454 21040
rect 1582 24268 1638 24304
rect 1582 24248 1584 24268
rect 1584 24248 1636 24268
rect 1636 24248 1638 24268
rect 1858 24520 1914 24576
rect 1858 23568 1914 23624
rect 1766 21664 1822 21720
rect 1766 21256 1822 21312
rect 2042 24112 2098 24168
rect 2042 23724 2098 23760
rect 2042 23704 2044 23724
rect 2044 23704 2096 23724
rect 2096 23704 2098 23724
rect 2410 22924 2412 22944
rect 2412 22924 2464 22944
rect 2464 22924 2466 22944
rect 2410 22888 2466 22924
rect 2870 23432 2926 23488
rect 2778 22752 2834 22808
rect 2318 21956 2374 21992
rect 2318 21936 2320 21956
rect 2320 21936 2372 21956
rect 2372 21936 2374 21956
rect 2410 21140 2466 21176
rect 2410 21120 2412 21140
rect 2412 21120 2464 21140
rect 2464 21120 2466 21140
rect 2318 20460 2374 20496
rect 2318 20440 2320 20460
rect 2320 20440 2372 20460
rect 2372 20440 2374 20460
rect 2778 20848 2834 20904
rect 2778 20304 2834 20360
rect 2686 20204 2688 20224
rect 2688 20204 2740 20224
rect 2740 20204 2742 20224
rect 2686 20168 2742 20204
rect 2962 22208 3018 22264
rect 3514 27104 3570 27160
rect 3422 26424 3478 26480
rect 3238 25880 3294 25936
rect 3514 25220 3570 25256
rect 3514 25200 3516 25220
rect 3516 25200 3568 25220
rect 3568 25200 3570 25220
rect 3146 22500 3202 22536
rect 3146 22480 3148 22500
rect 3148 22480 3200 22500
rect 3200 22480 3202 22500
rect 3054 21528 3110 21584
rect 2870 19896 2926 19952
rect 2318 19796 2320 19816
rect 2320 19796 2372 19816
rect 2372 19796 2374 19816
rect 2318 19760 2374 19796
rect 1490 17720 1546 17776
rect 2042 18944 2098 19000
rect 1766 18164 1768 18184
rect 1768 18164 1820 18184
rect 1820 18164 1822 18184
rect 1766 18128 1822 18164
rect 2410 17720 2466 17776
rect 1674 17448 1730 17504
rect 294 17040 350 17096
rect 1582 16632 1638 16688
rect 1490 15952 1546 16008
rect 2134 17584 2190 17640
rect 2318 17060 2374 17096
rect 2318 17040 2320 17060
rect 2320 17040 2372 17060
rect 2372 17040 2374 17060
rect 2962 19080 3018 19136
rect 3514 21528 3570 21584
rect 3422 21392 3478 21448
rect 3790 25200 3846 25256
rect 4250 24012 4252 24032
rect 4252 24012 4304 24032
rect 4304 24012 4306 24032
rect 4250 23976 4306 24012
rect 3330 19080 3386 19136
rect 3146 18536 3202 18592
rect 3514 18264 3570 18320
rect 3698 20984 3754 21040
rect 3422 17720 3478 17776
rect 3054 17312 3110 17368
rect 3330 17176 3386 17232
rect 2870 17040 2926 17096
rect 1674 13096 1730 13152
rect 1858 13776 1914 13832
rect 2134 12980 2190 13016
rect 2134 12960 2136 12980
rect 2136 12960 2188 12980
rect 2188 12960 2190 12980
rect 2778 14864 2834 14920
rect 1766 12164 1822 12200
rect 1766 12144 1768 12164
rect 1768 12144 1820 12164
rect 1820 12144 1822 12164
rect 1766 10240 1822 10296
rect 2502 10784 2558 10840
rect 2686 12824 2742 12880
rect 2594 10240 2650 10296
rect 3146 16904 3202 16960
rect 3606 17040 3662 17096
rect 4066 20168 4122 20224
rect 4526 23024 4582 23080
rect 4342 19352 4398 19408
rect 4066 18692 4122 18728
rect 4066 18672 4068 18692
rect 4068 18672 4120 18692
rect 4120 18672 4122 18692
rect 3790 17040 3846 17096
rect 3330 13776 3386 13832
rect 2962 9968 3018 10024
rect 2686 9016 2742 9072
rect 2042 3848 2098 3904
rect 2594 2916 2650 2952
rect 2594 2896 2596 2916
rect 2596 2896 2648 2916
rect 2648 2896 2650 2916
rect 3514 11192 3570 11248
rect 3514 10512 3570 10568
rect 3422 9016 3478 9072
rect 3698 11464 3754 11520
rect 3698 8200 3754 8256
rect 4066 16088 4122 16144
rect 3974 15544 4030 15600
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5998 24792 6054 24848
rect 5354 24384 5410 24440
rect 5170 24248 5226 24304
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5170 22888 5226 22944
rect 4986 22072 5042 22128
rect 4434 18964 4490 19000
rect 4434 18944 4436 18964
rect 4436 18944 4488 18964
rect 4488 18944 4490 18964
rect 4342 18164 4344 18184
rect 4344 18164 4396 18184
rect 4396 18164 4398 18184
rect 4342 18128 4398 18164
rect 4250 17448 4306 17504
rect 3974 12688 4030 12744
rect 3882 11736 3938 11792
rect 4066 12416 4122 12472
rect 4066 9988 4122 10024
rect 4066 9968 4068 9988
rect 4068 9968 4120 9988
rect 4120 9968 4122 9988
rect 3974 3304 4030 3360
rect 3790 2624 3846 2680
rect 4526 17856 4582 17912
rect 4434 15816 4490 15872
rect 4802 17856 4858 17912
rect 4802 17584 4858 17640
rect 5170 21256 5226 21312
rect 4894 17040 4950 17096
rect 5170 17584 5226 17640
rect 5078 16632 5134 16688
rect 5078 15408 5134 15464
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5538 22616 5594 22672
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5446 21664 5502 21720
rect 5630 21256 5686 21312
rect 6274 21120 6330 21176
rect 6182 20984 6238 21040
rect 5538 20848 5594 20904
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5998 20596 6054 20632
rect 5998 20576 6000 20596
rect 6000 20576 6052 20596
rect 6052 20576 6054 20596
rect 6826 24520 6882 24576
rect 7010 24656 7066 24712
rect 7102 23704 7158 23760
rect 7930 23568 7986 23624
rect 8114 23568 8170 23624
rect 7930 23432 7986 23488
rect 6918 23024 6974 23080
rect 6550 21256 6606 21312
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5538 19352 5594 19408
rect 5998 19080 6054 19136
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5354 15000 5410 15056
rect 4802 13912 4858 13968
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5262 12844 5318 12880
rect 5262 12824 5264 12844
rect 5264 12824 5316 12844
rect 5316 12824 5318 12844
rect 5446 12824 5502 12880
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5998 11736 6054 11792
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5630 10104 5686 10160
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 4894 9424 4950 9480
rect 5078 9444 5134 9480
rect 5078 9424 5080 9444
rect 5080 9424 5132 9444
rect 5132 9424 5134 9444
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 4618 3984 4674 4040
rect 4342 2080 4398 2136
rect 6274 19236 6330 19272
rect 6274 19216 6276 19236
rect 6276 19216 6328 19236
rect 6328 19216 6330 19236
rect 6642 18808 6698 18864
rect 6642 17448 6698 17504
rect 7010 19080 7066 19136
rect 6918 18808 6974 18864
rect 7286 18692 7342 18728
rect 7286 18672 7288 18692
rect 7288 18672 7340 18692
rect 7340 18672 7342 18692
rect 8850 24812 8906 24848
rect 8850 24792 8852 24812
rect 8852 24792 8904 24812
rect 8904 24792 8906 24812
rect 9770 24384 9826 24440
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 9954 24112 10010 24168
rect 9402 23432 9458 23488
rect 9494 21936 9550 21992
rect 8850 20984 8906 21040
rect 9034 20596 9090 20632
rect 9034 20576 9036 20596
rect 9036 20576 9088 20596
rect 9088 20576 9090 20596
rect 8390 19916 8446 19952
rect 8390 19896 8392 19916
rect 8392 19896 8444 19916
rect 8444 19896 8446 19916
rect 8022 19780 8078 19816
rect 8022 19760 8024 19780
rect 8024 19760 8076 19780
rect 8076 19760 8078 19780
rect 6550 14320 6606 14376
rect 6458 13640 6514 13696
rect 7194 16632 7250 16688
rect 9678 20440 9734 20496
rect 8850 19080 8906 19136
rect 7930 17620 7932 17640
rect 7932 17620 7984 17640
rect 7984 17620 7986 17640
rect 7930 17584 7986 17620
rect 7654 17448 7710 17504
rect 8482 17720 8538 17776
rect 8298 17484 8300 17504
rect 8300 17484 8352 17504
rect 8352 17484 8354 17504
rect 8298 17448 8354 17484
rect 8206 16940 8208 16960
rect 8208 16940 8260 16960
rect 8260 16940 8262 16960
rect 8206 16904 8262 16940
rect 7470 16632 7526 16688
rect 6826 15408 6882 15464
rect 6734 14884 6790 14920
rect 6734 14864 6736 14884
rect 6736 14864 6788 14884
rect 6788 14864 6790 14884
rect 7378 15020 7434 15056
rect 7378 15000 7380 15020
rect 7380 15000 7432 15020
rect 7432 15000 7434 15020
rect 10690 23568 10746 23624
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10874 23432 10930 23488
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10046 21528 10102 21584
rect 10690 21256 10746 21312
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10138 19116 10140 19136
rect 10140 19116 10192 19136
rect 10192 19116 10194 19136
rect 10138 19080 10194 19116
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 9310 17040 9366 17096
rect 7930 15544 7986 15600
rect 7470 13776 7526 13832
rect 8574 14184 8630 14240
rect 11702 23432 11758 23488
rect 11242 21392 11298 21448
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 9862 16088 9918 16144
rect 8942 14864 8998 14920
rect 6642 13368 6698 13424
rect 8022 13252 8078 13288
rect 8022 13232 8024 13252
rect 8024 13232 8076 13252
rect 8076 13232 8078 13252
rect 7470 12824 7526 12880
rect 6550 12316 6552 12336
rect 6552 12316 6604 12336
rect 6604 12316 6606 12336
rect 6550 12280 6606 12316
rect 6550 11500 6552 11520
rect 6552 11500 6604 11520
rect 6604 11500 6606 11520
rect 6550 11464 6606 11500
rect 7010 12008 7066 12064
rect 8298 12280 8354 12336
rect 7470 10648 7526 10704
rect 7746 10260 7802 10296
rect 7746 10240 7748 10260
rect 7748 10240 7800 10260
rect 7800 10240 7802 10260
rect 6826 9868 6828 9888
rect 6828 9868 6880 9888
rect 6880 9868 6882 9888
rect 6826 9832 6882 9868
rect 6642 9016 6698 9072
rect 6826 8336 6882 8392
rect 8298 8880 8354 8936
rect 8758 12008 8814 12064
rect 9218 14864 9274 14920
rect 8482 9832 8538 9888
rect 8390 3984 8446 4040
rect 6182 3440 6238 3496
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10690 16940 10692 16960
rect 10692 16940 10744 16960
rect 10744 16940 10746 16960
rect 10690 16904 10746 16940
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 11334 20032 11390 20088
rect 11150 18264 11206 18320
rect 11150 17176 11206 17232
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 11334 14864 11390 14920
rect 10138 13640 10194 13696
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 9770 13368 9826 13424
rect 10414 12860 10416 12880
rect 10416 12860 10468 12880
rect 10468 12860 10470 12880
rect 10414 12824 10470 12860
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10138 11328 10194 11384
rect 12438 23568 12494 23624
rect 13082 24792 13138 24848
rect 12990 23432 13046 23488
rect 11886 19352 11942 19408
rect 12714 19216 12770 19272
rect 12990 17196 13046 17232
rect 12990 17176 12992 17196
rect 12992 17176 13044 17196
rect 13044 17176 13046 17196
rect 11610 14220 11612 14240
rect 11612 14220 11664 14240
rect 11664 14220 11666 14240
rect 11610 14184 11666 14220
rect 13174 21004 13230 21040
rect 13174 20984 13176 21004
rect 13176 20984 13228 21004
rect 13228 20984 13230 21004
rect 14186 25200 14242 25256
rect 14554 17176 14610 17232
rect 13634 16668 13636 16688
rect 13636 16668 13688 16688
rect 13688 16668 13690 16688
rect 13634 16632 13690 16668
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15658 24792 15714 24848
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15382 22616 15438 22672
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15290 21256 15346 21312
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15290 19352 15346 19408
rect 15290 18828 15346 18864
rect 15290 18808 15292 18828
rect 15292 18808 15344 18828
rect 15344 18808 15346 18828
rect 15290 18672 15346 18728
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15934 23296 15990 23352
rect 15658 20032 15714 20088
rect 15750 16940 15752 16960
rect 15752 16940 15804 16960
rect 15804 16940 15806 16960
rect 15750 16904 15806 16940
rect 15290 15408 15346 15464
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 11518 12688 11574 12744
rect 12162 12724 12164 12744
rect 12164 12724 12216 12744
rect 12216 12724 12218 12744
rect 12162 12688 12218 12724
rect 10874 11192 10930 11248
rect 10230 11076 10286 11112
rect 10230 11056 10232 11076
rect 10232 11056 10284 11076
rect 10284 11056 10286 11076
rect 9954 10412 9956 10432
rect 9956 10412 10008 10432
rect 10008 10412 10010 10432
rect 9954 10376 10010 10412
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 12162 10532 12218 10568
rect 12162 10512 12164 10532
rect 12164 10512 12216 10532
rect 12216 10512 12218 10532
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 11886 9424 11942 9480
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 9310 1400 9366 1456
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 16118 13912 16174 13968
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 16762 24404 16818 24440
rect 16762 24384 16764 24404
rect 16764 24384 16816 24404
rect 16816 24384 16818 24404
rect 16302 22480 16358 22536
rect 16302 19896 16358 19952
rect 16302 15988 16304 16008
rect 16304 15988 16356 16008
rect 16356 15988 16358 16008
rect 16302 15952 16358 15988
rect 16670 23432 16726 23488
rect 17866 24792 17922 24848
rect 17590 23568 17646 23624
rect 17406 23296 17462 23352
rect 19062 24792 19118 24848
rect 19062 24656 19118 24712
rect 18510 24384 18566 24440
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19982 24792 20038 24848
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 16762 12860 16764 12880
rect 16764 12860 16816 12880
rect 16816 12860 16818 12880
rect 16762 12824 16818 12860
rect 16946 12844 17002 12880
rect 19154 23604 19156 23624
rect 19156 23604 19208 23624
rect 19208 23604 19210 23624
rect 19154 23568 19210 23604
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 21362 24792 21418 24848
rect 20810 24656 20866 24712
rect 20442 23976 20498 24032
rect 16946 12824 16948 12844
rect 16948 12824 17000 12844
rect 17000 12824 17002 12844
rect 18602 12824 18658 12880
rect 13266 12688 13322 12744
rect 18050 12724 18052 12744
rect 18052 12724 18104 12744
rect 18104 12724 18106 12744
rect 14002 12144 14058 12200
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 12714 10920 12770 10976
rect 14094 11192 14150 11248
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 18050 12688 18106 12724
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 18786 11212 18842 11248
rect 18786 11192 18788 11212
rect 18788 11192 18840 11212
rect 18840 11192 18842 11212
rect 19430 11192 19486 11248
rect 18510 11056 18566 11112
rect 20166 10648 20222 10704
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 21914 23976 21970 24032
rect 21546 23860 21602 23896
rect 21546 23840 21548 23860
rect 21548 23840 21600 23860
rect 21600 23840 21602 23860
rect 23110 23840 23166 23896
rect 20718 13232 20774 13288
rect 16670 10104 16726 10160
rect 19154 10124 19210 10160
rect 19154 10104 19156 10124
rect 19156 10104 19208 10124
rect 19208 10104 19210 10124
rect 20258 10104 20314 10160
rect 18878 9968 18934 10024
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 21822 15156 21878 15192
rect 21822 15136 21824 15156
rect 21824 15136 21876 15156
rect 21876 15136 21878 15156
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19338 8336 19394 8392
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 22282 7284 22284 7304
rect 22284 7284 22336 7304
rect 22336 7284 22338 7304
rect 22282 7248 22338 7284
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 22742 6860 22798 6896
rect 22742 6840 22744 6860
rect 22744 6840 22796 6860
rect 22796 6840 22798 6860
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 23432 24822 23488
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 23662 15136 23718 15192
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 23846 6840 23902 6896
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 23662 6196 23664 6216
rect 23664 6196 23716 6216
rect 23716 6196 23718 6216
rect 23662 6160 23718 6196
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 24030 5772 24086 5808
rect 24030 5752 24032 5772
rect 24032 5752 24084 5772
rect 24084 5752 24086 5772
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 26514 23432 26570 23488
rect 24950 6840 25006 6896
rect 24582 5208 24638 5264
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 27618 17584 27674 17640
rect 24766 4820 24822 4856
rect 24766 4800 24768 4820
rect 24768 4800 24820 4820
rect 24820 4800 24822 4820
rect 26238 4800 26294 4856
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24582 4156 24584 4176
rect 24584 4156 24636 4176
rect 24636 4156 24638 4176
rect 24582 4120 24638 4156
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 23202 3440 23258 3496
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 13910 2896 13966 2952
rect 12622 1264 12678 1320
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 3330 312 3386 368
<< metal3 >>
rect 0 27706 480 27736
rect 3417 27706 3483 27709
rect 0 27704 3483 27706
rect 0 27648 3422 27704
rect 3478 27648 3483 27704
rect 0 27646 3483 27648
rect 0 27616 480 27646
rect 3417 27643 3483 27646
rect 0 27162 480 27192
rect 3509 27162 3575 27165
rect 0 27160 3575 27162
rect 0 27104 3514 27160
rect 3570 27104 3575 27160
rect 0 27102 3575 27104
rect 0 27072 480 27102
rect 3509 27099 3575 27102
rect 0 26482 480 26512
rect 3417 26482 3483 26485
rect 0 26480 3483 26482
rect 0 26424 3422 26480
rect 3478 26424 3483 26480
rect 0 26422 3483 26424
rect 0 26392 480 26422
rect 3417 26419 3483 26422
rect 0 25938 480 25968
rect 3233 25938 3299 25941
rect 0 25936 3299 25938
rect 0 25880 3238 25936
rect 3294 25880 3299 25936
rect 0 25878 3299 25880
rect 0 25848 480 25878
rect 3233 25875 3299 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25258 480 25288
rect 3509 25258 3575 25261
rect 0 25256 3575 25258
rect 0 25200 3514 25256
rect 3570 25200 3575 25256
rect 0 25198 3575 25200
rect 0 25168 480 25198
rect 3509 25195 3575 25198
rect 3785 25258 3851 25261
rect 14181 25258 14247 25261
rect 3785 25256 14247 25258
rect 3785 25200 3790 25256
rect 3846 25200 14186 25256
rect 14242 25200 14247 25256
rect 3785 25198 14247 25200
rect 3785 25195 3851 25198
rect 14181 25195 14247 25198
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 5993 24850 6059 24853
rect 8845 24850 8911 24853
rect 5993 24848 8911 24850
rect 5993 24792 5998 24848
rect 6054 24792 8850 24848
rect 8906 24792 8911 24848
rect 5993 24790 8911 24792
rect 5993 24787 6059 24790
rect 8845 24787 8911 24790
rect 13077 24850 13143 24853
rect 15653 24850 15719 24853
rect 13077 24848 15719 24850
rect 13077 24792 13082 24848
rect 13138 24792 15658 24848
rect 15714 24792 15719 24848
rect 13077 24790 15719 24792
rect 13077 24787 13143 24790
rect 15653 24787 15719 24790
rect 17861 24850 17927 24853
rect 19057 24850 19123 24853
rect 17861 24848 19123 24850
rect 17861 24792 17866 24848
rect 17922 24792 19062 24848
rect 19118 24792 19123 24848
rect 17861 24790 19123 24792
rect 17861 24787 17927 24790
rect 19057 24787 19123 24790
rect 19977 24850 20043 24853
rect 21357 24850 21423 24853
rect 19977 24848 21423 24850
rect 19977 24792 19982 24848
rect 20038 24792 21362 24848
rect 21418 24792 21423 24848
rect 19977 24790 21423 24792
rect 19977 24787 20043 24790
rect 21357 24787 21423 24790
rect 0 24714 480 24744
rect 7005 24714 7071 24717
rect 0 24712 7071 24714
rect 0 24656 7010 24712
rect 7066 24656 7071 24712
rect 0 24654 7071 24656
rect 0 24624 480 24654
rect 7005 24651 7071 24654
rect 19057 24714 19123 24717
rect 20805 24714 20871 24717
rect 19057 24712 20871 24714
rect 19057 24656 19062 24712
rect 19118 24656 20810 24712
rect 20866 24656 20871 24712
rect 19057 24654 20871 24656
rect 19057 24651 19123 24654
rect 20805 24651 20871 24654
rect 1853 24578 1919 24581
rect 6821 24578 6887 24581
rect 1853 24576 6887 24578
rect 1853 24520 1858 24576
rect 1914 24520 6826 24576
rect 6882 24520 6887 24576
rect 1853 24518 6887 24520
rect 1853 24515 1919 24518
rect 6821 24515 6887 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 5349 24442 5415 24445
rect 9765 24442 9831 24445
rect 5349 24440 9831 24442
rect 5349 24384 5354 24440
rect 5410 24384 9770 24440
rect 9826 24384 9831 24440
rect 5349 24382 9831 24384
rect 5349 24379 5415 24382
rect 9765 24379 9831 24382
rect 16757 24442 16823 24445
rect 18505 24442 18571 24445
rect 16757 24440 18571 24442
rect 16757 24384 16762 24440
rect 16818 24384 18510 24440
rect 18566 24384 18571 24440
rect 16757 24382 18571 24384
rect 16757 24379 16823 24382
rect 18505 24379 18571 24382
rect 1577 24306 1643 24309
rect 5165 24306 5231 24309
rect 1577 24304 5231 24306
rect 1577 24248 1582 24304
rect 1638 24248 5170 24304
rect 5226 24248 5231 24304
rect 1577 24246 5231 24248
rect 1577 24243 1643 24246
rect 5165 24243 5231 24246
rect 2037 24170 2103 24173
rect 9949 24170 10015 24173
rect 2037 24168 10015 24170
rect 2037 24112 2042 24168
rect 2098 24112 9954 24168
rect 10010 24112 10015 24168
rect 2037 24110 10015 24112
rect 2037 24107 2103 24110
rect 9949 24107 10015 24110
rect 0 24034 480 24064
rect 4245 24034 4311 24037
rect 0 24032 4311 24034
rect 0 23976 4250 24032
rect 4306 23976 4311 24032
rect 0 23974 4311 23976
rect 0 23944 480 23974
rect 4245 23971 4311 23974
rect 20437 24034 20503 24037
rect 21909 24034 21975 24037
rect 20437 24032 21975 24034
rect 20437 23976 20442 24032
rect 20498 23976 21914 24032
rect 21970 23976 21975 24032
rect 20437 23974 21975 23976
rect 20437 23971 20503 23974
rect 21909 23971 21975 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 21541 23898 21607 23901
rect 23105 23898 23171 23901
rect 21541 23896 23171 23898
rect 21541 23840 21546 23896
rect 21602 23840 23110 23896
rect 23166 23840 23171 23896
rect 21541 23838 23171 23840
rect 21541 23835 21607 23838
rect 23105 23835 23171 23838
rect 2037 23762 2103 23765
rect 7097 23762 7163 23765
rect 2037 23760 7163 23762
rect 2037 23704 2042 23760
rect 2098 23704 7102 23760
rect 7158 23704 7163 23760
rect 2037 23702 7163 23704
rect 2037 23699 2103 23702
rect 7097 23699 7163 23702
rect 1853 23626 1919 23629
rect 7925 23626 7991 23629
rect 1853 23624 7991 23626
rect 1853 23568 1858 23624
rect 1914 23568 7930 23624
rect 7986 23568 7991 23624
rect 1853 23566 7991 23568
rect 1853 23563 1919 23566
rect 7925 23563 7991 23566
rect 8109 23626 8175 23629
rect 10685 23626 10751 23629
rect 12433 23626 12499 23629
rect 8109 23624 12499 23626
rect 8109 23568 8114 23624
rect 8170 23568 10690 23624
rect 10746 23568 12438 23624
rect 12494 23568 12499 23624
rect 8109 23566 12499 23568
rect 8109 23563 8175 23566
rect 10685 23563 10751 23566
rect 12433 23563 12499 23566
rect 17585 23626 17651 23629
rect 19149 23626 19215 23629
rect 17585 23624 19215 23626
rect 17585 23568 17590 23624
rect 17646 23568 19154 23624
rect 19210 23568 19215 23624
rect 17585 23566 19215 23568
rect 17585 23563 17651 23566
rect 19149 23563 19215 23566
rect 0 23490 480 23520
rect 2865 23490 2931 23493
rect 0 23488 2931 23490
rect 0 23432 2870 23488
rect 2926 23432 2931 23488
rect 0 23430 2931 23432
rect 0 23400 480 23430
rect 2865 23427 2931 23430
rect 7925 23490 7991 23493
rect 9397 23490 9463 23493
rect 7925 23488 9463 23490
rect 7925 23432 7930 23488
rect 7986 23432 9402 23488
rect 9458 23432 9463 23488
rect 7925 23430 9463 23432
rect 7925 23427 7991 23430
rect 9397 23427 9463 23430
rect 10869 23490 10935 23493
rect 11697 23490 11763 23493
rect 10869 23488 11763 23490
rect 10869 23432 10874 23488
rect 10930 23432 11702 23488
rect 11758 23432 11763 23488
rect 10869 23430 11763 23432
rect 10869 23427 10935 23430
rect 11697 23427 11763 23430
rect 12985 23490 13051 23493
rect 16665 23490 16731 23493
rect 12985 23488 16731 23490
rect 12985 23432 12990 23488
rect 13046 23432 16670 23488
rect 16726 23432 16731 23488
rect 12985 23430 16731 23432
rect 12985 23427 13051 23430
rect 16665 23427 16731 23430
rect 24761 23490 24827 23493
rect 26509 23490 26575 23493
rect 24761 23488 26575 23490
rect 24761 23432 24766 23488
rect 24822 23432 26514 23488
rect 26570 23432 26575 23488
rect 24761 23430 26575 23432
rect 24761 23427 24827 23430
rect 26509 23427 26575 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 15929 23354 15995 23357
rect 17401 23354 17467 23357
rect 15929 23352 17467 23354
rect 15929 23296 15934 23352
rect 15990 23296 17406 23352
rect 17462 23296 17467 23352
rect 15929 23294 17467 23296
rect 15929 23291 15995 23294
rect 17401 23291 17467 23294
rect 4521 23082 4587 23085
rect 6913 23082 6979 23085
rect 4521 23080 6979 23082
rect 4521 23024 4526 23080
rect 4582 23024 6918 23080
rect 6974 23024 6979 23080
rect 4521 23022 6979 23024
rect 4521 23019 4587 23022
rect 6913 23019 6979 23022
rect 2405 22946 2471 22949
rect 5165 22946 5231 22949
rect 2405 22944 5231 22946
rect 2405 22888 2410 22944
rect 2466 22888 5170 22944
rect 5226 22888 5231 22944
rect 2405 22886 5231 22888
rect 2405 22883 2471 22886
rect 5165 22883 5231 22886
rect 5610 22880 5930 22881
rect 0 22810 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 2773 22810 2839 22813
rect 0 22808 2839 22810
rect 0 22752 2778 22808
rect 2834 22752 2839 22808
rect 0 22750 2839 22752
rect 0 22720 480 22750
rect 2773 22747 2839 22750
rect 5533 22674 5599 22677
rect 15377 22674 15443 22677
rect 5533 22672 15443 22674
rect 5533 22616 5538 22672
rect 5594 22616 15382 22672
rect 15438 22616 15443 22672
rect 5533 22614 15443 22616
rect 5533 22611 5599 22614
rect 15377 22611 15443 22614
rect 3141 22538 3207 22541
rect 16297 22538 16363 22541
rect 3141 22536 16363 22538
rect 3141 22480 3146 22536
rect 3202 22480 16302 22536
rect 16358 22480 16363 22536
rect 3141 22478 16363 22480
rect 3141 22475 3207 22478
rect 16297 22475 16363 22478
rect 10277 22336 10597 22337
rect 0 22266 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 2957 22266 3023 22269
rect 0 22264 3023 22266
rect 0 22208 2962 22264
rect 3018 22208 3023 22264
rect 0 22206 3023 22208
rect 0 22176 480 22206
rect 2957 22203 3023 22206
rect 841 22130 907 22133
rect 4981 22130 5047 22133
rect 841 22128 5047 22130
rect 841 22072 846 22128
rect 902 22072 4986 22128
rect 5042 22072 5047 22128
rect 841 22070 5047 22072
rect 841 22067 907 22070
rect 4981 22067 5047 22070
rect 2313 21994 2379 21997
rect 9489 21994 9555 21997
rect 2313 21992 9555 21994
rect 2313 21936 2318 21992
rect 2374 21936 9494 21992
rect 9550 21936 9555 21992
rect 2313 21934 9555 21936
rect 2313 21931 2379 21934
rect 9489 21931 9555 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 1761 21722 1827 21725
rect 5441 21722 5507 21725
rect 1761 21720 5507 21722
rect 1761 21664 1766 21720
rect 1822 21664 5446 21720
rect 5502 21664 5507 21720
rect 1761 21662 5507 21664
rect 1761 21659 1827 21662
rect 5441 21659 5507 21662
rect 0 21586 480 21616
rect 3049 21586 3115 21589
rect 0 21584 3115 21586
rect 0 21528 3054 21584
rect 3110 21528 3115 21584
rect 0 21526 3115 21528
rect 0 21496 480 21526
rect 3049 21523 3115 21526
rect 3509 21586 3575 21589
rect 10041 21586 10107 21589
rect 3509 21584 10107 21586
rect 3509 21528 3514 21584
rect 3570 21528 10046 21584
rect 10102 21528 10107 21584
rect 3509 21526 10107 21528
rect 3509 21523 3575 21526
rect 10041 21523 10107 21526
rect 3417 21450 3483 21453
rect 11237 21450 11303 21453
rect 3417 21448 11303 21450
rect 3417 21392 3422 21448
rect 3478 21392 11242 21448
rect 11298 21392 11303 21448
rect 3417 21390 11303 21392
rect 3417 21387 3483 21390
rect 11237 21387 11303 21390
rect 1761 21314 1827 21317
rect 5165 21314 5231 21317
rect 1761 21312 5231 21314
rect 1761 21256 1766 21312
rect 1822 21256 5170 21312
rect 5226 21256 5231 21312
rect 1761 21254 5231 21256
rect 1761 21251 1827 21254
rect 5165 21251 5231 21254
rect 5625 21314 5691 21317
rect 6545 21314 6611 21317
rect 5625 21312 6611 21314
rect 5625 21256 5630 21312
rect 5686 21256 6550 21312
rect 6606 21256 6611 21312
rect 5625 21254 6611 21256
rect 5625 21251 5691 21254
rect 6545 21251 6611 21254
rect 10685 21314 10751 21317
rect 15285 21314 15351 21317
rect 10685 21312 15351 21314
rect 10685 21256 10690 21312
rect 10746 21256 15290 21312
rect 15346 21256 15351 21312
rect 10685 21254 15351 21256
rect 10685 21251 10751 21254
rect 15285 21251 15351 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 2405 21178 2471 21181
rect 6269 21178 6335 21181
rect 2405 21176 6335 21178
rect 2405 21120 2410 21176
rect 2466 21120 6274 21176
rect 6330 21120 6335 21176
rect 2405 21118 6335 21120
rect 2405 21115 2471 21118
rect 6269 21115 6335 21118
rect 0 21042 480 21072
rect 1393 21042 1459 21045
rect 0 21040 1459 21042
rect 0 20984 1398 21040
rect 1454 20984 1459 21040
rect 0 20982 1459 20984
rect 0 20952 480 20982
rect 1393 20979 1459 20982
rect 3693 21042 3759 21045
rect 6177 21042 6243 21045
rect 3693 21040 6243 21042
rect 3693 20984 3698 21040
rect 3754 20984 6182 21040
rect 6238 20984 6243 21040
rect 3693 20982 6243 20984
rect 3693 20979 3759 20982
rect 6177 20979 6243 20982
rect 8845 21042 8911 21045
rect 13169 21042 13235 21045
rect 8845 21040 13235 21042
rect 8845 20984 8850 21040
rect 8906 20984 13174 21040
rect 13230 20984 13235 21040
rect 8845 20982 13235 20984
rect 8845 20979 8911 20982
rect 13169 20979 13235 20982
rect 2773 20906 2839 20909
rect 5533 20906 5599 20909
rect 2773 20904 5599 20906
rect 2773 20848 2778 20904
rect 2834 20848 5538 20904
rect 5594 20848 5599 20904
rect 2773 20846 5599 20848
rect 2773 20843 2839 20846
rect 5533 20843 5599 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 5993 20634 6059 20637
rect 9029 20634 9095 20637
rect 5993 20632 9095 20634
rect 5993 20576 5998 20632
rect 6054 20576 9034 20632
rect 9090 20576 9095 20632
rect 5993 20574 9095 20576
rect 5993 20571 6059 20574
rect 9029 20571 9095 20574
rect 2313 20498 2379 20501
rect 9673 20498 9739 20501
rect 2313 20496 9739 20498
rect 2313 20440 2318 20496
rect 2374 20440 9678 20496
rect 9734 20440 9739 20496
rect 2313 20438 9739 20440
rect 2313 20435 2379 20438
rect 9673 20435 9739 20438
rect 0 20362 480 20392
rect 2773 20362 2839 20365
rect 0 20360 2839 20362
rect 0 20304 2778 20360
rect 2834 20304 2839 20360
rect 0 20302 2839 20304
rect 0 20272 480 20302
rect 2773 20299 2839 20302
rect 2681 20226 2747 20229
rect 4061 20226 4127 20229
rect 2681 20224 4127 20226
rect 2681 20168 2686 20224
rect 2742 20168 4066 20224
rect 4122 20168 4127 20224
rect 2681 20166 4127 20168
rect 2681 20163 2747 20166
rect 4061 20163 4127 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 11329 20090 11395 20093
rect 15653 20090 15719 20093
rect 11329 20088 15719 20090
rect 11329 20032 11334 20088
rect 11390 20032 15658 20088
rect 15714 20032 15719 20088
rect 11329 20030 15719 20032
rect 11329 20027 11395 20030
rect 15653 20027 15719 20030
rect 2865 19954 2931 19957
rect 1534 19952 2931 19954
rect 1534 19896 2870 19952
rect 2926 19896 2931 19952
rect 1534 19894 2931 19896
rect 0 19818 480 19848
rect 1534 19818 1594 19894
rect 2865 19891 2931 19894
rect 8385 19954 8451 19957
rect 16297 19954 16363 19957
rect 8385 19952 16363 19954
rect 8385 19896 8390 19952
rect 8446 19896 16302 19952
rect 16358 19896 16363 19952
rect 8385 19894 16363 19896
rect 8385 19891 8451 19894
rect 16297 19891 16363 19894
rect 0 19758 1594 19818
rect 2313 19818 2379 19821
rect 8017 19818 8083 19821
rect 2313 19816 8083 19818
rect 2313 19760 2318 19816
rect 2374 19760 8022 19816
rect 8078 19760 8083 19816
rect 2313 19758 8083 19760
rect 0 19728 480 19758
rect 2313 19755 2379 19758
rect 8017 19755 8083 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 4337 19410 4403 19413
rect 5533 19410 5599 19413
rect 4337 19408 5599 19410
rect 4337 19352 4342 19408
rect 4398 19352 5538 19408
rect 5594 19352 5599 19408
rect 4337 19350 5599 19352
rect 4337 19347 4403 19350
rect 5533 19347 5599 19350
rect 11881 19410 11947 19413
rect 15285 19410 15351 19413
rect 11881 19408 15351 19410
rect 11881 19352 11886 19408
rect 11942 19352 15290 19408
rect 15346 19352 15351 19408
rect 11881 19350 15351 19352
rect 11881 19347 11947 19350
rect 15285 19347 15351 19350
rect 6269 19274 6335 19277
rect 12709 19274 12775 19277
rect 6269 19272 12775 19274
rect 6269 19216 6274 19272
rect 6330 19216 12714 19272
rect 12770 19216 12775 19272
rect 6269 19214 12775 19216
rect 6269 19211 6335 19214
rect 12709 19211 12775 19214
rect 0 19138 480 19168
rect 2957 19138 3023 19141
rect 0 19136 3023 19138
rect 0 19080 2962 19136
rect 3018 19080 3023 19136
rect 0 19078 3023 19080
rect 0 19048 480 19078
rect 2957 19075 3023 19078
rect 3325 19138 3391 19141
rect 5993 19138 6059 19141
rect 3325 19136 6059 19138
rect 3325 19080 3330 19136
rect 3386 19080 5998 19136
rect 6054 19080 6059 19136
rect 3325 19078 6059 19080
rect 3325 19075 3391 19078
rect 5993 19075 6059 19078
rect 7005 19138 7071 19141
rect 8845 19138 8911 19141
rect 10133 19138 10199 19141
rect 7005 19136 10199 19138
rect 7005 19080 7010 19136
rect 7066 19080 8850 19136
rect 8906 19080 10138 19136
rect 10194 19080 10199 19136
rect 7005 19078 10199 19080
rect 7005 19075 7071 19078
rect 8845 19075 8911 19078
rect 10133 19075 10199 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 2037 19002 2103 19005
rect 4429 19002 4495 19005
rect 2037 19000 4495 19002
rect 2037 18944 2042 19000
rect 2098 18944 4434 19000
rect 4490 18944 4495 19000
rect 2037 18942 4495 18944
rect 2037 18939 2103 18942
rect 4429 18939 4495 18942
rect 6637 18866 6703 18869
rect 6913 18866 6979 18869
rect 15285 18866 15351 18869
rect 6637 18864 6979 18866
rect 6637 18808 6642 18864
rect 6698 18808 6918 18864
rect 6974 18808 6979 18864
rect 6637 18806 6979 18808
rect 6637 18803 6703 18806
rect 6913 18803 6979 18806
rect 7054 18864 15351 18866
rect 7054 18808 15290 18864
rect 15346 18808 15351 18864
rect 7054 18806 15351 18808
rect 4061 18730 4127 18733
rect 7054 18730 7114 18806
rect 15285 18803 15351 18806
rect 4061 18728 7114 18730
rect 4061 18672 4066 18728
rect 4122 18672 7114 18728
rect 4061 18670 7114 18672
rect 7281 18730 7347 18733
rect 15285 18730 15351 18733
rect 7281 18728 15351 18730
rect 7281 18672 7286 18728
rect 7342 18672 15290 18728
rect 15346 18672 15351 18728
rect 7281 18670 15351 18672
rect 4061 18667 4127 18670
rect 7281 18667 7347 18670
rect 15285 18667 15351 18670
rect 0 18594 480 18624
rect 3141 18594 3207 18597
rect 0 18592 3207 18594
rect 0 18536 3146 18592
rect 3202 18536 3207 18592
rect 0 18534 3207 18536
rect 0 18504 480 18534
rect 3141 18531 3207 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 3509 18322 3575 18325
rect 11145 18322 11211 18325
rect 3509 18320 11211 18322
rect 3509 18264 3514 18320
rect 3570 18264 11150 18320
rect 11206 18264 11211 18320
rect 3509 18262 11211 18264
rect 3509 18259 3575 18262
rect 11145 18259 11211 18262
rect 1761 18186 1827 18189
rect 4337 18186 4403 18189
rect 1761 18184 4403 18186
rect 1761 18128 1766 18184
rect 1822 18128 4342 18184
rect 4398 18128 4403 18184
rect 1761 18126 4403 18128
rect 1761 18123 1827 18126
rect 4337 18123 4403 18126
rect 10277 17984 10597 17985
rect 0 17914 480 17944
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 4521 17914 4587 17917
rect 0 17912 4587 17914
rect 0 17856 4526 17912
rect 4582 17856 4587 17912
rect 0 17854 4587 17856
rect 0 17824 480 17854
rect 4521 17851 4587 17854
rect 4797 17914 4863 17917
rect 4797 17912 10058 17914
rect 4797 17856 4802 17912
rect 4858 17856 10058 17912
rect 4797 17854 10058 17856
rect 4797 17851 4863 17854
rect 1485 17778 1551 17781
rect 2405 17778 2471 17781
rect 1485 17776 2471 17778
rect 1485 17720 1490 17776
rect 1546 17720 2410 17776
rect 2466 17720 2471 17776
rect 1485 17718 2471 17720
rect 1485 17715 1551 17718
rect 2405 17715 2471 17718
rect 3417 17778 3483 17781
rect 8477 17778 8543 17781
rect 3417 17776 8543 17778
rect 3417 17720 3422 17776
rect 3478 17720 8482 17776
rect 8538 17720 8543 17776
rect 3417 17718 8543 17720
rect 3417 17715 3483 17718
rect 8477 17715 8543 17718
rect 2129 17642 2195 17645
rect 4797 17642 4863 17645
rect 2129 17640 4863 17642
rect 2129 17584 2134 17640
rect 2190 17584 4802 17640
rect 4858 17584 4863 17640
rect 2129 17582 4863 17584
rect 2129 17579 2195 17582
rect 4797 17579 4863 17582
rect 5165 17642 5231 17645
rect 7925 17642 7991 17645
rect 5165 17640 7991 17642
rect 5165 17584 5170 17640
rect 5226 17584 7930 17640
rect 7986 17584 7991 17640
rect 5165 17582 7991 17584
rect 9998 17642 10058 17854
rect 27613 17642 27679 17645
rect 9998 17640 27679 17642
rect 9998 17584 27618 17640
rect 27674 17584 27679 17640
rect 9998 17582 27679 17584
rect 5165 17579 5231 17582
rect 7925 17579 7991 17582
rect 27613 17579 27679 17582
rect 1669 17506 1735 17509
rect 4245 17506 4311 17509
rect 1669 17504 4311 17506
rect 1669 17448 1674 17504
rect 1730 17448 4250 17504
rect 4306 17448 4311 17504
rect 1669 17446 4311 17448
rect 1669 17443 1735 17446
rect 4245 17443 4311 17446
rect 6637 17506 6703 17509
rect 7649 17506 7715 17509
rect 8293 17506 8359 17509
rect 6637 17504 8359 17506
rect 6637 17448 6642 17504
rect 6698 17448 7654 17504
rect 7710 17448 8298 17504
rect 8354 17448 8359 17504
rect 6637 17446 8359 17448
rect 6637 17443 6703 17446
rect 7649 17443 7715 17446
rect 8293 17443 8359 17446
rect 5610 17440 5930 17441
rect 0 17370 480 17400
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 3049 17370 3115 17373
rect 0 17368 3115 17370
rect 0 17312 3054 17368
rect 3110 17312 3115 17368
rect 0 17310 3115 17312
rect 0 17280 480 17310
rect 3049 17307 3115 17310
rect 3325 17234 3391 17237
rect 11145 17234 11211 17237
rect 3325 17232 11211 17234
rect 3325 17176 3330 17232
rect 3386 17176 11150 17232
rect 11206 17176 11211 17232
rect 3325 17174 11211 17176
rect 3325 17171 3391 17174
rect 11145 17171 11211 17174
rect 12985 17234 13051 17237
rect 14549 17234 14615 17237
rect 12985 17232 14615 17234
rect 12985 17176 12990 17232
rect 13046 17176 14554 17232
rect 14610 17176 14615 17232
rect 12985 17174 14615 17176
rect 12985 17171 13051 17174
rect 14549 17171 14615 17174
rect 289 17098 355 17101
rect 2313 17098 2379 17101
rect 289 17096 2379 17098
rect 289 17040 294 17096
rect 350 17040 2318 17096
rect 2374 17040 2379 17096
rect 289 17038 2379 17040
rect 289 17035 355 17038
rect 2313 17035 2379 17038
rect 2865 17098 2931 17101
rect 3601 17098 3667 17101
rect 2865 17096 3667 17098
rect 2865 17040 2870 17096
rect 2926 17040 3606 17096
rect 3662 17040 3667 17096
rect 2865 17038 3667 17040
rect 2865 17035 2931 17038
rect 3601 17035 3667 17038
rect 3785 17098 3851 17101
rect 4889 17098 4955 17101
rect 9305 17098 9371 17101
rect 3785 17096 9371 17098
rect 3785 17040 3790 17096
rect 3846 17040 4894 17096
rect 4950 17040 9310 17096
rect 9366 17040 9371 17096
rect 3785 17038 9371 17040
rect 3785 17035 3851 17038
rect 4889 17035 4955 17038
rect 9305 17035 9371 17038
rect 3141 16962 3207 16965
rect 8201 16962 8267 16965
rect 3141 16960 8267 16962
rect 3141 16904 3146 16960
rect 3202 16904 8206 16960
rect 8262 16904 8267 16960
rect 3141 16902 8267 16904
rect 3141 16899 3207 16902
rect 8201 16899 8267 16902
rect 10685 16962 10751 16965
rect 15745 16962 15811 16965
rect 10685 16960 15811 16962
rect 10685 16904 10690 16960
rect 10746 16904 15750 16960
rect 15806 16904 15811 16960
rect 10685 16902 15811 16904
rect 10685 16899 10751 16902
rect 15745 16899 15811 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 0 16690 480 16720
rect 1577 16690 1643 16693
rect 0 16688 1643 16690
rect 0 16632 1582 16688
rect 1638 16632 1643 16688
rect 0 16630 1643 16632
rect 0 16600 480 16630
rect 1577 16627 1643 16630
rect 5073 16690 5139 16693
rect 7189 16690 7255 16693
rect 5073 16688 7255 16690
rect 5073 16632 5078 16688
rect 5134 16632 7194 16688
rect 7250 16632 7255 16688
rect 5073 16630 7255 16632
rect 5073 16627 5139 16630
rect 7189 16627 7255 16630
rect 7465 16690 7531 16693
rect 13629 16690 13695 16693
rect 7465 16688 13695 16690
rect 7465 16632 7470 16688
rect 7526 16632 13634 16688
rect 13690 16632 13695 16688
rect 7465 16630 13695 16632
rect 7465 16627 7531 16630
rect 13629 16627 13695 16630
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 16146 480 16176
rect 4061 16146 4127 16149
rect 9857 16146 9923 16149
rect 0 16086 1410 16146
rect 0 16056 480 16086
rect 1350 15874 1410 16086
rect 4061 16144 9923 16146
rect 4061 16088 4066 16144
rect 4122 16088 9862 16144
rect 9918 16088 9923 16144
rect 4061 16086 9923 16088
rect 4061 16083 4127 16086
rect 9857 16083 9923 16086
rect 1485 16010 1551 16013
rect 16297 16010 16363 16013
rect 1485 16008 16363 16010
rect 1485 15952 1490 16008
rect 1546 15952 16302 16008
rect 16358 15952 16363 16008
rect 1485 15950 16363 15952
rect 1485 15947 1551 15950
rect 16297 15947 16363 15950
rect 4429 15874 4495 15877
rect 1350 15872 4495 15874
rect 1350 15816 4434 15872
rect 4490 15816 4495 15872
rect 1350 15814 4495 15816
rect 4429 15811 4495 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 3969 15602 4035 15605
rect 7925 15602 7991 15605
rect 3969 15600 7991 15602
rect 3969 15544 3974 15600
rect 4030 15544 7930 15600
rect 7986 15544 7991 15600
rect 3969 15542 7991 15544
rect 3969 15539 4035 15542
rect 7925 15539 7991 15542
rect 0 15466 480 15496
rect 5073 15466 5139 15469
rect 0 15464 5139 15466
rect 0 15408 5078 15464
rect 5134 15408 5139 15464
rect 0 15406 5139 15408
rect 0 15376 480 15406
rect 5073 15403 5139 15406
rect 6821 15466 6887 15469
rect 15285 15466 15351 15469
rect 6821 15464 15351 15466
rect 6821 15408 6826 15464
rect 6882 15408 15290 15464
rect 15346 15408 15351 15464
rect 6821 15406 15351 15408
rect 6821 15403 6887 15406
rect 15285 15403 15351 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 21817 15194 21883 15197
rect 23657 15194 23723 15197
rect 21817 15192 23723 15194
rect 21817 15136 21822 15192
rect 21878 15136 23662 15192
rect 23718 15136 23723 15192
rect 21817 15134 23723 15136
rect 21817 15131 21883 15134
rect 23657 15131 23723 15134
rect 5349 15058 5415 15061
rect 7373 15058 7439 15061
rect 5349 15056 7439 15058
rect 5349 15000 5354 15056
rect 5410 15000 7378 15056
rect 7434 15000 7439 15056
rect 5349 14998 7439 15000
rect 5349 14995 5415 14998
rect 7373 14995 7439 14998
rect 0 14922 480 14952
rect 2773 14922 2839 14925
rect 0 14920 2839 14922
rect 0 14864 2778 14920
rect 2834 14864 2839 14920
rect 0 14862 2839 14864
rect 0 14832 480 14862
rect 2773 14859 2839 14862
rect 6729 14922 6795 14925
rect 8937 14922 9003 14925
rect 9213 14922 9279 14925
rect 11329 14922 11395 14925
rect 6729 14920 11395 14922
rect 6729 14864 6734 14920
rect 6790 14864 8942 14920
rect 8998 14864 9218 14920
rect 9274 14864 11334 14920
rect 11390 14864 11395 14920
rect 6729 14862 11395 14864
rect 6729 14859 6795 14862
rect 8937 14859 9003 14862
rect 9213 14859 9279 14862
rect 11329 14859 11395 14862
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 0 14378 480 14408
rect 6545 14378 6611 14381
rect 0 14376 6611 14378
rect 0 14320 6550 14376
rect 6606 14320 6611 14376
rect 0 14318 6611 14320
rect 0 14288 480 14318
rect 6545 14315 6611 14318
rect 8569 14242 8635 14245
rect 11605 14242 11671 14245
rect 8569 14240 11671 14242
rect 8569 14184 8574 14240
rect 8630 14184 11610 14240
rect 11666 14184 11671 14240
rect 8569 14182 11671 14184
rect 8569 14179 8635 14182
rect 11605 14179 11671 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 4797 13970 4863 13973
rect 16113 13970 16179 13973
rect 4797 13968 16179 13970
rect 4797 13912 4802 13968
rect 4858 13912 16118 13968
rect 16174 13912 16179 13968
rect 4797 13910 16179 13912
rect 4797 13907 4863 13910
rect 16113 13907 16179 13910
rect 1853 13834 1919 13837
rect 1718 13832 1919 13834
rect 1718 13776 1858 13832
rect 1914 13776 1919 13832
rect 1718 13774 1919 13776
rect 0 13698 480 13728
rect 1718 13698 1778 13774
rect 1853 13771 1919 13774
rect 3325 13834 3391 13837
rect 7465 13834 7531 13837
rect 3325 13832 7531 13834
rect 3325 13776 3330 13832
rect 3386 13776 7470 13832
rect 7526 13776 7531 13832
rect 3325 13774 7531 13776
rect 3325 13771 3391 13774
rect 7465 13771 7531 13774
rect 0 13638 1778 13698
rect 6453 13698 6519 13701
rect 10133 13698 10199 13701
rect 6453 13696 10199 13698
rect 6453 13640 6458 13696
rect 6514 13640 10138 13696
rect 10194 13640 10199 13696
rect 6453 13638 10199 13640
rect 0 13608 480 13638
rect 6453 13635 6519 13638
rect 10133 13635 10199 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 6637 13426 6703 13429
rect 9765 13426 9831 13429
rect 6637 13424 9831 13426
rect 6637 13368 6642 13424
rect 6698 13368 9770 13424
rect 9826 13368 9831 13424
rect 6637 13366 9831 13368
rect 6637 13363 6703 13366
rect 9765 13363 9831 13366
rect 8017 13290 8083 13293
rect 20713 13290 20779 13293
rect 8017 13288 20779 13290
rect 8017 13232 8022 13288
rect 8078 13232 20718 13288
rect 20774 13232 20779 13288
rect 8017 13230 20779 13232
rect 8017 13227 8083 13230
rect 20713 13227 20779 13230
rect 0 13154 480 13184
rect 1669 13154 1735 13157
rect 0 13152 1735 13154
rect 0 13096 1674 13152
rect 1730 13096 1735 13152
rect 0 13094 1735 13096
rect 0 13064 480 13094
rect 1669 13091 1735 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 2129 13018 2195 13021
rect 2129 13016 5458 13018
rect 2129 12960 2134 13016
rect 2190 12960 5458 13016
rect 2129 12958 5458 12960
rect 2129 12955 2195 12958
rect 5398 12885 5458 12958
rect 2681 12882 2747 12885
rect 5257 12882 5323 12885
rect 2681 12880 5323 12882
rect 2681 12824 2686 12880
rect 2742 12824 5262 12880
rect 5318 12824 5323 12880
rect 2681 12822 5323 12824
rect 5398 12882 5507 12885
rect 7465 12882 7531 12885
rect 5398 12880 7531 12882
rect 5398 12824 5446 12880
rect 5502 12824 7470 12880
rect 7526 12824 7531 12880
rect 5398 12822 7531 12824
rect 2681 12819 2747 12822
rect 5257 12819 5323 12822
rect 5441 12819 5507 12822
rect 7465 12819 7531 12822
rect 10409 12882 10475 12885
rect 16757 12882 16823 12885
rect 10409 12880 16823 12882
rect 10409 12824 10414 12880
rect 10470 12824 16762 12880
rect 16818 12824 16823 12880
rect 10409 12822 16823 12824
rect 10409 12819 10475 12822
rect 16757 12819 16823 12822
rect 16941 12882 17007 12885
rect 18597 12882 18663 12885
rect 16941 12880 18663 12882
rect 16941 12824 16946 12880
rect 17002 12824 18602 12880
rect 18658 12824 18663 12880
rect 16941 12822 18663 12824
rect 16941 12819 17007 12822
rect 18597 12819 18663 12822
rect 3969 12746 4035 12749
rect 11513 12746 11579 12749
rect 12157 12746 12223 12749
rect 3969 12744 12223 12746
rect 3969 12688 3974 12744
rect 4030 12688 11518 12744
rect 11574 12688 12162 12744
rect 12218 12688 12223 12744
rect 3969 12686 12223 12688
rect 3969 12683 4035 12686
rect 11513 12683 11579 12686
rect 12157 12683 12223 12686
rect 13261 12746 13327 12749
rect 18045 12746 18111 12749
rect 13261 12744 18111 12746
rect 13261 12688 13266 12744
rect 13322 12688 18050 12744
rect 18106 12688 18111 12744
rect 13261 12686 18111 12688
rect 13261 12683 13327 12686
rect 18045 12683 18111 12686
rect 10277 12544 10597 12545
rect 0 12474 480 12504
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 4061 12474 4127 12477
rect 0 12472 4127 12474
rect 0 12416 4066 12472
rect 4122 12416 4127 12472
rect 0 12414 4127 12416
rect 0 12384 480 12414
rect 4061 12411 4127 12414
rect 6545 12338 6611 12341
rect 8293 12338 8359 12341
rect 6545 12336 8359 12338
rect 6545 12280 6550 12336
rect 6606 12280 8298 12336
rect 8354 12280 8359 12336
rect 6545 12278 8359 12280
rect 6545 12275 6611 12278
rect 8293 12275 8359 12278
rect 1761 12202 1827 12205
rect 13997 12202 14063 12205
rect 1761 12200 14063 12202
rect 1761 12144 1766 12200
rect 1822 12144 14002 12200
rect 14058 12144 14063 12200
rect 1761 12142 14063 12144
rect 1761 12139 1827 12142
rect 13997 12139 14063 12142
rect 7005 12066 7071 12069
rect 8753 12066 8819 12069
rect 7005 12064 8819 12066
rect 7005 12008 7010 12064
rect 7066 12008 8758 12064
rect 8814 12008 8819 12064
rect 7005 12006 8819 12008
rect 7005 12003 7071 12006
rect 8753 12003 8819 12006
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 0 11870 3618 11930
rect 0 11840 480 11870
rect 3558 11386 3618 11870
rect 3877 11794 3943 11797
rect 5993 11794 6059 11797
rect 3877 11792 6059 11794
rect 3877 11736 3882 11792
rect 3938 11736 5998 11792
rect 6054 11736 6059 11792
rect 3877 11734 6059 11736
rect 3877 11731 3943 11734
rect 5993 11731 6059 11734
rect 3693 11522 3759 11525
rect 6545 11522 6611 11525
rect 3693 11520 6611 11522
rect 3693 11464 3698 11520
rect 3754 11464 6550 11520
rect 6606 11464 6611 11520
rect 3693 11462 6611 11464
rect 3693 11459 3759 11462
rect 6545 11459 6611 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 10133 11386 10199 11389
rect 3558 11384 10199 11386
rect 3558 11328 10138 11384
rect 10194 11328 10199 11384
rect 3558 11326 10199 11328
rect 10133 11323 10199 11326
rect 0 11250 480 11280
rect 3509 11250 3575 11253
rect 0 11248 3575 11250
rect 0 11192 3514 11248
rect 3570 11192 3575 11248
rect 0 11190 3575 11192
rect 0 11160 480 11190
rect 3509 11187 3575 11190
rect 10869 11250 10935 11253
rect 14089 11250 14155 11253
rect 10869 11248 14155 11250
rect 10869 11192 10874 11248
rect 10930 11192 14094 11248
rect 14150 11192 14155 11248
rect 10869 11190 14155 11192
rect 10869 11187 10935 11190
rect 14089 11187 14155 11190
rect 18781 11250 18847 11253
rect 19425 11250 19491 11253
rect 18781 11248 19491 11250
rect 18781 11192 18786 11248
rect 18842 11192 19430 11248
rect 19486 11192 19491 11248
rect 18781 11190 19491 11192
rect 18781 11187 18847 11190
rect 19425 11187 19491 11190
rect 10225 11114 10291 11117
rect 18505 11114 18571 11117
rect 10225 11112 18571 11114
rect 10225 11056 10230 11112
rect 10286 11056 18510 11112
rect 18566 11056 18571 11112
rect 10225 11054 18571 11056
rect 10225 11051 10291 11054
rect 18505 11051 18571 11054
rect 12709 10978 12775 10981
rect 6134 10976 12775 10978
rect 6134 10920 12714 10976
rect 12770 10920 12775 10976
rect 6134 10918 12775 10920
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 2497 10842 2563 10845
rect 2497 10840 5458 10842
rect 2497 10784 2502 10840
rect 2558 10784 5458 10840
rect 2497 10782 5458 10784
rect 2497 10779 2563 10782
rect 0 10706 480 10736
rect 5398 10706 5458 10782
rect 6134 10706 6194 10918
rect 12709 10915 12775 10918
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 0 10646 3434 10706
rect 5398 10646 6194 10706
rect 7465 10706 7531 10709
rect 20161 10706 20227 10709
rect 7465 10704 20227 10706
rect 7465 10648 7470 10704
rect 7526 10648 20166 10704
rect 20222 10648 20227 10704
rect 7465 10646 20227 10648
rect 0 10616 480 10646
rect 3374 10434 3434 10646
rect 7465 10643 7531 10646
rect 20161 10643 20227 10646
rect 3509 10570 3575 10573
rect 12157 10570 12223 10573
rect 3509 10568 12223 10570
rect 3509 10512 3514 10568
rect 3570 10512 12162 10568
rect 12218 10512 12223 10568
rect 3509 10510 12223 10512
rect 3509 10507 3575 10510
rect 12157 10507 12223 10510
rect 9949 10434 10015 10437
rect 3374 10432 10015 10434
rect 3374 10376 9954 10432
rect 10010 10376 10015 10432
rect 3374 10374 10015 10376
rect 9949 10371 10015 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 1761 10298 1827 10301
rect 2589 10298 2655 10301
rect 7741 10298 7807 10301
rect 1761 10296 7807 10298
rect 1761 10240 1766 10296
rect 1822 10240 2594 10296
rect 2650 10240 7746 10296
rect 7802 10240 7807 10296
rect 1761 10238 7807 10240
rect 1761 10235 1827 10238
rect 2589 10235 2655 10238
rect 7741 10235 7807 10238
rect 5625 10162 5691 10165
rect 16665 10162 16731 10165
rect 5625 10160 16731 10162
rect 5625 10104 5630 10160
rect 5686 10104 16670 10160
rect 16726 10104 16731 10160
rect 5625 10102 16731 10104
rect 5625 10099 5691 10102
rect 16665 10099 16731 10102
rect 19149 10162 19215 10165
rect 20253 10162 20319 10165
rect 19149 10160 20319 10162
rect 19149 10104 19154 10160
rect 19210 10104 20258 10160
rect 20314 10104 20319 10160
rect 19149 10102 20319 10104
rect 19149 10099 19215 10102
rect 20253 10099 20319 10102
rect 0 10026 480 10056
rect 2957 10026 3023 10029
rect 0 10024 3023 10026
rect 0 9968 2962 10024
rect 3018 9968 3023 10024
rect 0 9966 3023 9968
rect 0 9936 480 9966
rect 2957 9963 3023 9966
rect 4061 10026 4127 10029
rect 18873 10026 18939 10029
rect 4061 10024 18939 10026
rect 4061 9968 4066 10024
rect 4122 9968 18878 10024
rect 18934 9968 18939 10024
rect 4061 9966 18939 9968
rect 4061 9963 4127 9966
rect 18873 9963 18939 9966
rect 6821 9890 6887 9893
rect 8477 9890 8543 9893
rect 6821 9888 8543 9890
rect 6821 9832 6826 9888
rect 6882 9832 8482 9888
rect 8538 9832 8543 9888
rect 6821 9830 8543 9832
rect 6821 9827 6887 9830
rect 8477 9827 8543 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 0 9482 480 9512
rect 4889 9482 4955 9485
rect 0 9480 4955 9482
rect 0 9424 4894 9480
rect 4950 9424 4955 9480
rect 0 9422 4955 9424
rect 0 9392 480 9422
rect 4889 9419 4955 9422
rect 5073 9482 5139 9485
rect 11881 9482 11947 9485
rect 5073 9480 11947 9482
rect 5073 9424 5078 9480
rect 5134 9424 11886 9480
rect 11942 9424 11947 9480
rect 5073 9422 11947 9424
rect 5073 9419 5139 9422
rect 11881 9419 11947 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 2681 9074 2747 9077
rect 3417 9074 3483 9077
rect 6637 9074 6703 9077
rect 2681 9072 6703 9074
rect 2681 9016 2686 9072
rect 2742 9016 3422 9072
rect 3478 9016 6642 9072
rect 6698 9016 6703 9072
rect 2681 9014 6703 9016
rect 2681 9011 2747 9014
rect 3417 9011 3483 9014
rect 6637 9011 6703 9014
rect 8293 8938 8359 8941
rect 3374 8936 8359 8938
rect 3374 8880 8298 8936
rect 8354 8880 8359 8936
rect 3374 8878 8359 8880
rect 0 8802 480 8832
rect 3374 8802 3434 8878
rect 8293 8875 8359 8878
rect 0 8742 3434 8802
rect 0 8712 480 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 6821 8394 6887 8397
rect 19333 8394 19399 8397
rect 6821 8392 19480 8394
rect 6821 8336 6826 8392
rect 6882 8336 19338 8392
rect 19394 8336 19480 8392
rect 6821 8334 19480 8336
rect 6821 8331 6887 8334
rect 19333 8331 19399 8334
rect 0 8258 480 8288
rect 3693 8258 3759 8261
rect 0 8256 3759 8258
rect 0 8200 3698 8256
rect 3754 8200 3759 8256
rect 0 8198 3759 8200
rect 0 8168 480 8198
rect 3693 8195 3759 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 5610 7648 5930 7649
rect 0 7578 480 7608
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 0 7518 3434 7578
rect 0 7488 480 7518
rect 3374 7306 3434 7518
rect 22277 7306 22343 7309
rect 3374 7304 22343 7306
rect 3374 7248 22282 7304
rect 22338 7248 22343 7304
rect 3374 7246 22343 7248
rect 22277 7243 22343 7246
rect 10277 7104 10597 7105
rect 0 7034 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 0 6974 3986 7034
rect 0 6944 480 6974
rect 3926 6898 3986 6974
rect 22737 6898 22803 6901
rect 3926 6896 22803 6898
rect 3926 6840 22742 6896
rect 22798 6840 22803 6896
rect 3926 6838 22803 6840
rect 22737 6835 22803 6838
rect 23841 6898 23907 6901
rect 24945 6898 25011 6901
rect 23841 6896 25011 6898
rect 23841 6840 23846 6896
rect 23902 6840 24950 6896
rect 25006 6840 25011 6896
rect 23841 6838 25011 6840
rect 23841 6835 23907 6838
rect 24945 6835 25011 6838
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 0 6354 480 6384
rect 0 6294 674 6354
rect 0 6264 480 6294
rect 614 6218 674 6294
rect 23657 6218 23723 6221
rect 614 6216 23723 6218
rect 614 6160 23662 6216
rect 23718 6160 23723 6216
rect 614 6158 23723 6160
rect 23657 6155 23723 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 0 5810 480 5840
rect 24025 5810 24091 5813
rect 0 5808 24091 5810
rect 0 5752 24030 5808
rect 24086 5752 24091 5808
rect 0 5750 24091 5752
rect 0 5720 480 5750
rect 24025 5747 24091 5750
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 24577 5266 24643 5269
rect 614 5264 24643 5266
rect 614 5208 24582 5264
rect 24638 5208 24643 5264
rect 614 5206 24643 5208
rect 0 5130 480 5160
rect 614 5130 674 5206
rect 24577 5203 24643 5206
rect 0 5070 674 5130
rect 0 5040 480 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 24761 4858 24827 4861
rect 26233 4858 26299 4861
rect 24761 4856 26299 4858
rect 24761 4800 24766 4856
rect 24822 4800 26238 4856
rect 26294 4800 26299 4856
rect 24761 4798 26299 4800
rect 24761 4795 24827 4798
rect 26233 4795 26299 4798
rect 0 4586 480 4616
rect 0 4526 674 4586
rect 0 4496 480 4526
rect 614 4178 674 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 24577 4178 24643 4181
rect 614 4176 24643 4178
rect 614 4120 24582 4176
rect 24638 4120 24643 4176
rect 614 4118 24643 4120
rect 24577 4115 24643 4118
rect 4613 4042 4679 4045
rect 8385 4042 8451 4045
rect 4613 4040 8451 4042
rect 4613 3984 4618 4040
rect 4674 3984 8390 4040
rect 8446 3984 8451 4040
rect 4613 3982 8451 3984
rect 4613 3979 4679 3982
rect 8385 3979 8451 3982
rect 0 3906 480 3936
rect 2037 3906 2103 3909
rect 0 3904 2103 3906
rect 0 3848 2042 3904
rect 2098 3848 2103 3904
rect 0 3846 2103 3848
rect 0 3816 480 3846
rect 2037 3843 2103 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 6177 3498 6243 3501
rect 23197 3498 23263 3501
rect 6177 3496 23263 3498
rect 6177 3440 6182 3496
rect 6238 3440 23202 3496
rect 23258 3440 23263 3496
rect 6177 3438 23263 3440
rect 6177 3435 6243 3438
rect 23197 3435 23263 3438
rect 0 3362 480 3392
rect 3969 3362 4035 3365
rect 0 3360 4035 3362
rect 0 3304 3974 3360
rect 4030 3304 4035 3360
rect 0 3302 4035 3304
rect 0 3272 480 3302
rect 3969 3299 4035 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 2589 2954 2655 2957
rect 13905 2954 13971 2957
rect 2589 2952 13971 2954
rect 2589 2896 2594 2952
rect 2650 2896 13910 2952
rect 13966 2896 13971 2952
rect 2589 2894 13971 2896
rect 2589 2891 2655 2894
rect 13905 2891 13971 2894
rect 10277 2752 10597 2753
rect 0 2682 480 2712
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 3785 2682 3851 2685
rect 0 2680 3851 2682
rect 0 2624 3790 2680
rect 3846 2624 3851 2680
rect 0 2622 3851 2624
rect 0 2592 480 2622
rect 3785 2619 3851 2622
rect 5610 2208 5930 2209
rect 0 2138 480 2168
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 4337 2138 4403 2141
rect 0 2136 4403 2138
rect 0 2080 4342 2136
rect 4398 2080 4403 2136
rect 0 2078 4403 2080
rect 0 2048 480 2078
rect 4337 2075 4403 2078
rect 0 1458 480 1488
rect 9305 1458 9371 1461
rect 0 1456 9371 1458
rect 0 1400 9310 1456
rect 9366 1400 9371 1456
rect 0 1398 9371 1400
rect 0 1368 480 1398
rect 9305 1395 9371 1398
rect 12617 1322 12683 1325
rect 614 1320 12683 1322
rect 614 1264 12622 1320
rect 12678 1264 12683 1320
rect 614 1262 12683 1264
rect 0 914 480 944
rect 614 914 674 1262
rect 12617 1259 12683 1262
rect 0 854 674 914
rect 0 824 480 854
rect 0 370 480 400
rect 3325 370 3391 373
rect 0 368 3391 370
rect 0 312 3330 368
rect 3386 312 3391 368
rect 0 310 3391 312
rect 0 280 480 310
rect 3325 307 3391 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2300 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1604681595
transform 1 0 4048 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1604681595
transform 1 0 5152 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_56
timestamp 1604681595
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604681595
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604681595
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604681595
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1604681595
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_273
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604681595
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604681595
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1604681595
transform 1 0 24564 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_253
timestamp 1604681595
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _80_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24564 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_251
timestamp 1604681595
transform 1 0 24196 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_259
timestamp 1604681595
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1604681595
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604681595
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1604681595
transform 1 0 24012 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1604681595
transform 1 0 24564 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1604681595
transform 1 0 25116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_251
timestamp 1604681595
transform 1 0 24196 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_259
timestamp 1604681595
transform 1 0 24932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_263
timestamp 1604681595
transform 1 0 25300 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_275
timestamp 1604681595
transform 1 0 26404 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604681595
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604681595
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_237
timestamp 1604681595
transform 1 0 22908 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_232
timestamp 1604681595
transform 1 0 22448 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1604681595
transform 1 0 22724 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1604681595
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_249
timestamp 1604681595
transform 1 0 24012 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_247
timestamp 1604681595
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1604681595
transform 1 0 24012 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1604681595
transform 1 0 24196 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1604681595
transform 1 0 24380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1604681595
transform 1 0 25484 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_253
timestamp 1604681595
transform 1 0 24380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_265
timestamp 1604681595
transform 1 0 25484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp 1604681595
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1604681595
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_227
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1604681595
transform 1 0 22724 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1604681595
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1604681595
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1604681595
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_35
timestamp 1604681595
transform 1 0 4324 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_38
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _41_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5612 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_46
timestamp 1604681595
transform 1 0 5336 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_55
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8096 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_65
timestamp 1604681595
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_69
timestamp 1604681595
transform 1 0 7452 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_75
timestamp 1604681595
transform 1 0 8004 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1604681595
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_83
timestamp 1604681595
transform 1 0 8740 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_95
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_107
timestamp 1604681595
transform 1 0 10948 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp 1604681595
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1604681595
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_228
timestamp 1604681595
transform 1 0 22080 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1604681595
transform 1 0 22264 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1604681595
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_234
timestamp 1604681595
transform 1 0 22632 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_238
timestamp 1604681595
transform 1 0 23000 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 1564 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_8
timestamp 1604681595
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_12
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_16
timestamp 1604681595
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_20
timestamp 1604681595
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_24
timestamp 1604681595
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_28
timestamp 1604681595
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_36
timestamp 1604681595
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1604681595
transform 1 0 4140 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_40
timestamp 1604681595
transform 1 0 4784 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5612 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_45
timestamp 1604681595
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1604681595
transform 1 0 8096 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_72
timestamp 1604681595
transform 1 0 7728 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_79
timestamp 1604681595
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_83
timestamp 1604681595
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1604681595
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1604681595
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1564 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_14
timestamp 1604681595
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_18
timestamp 1604681595
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3128 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_31
timestamp 1604681595
transform 1 0 3956 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_35
timestamp 1604681595
transform 1 0 4324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_38
timestamp 1604681595
transform 1 0 4600 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5060 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_52
timestamp 1604681595
transform 1 0 5888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1604681595
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_75
timestamp 1604681595
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_88
timestamp 1604681595
transform 1 0 9200 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_100
timestamp 1604681595
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_104
timestamp 1604681595
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_108
timestamp 1604681595
transform 1 0 11040 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1604681595
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 1564 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_14
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_18
timestamp 1604681595
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4416 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_22
timestamp 1604681595
transform 1 0 3128 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_28
timestamp 1604681595
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_55
timestamp 1604681595
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1604681595
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6900 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_12_82
timestamp 1604681595
transform 1 0 8648 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1604681595
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_101
timestamp 1604681595
transform 1 0 10396 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1604681595
transform 1 0 12236 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_133
timestamp 1604681595
transform 1 0 13340 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1564 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2208 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_9
timestamp 1604681595
transform 1 0 1932 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_25
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_21
timestamp 1604681595
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_28
timestamp 1604681595
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_24
timestamp 1604681595
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4048 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_45
timestamp 1604681595
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5612 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_58
timestamp 1604681595
transform 1 0 6440 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_55
timestamp 1604681595
transform 1 0 6164 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1604681595
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_69
timestamp 1604681595
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_66
timestamp 1604681595
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_76
timestamp 1604681595
transform 1 0 8096 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7636 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1604681595
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1604681595
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_104
timestamp 1604681595
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_100
timestamp 1604681595
transform 1 0 10304 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_94
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604681595
transform 1 0 10396 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10120 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_108
timestamp 1604681595
transform 1 0 11040 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_117
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_125
timestamp 1604681595
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_129
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_133
timestamp 1604681595
transform 1 0 13340 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1604681595
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1604681595
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1604681595
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_195
timestamp 1604681595
transform 1 0 19044 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_192
timestamp 1604681595
transform 1 0 18768 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18860 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_204
timestamp 1604681595
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19320 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_199
timestamp 1604681595
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1604681595
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604681595
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1840 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4324 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_31
timestamp 1604681595
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_44
timestamp 1604681595
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1604681595
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_52
timestamp 1604681595
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5704 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_56
timestamp 1604681595
transform 1 0 6256 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_67
timestamp 1604681595
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1604681595
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_94
timestamp 1604681595
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_107
timestamp 1604681595
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_111
timestamp 1604681595
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1604681595
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1604681595
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_136
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_148
timestamp 1604681595
transform 1 0 14720 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_160
timestamp 1604681595
transform 1 0 15824 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_172
timestamp 1604681595
transform 1 0 16928 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1604681595
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20148 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18492 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_188
timestamp 1604681595
transform 1 0 18400 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_191
timestamp 1604681595
transform 1 0 18676 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_203
timestamp 1604681595
transform 1 0 19780 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_213
timestamp 1604681595
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_217
timestamp 1604681595
transform 1 0 21068 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_229
timestamp 1604681595
transform 1 0 22172 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_241
timestamp 1604681595
transform 1 0 23276 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_16
timestamp 1604681595
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_20
timestamp 1604681595
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_24
timestamp 1604681595
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_28
timestamp 1604681595
transform 1 0 3680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4324 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_37
timestamp 1604681595
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4692 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4968 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_16_61
timestamp 1604681595
transform 1 0 6716 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7452 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_66
timestamp 1604681595
transform 1 0 7176 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_78
timestamp 1604681595
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1604681595
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10212 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 9016 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_89
timestamp 1604681595
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11224 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11592 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_108
timestamp 1604681595
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_112
timestamp 1604681595
transform 1 0 11408 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_116
timestamp 1604681595
transform 1 0 11776 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_120
timestamp 1604681595
transform 1 0 12144 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_125
timestamp 1604681595
transform 1 0 12604 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12696 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_178
timestamp 1604681595
transform 1 0 17480 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_186
timestamp 1604681595
transform 1 0 18216 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18492 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_195
timestamp 1604681595
transform 1 0 19044 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_207
timestamp 1604681595
transform 1 0 20148 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604681595
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1656 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_19
timestamp 1604681595
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 3680 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_23
timestamp 1604681595
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_50
timestamp 1604681595
transform 1 0 5704 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_54
timestamp 1604681595
transform 1 0 6072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1604681595
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9292 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_85
timestamp 1604681595
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_108
timestamp 1604681595
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_112
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_142
timestamp 1604681595
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 14904 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_146
timestamp 1604681595
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_153
timestamp 1604681595
transform 1 0 15180 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_165
timestamp 1604681595
transform 1 0 16284 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_177
timestamp 1604681595
transform 1 0 17388 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1604681595
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_232
timestamp 1604681595
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_16
timestamp 1604681595
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1604681595
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3496 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_24
timestamp 1604681595
transform 1 0 3312 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_28
timestamp 1604681595
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_51
timestamp 1604681595
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_55
timestamp 1604681595
transform 1 0 6164 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp 1604681595
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_26.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7820 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6992 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 9752 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1604681595
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_101
timestamp 1604681595
transform 1 0 10396 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_18_124
timestamp 1604681595
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13248 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_128
timestamp 1604681595
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1604681595
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1604681595
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1604681595
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1604681595
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1604681595
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1604681595
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_8
timestamp 1604681595
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1656 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_19
timestamp 1604681595
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_12
timestamp 1604681595
transform 1 0 2208 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2300 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1604681595
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_32
timestamp 1604681595
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_35
timestamp 1604681595
transform 1 0 4324 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1604681595
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_39
timestamp 1604681595
transform 1 0 4692 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4784 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_42
timestamp 1604681595
transform 1 0 4968 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_49
timestamp 1604681595
transform 1 0 5612 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5244 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1604681595
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_54
timestamp 1604681595
transform 1 0 6072 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_71
timestamp 1604681595
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_67
timestamp 1604681595
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_72
timestamp 1604681595
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_69
timestamp 1604681595
transform 1 0 7452 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_65
timestamp 1604681595
transform 1 0 7084 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1604681595
transform 1 0 6992 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 8096 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_98
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_114
timestamp 1604681595
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_106
timestamp 1604681595
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_122
timestamp 1604681595
transform 1 0 12328 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_118
timestamp 1604681595
transform 1 0 11960 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13984 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1604681595
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_136
timestamp 1604681595
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_132
timestamp 1604681595
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_136
timestamp 1604681595
transform 1 0 13616 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1604681595
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1604681595
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_150
timestamp 1604681595
transform 1 0 14904 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_146
timestamp 1604681595
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _99_
timestamp 1604681595
transform 1 0 15272 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_166
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1604681595
transform 1 0 16008 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_158
timestamp 1604681595
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__99__A
timestamp 1604681595
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_174
timestamp 1604681595
transform 1 0 17112 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_168
timestamp 1604681595
transform 1 0 16560 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17388 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_183
timestamp 1604681595
transform 1 0 17940 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18768 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_190
timestamp 1604681595
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_194
timestamp 1604681595
transform 1 0 18952 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_206
timestamp 1604681595
transform 1 0 20056 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_195
timestamp 1604681595
transform 1 0 19044 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_207
timestamp 1604681595
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_218
timestamp 1604681595
transform 1 0 21160 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604681595
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_230
timestamp 1604681595
transform 1 0 22264 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_242
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1604681595
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_251
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_263
timestamp 1604681595
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 1656 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1604681595
transform 1 0 4140 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_25
timestamp 1604681595
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1604681595
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_36
timestamp 1604681595
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8372 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_75
timestamp 1604681595
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1604681595
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_103
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1604681595
transform 1 0 10856 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_109
timestamp 1604681595
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1604681595
transform 1 0 11500 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_142
timestamp 1604681595
transform 1 0 14168 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16100 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_154
timestamp 1604681595
transform 1 0 15272 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_162
timestamp 1604681595
transform 1 0 16008 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1604681595
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_173
timestamp 1604681595
transform 1 0 17020 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20700 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_212
timestamp 1604681595
transform 1 0 20608 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_219
timestamp 1604681595
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_223
timestamp 1604681595
transform 1 0 21620 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_235
timestamp 1604681595
transform 1 0 22724 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_243
timestamp 1604681595
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1604681595
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1604681595
transform 1 0 2944 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_12
timestamp 1604681595
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_16
timestamp 1604681595
transform 1 0 2576 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_36
timestamp 1604681595
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_40
timestamp 1604681595
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_63
timestamp 1604681595
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_67
timestamp 1604681595
transform 1 0 7268 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_72
timestamp 1604681595
transform 1 0 7728 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10212 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1604681595
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_97
timestamp 1604681595
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_118
timestamp 1604681595
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_122
timestamp 1604681595
transform 1 0 12328 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12696 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1604681595
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1472 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4232 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1604681595
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_31
timestamp 1604681595
transform 1 0 3956 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7544 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_66
timestamp 1604681595
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_79
timestamp 1604681595
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_83
timestamp 1604681595
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9108 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_106
timestamp 1604681595
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1604681595
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1604681595
transform 1 0 12512 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_127
timestamp 1604681595
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1604681595
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_154
timestamp 1604681595
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_158
timestamp 1604681595
transform 1 0 15640 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_170
timestamp 1604681595
transform 1 0 16744 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1604681595
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1604681595
transform 1 0 21620 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1604681595
transform 1 0 22172 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_227
timestamp 1604681595
transform 1 0 21988 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_231
timestamp 1604681595
transform 1 0 22356 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_243
timestamp 1604681595
transform 1 0 23460 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2024 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1604681595
transform 1 0 1748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1604681595
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_40
timestamp 1604681595
transform 1 0 4784 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_36
timestamp 1604681595
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5244 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7728 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_64
timestamp 1604681595
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_78
timestamp 1604681595
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1604681595
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_86
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_102
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 11316 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12328 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_106
timestamp 1604681595
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_110
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_120
timestamp 1604681595
transform 1 0 12144 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_124
timestamp 1604681595
transform 1 0 12512 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13892 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_137
timestamp 1604681595
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_145
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1604681595
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_160
timestamp 1604681595
transform 1 0 15824 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_172
timestamp 1604681595
transform 1 0 16928 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_184
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_196
timestamp 1604681595
transform 1 0 19136 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_208
timestamp 1604681595
transform 1 0 20240 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604681595
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1472 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_13
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_17
timestamp 1604681595
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3036 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_25_40
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 5520 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_45
timestamp 1604681595
transform 1 0 5244 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_71
timestamp 1604681595
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_75
timestamp 1604681595
transform 1 0 8004 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_80
timestamp 1604681595
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8832 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1604681595
transform 1 0 9660 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_97
timestamp 1604681595
transform 1 0 10028 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1604681595
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1604681595
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1604681595
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13892 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_127
timestamp 1604681595
transform 1 0 12788 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_130
timestamp 1604681595
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_134
timestamp 1604681595
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_138
timestamp 1604681595
transform 1 0 13800 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16376 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_158
timestamp 1604681595
transform 1 0 15640 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1604681595
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_176
timestamp 1604681595
transform 1 0 17296 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1604681595
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1604681595
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1604681595
transform 1 0 1748 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 1840 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_17
timestamp 1604681595
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2300 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2852 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_25
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_21
timestamp 1604681595
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_28
timestamp 1604681595
transform 1 0 3680 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_34
timestamp 1604681595
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_35
timestamp 1604681595
transform 1 0 4324 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1604681595
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_39
timestamp 1604681595
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_42
timestamp 1604681595
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_52
timestamp 1604681595
transform 1 0 5888 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5060 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1604681595
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_53
timestamp 1604681595
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1604681595
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6072 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6624 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8280 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 8004 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_69
timestamp 1604681595
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_73
timestamp 1604681595
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_77
timestamp 1604681595
transform 1 0 8188 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_81
timestamp 1604681595
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_85
timestamp 1604681595
transform 1 0 8924 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_88
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_84
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9384 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_103
timestamp 1604681595
transform 1 0 10580 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1604681595
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1604681595
transform 1 0 10028 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10120 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_109
timestamp 1604681595
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_111
timestamp 1604681595
transform 1 0 11316 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_107
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 11500 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_118
timestamp 1604681595
transform 1 0 11960 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 11684 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12512 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_133
timestamp 1604681595
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_132
timestamp 1604681595
transform 1 0 13248 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_128
timestamp 1604681595
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_137
timestamp 1604681595
transform 1 0 13708 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14352 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_163
timestamp 1604681595
transform 1 0 16100 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604681595
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1604681595
transform 1 0 17204 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1604681595
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604681595
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1604681595
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1472 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1604681595
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5980 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 5612 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_45
timestamp 1604681595
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_52
timestamp 1604681595
transform 1 0 5888 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 8556 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8280 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_72
timestamp 1604681595
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_76
timestamp 1604681595
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12144 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11592 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_112
timestamp 1604681595
transform 1 0 11408 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_116
timestamp 1604681595
transform 1 0 11776 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_139
timestamp 1604681595
transform 1 0 13892 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_143
timestamp 1604681595
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_146
timestamp 1604681595
transform 1 0 14536 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1604681595
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4232 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_26
timestamp 1604681595
transform 1 0 3496 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_30
timestamp 1604681595
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_71
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_75
timestamp 1604681595
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_79
timestamp 1604681595
transform 1 0 8372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9200 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_84
timestamp 1604681595
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_97
timestamp 1604681595
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1604681595
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_142
timestamp 1604681595
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15364 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16100 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_146
timestamp 1604681595
transform 1 0 14536 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_152
timestamp 1604681595
transform 1 0 15088 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_161
timestamp 1604681595
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_165
timestamp 1604681595
transform 1 0 16284 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_177
timestamp 1604681595
transform 1 0 17388 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_6
timestamp 1604681595
transform 1 0 1656 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1604681595
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_41
timestamp 1604681595
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5704 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_45
timestamp 1604681595
transform 1 0 5244 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_59
timestamp 1604681595
transform 1 0 6532 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8280 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8648 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_64
timestamp 1604681595
transform 1 0 6992 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_76
timestamp 1604681595
transform 1 0 8096 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_84
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_99
timestamp 1604681595
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_103
timestamp 1604681595
transform 1 0 10580 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12512 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10948 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_116
timestamp 1604681595
transform 1 0 11776 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_120
timestamp 1604681595
transform 1 0 12144 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_143
timestamp 1604681595
transform 1 0 14260 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16008 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1604681595
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_160
timestamp 1604681595
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_164
timestamp 1604681595
transform 1 0 16192 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_176
timestamp 1604681595
transform 1 0 17296 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_188
timestamp 1604681595
transform 1 0 18400 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_200
timestamp 1604681595
transform 1 0 19504 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2024 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_19
timestamp 1604681595
transform 1 0 2852 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3128 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_24
timestamp 1604681595
transform 1 0 3312 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_28
timestamp 1604681595
transform 1 0 3680 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_41
timestamp 1604681595
transform 1 0 4876 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_45
timestamp 1604681595
transform 1 0 5244 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5060 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5428 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 5612 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_53
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7728 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_65
timestamp 1604681595
transform 1 0 7084 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_70
timestamp 1604681595
transform 1 0 7544 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_93
timestamp 1604681595
transform 1 0 9660 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_99
timestamp 1604681595
transform 1 0 10212 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 10764 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604681595
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13248 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_128
timestamp 1604681595
transform 1 0 12880 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _97_
timestamp 1604681595
transform 1 0 15732 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16284 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_151
timestamp 1604681595
transform 1 0 14996 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_156
timestamp 1604681595
transform 1 0 15456 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_163
timestamp 1604681595
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__97__A
timestamp 1604681595
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_167
timestamp 1604681595
transform 1 0 16468 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 2760 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 2576 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_10
timestamp 1604681595
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_14
timestamp 1604681595
transform 1 0 2392 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1604681595
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1604681595
transform 1 0 3496 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_22
timestamp 1604681595
transform 1 0 3128 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3680 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 3312 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_36
timestamp 1604681595
transform 1 0 4416 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4508 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4692 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_58
timestamp 1604681595
transform 1 0 6440 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_64
timestamp 1604681595
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_71
timestamp 1604681595
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_88
timestamp 1604681595
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_116
timestamp 1604681595
transform 1 0 11776 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13156 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14168 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_126
timestamp 1604681595
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_130
timestamp 1604681595
transform 1 0 13064 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_140
timestamp 1604681595
transform 1 0 13984 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_144
timestamp 1604681595
transform 1 0 14352 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1604681595
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_163
timestamp 1604681595
transform 1 0 16100 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_175
timestamp 1604681595
transform 1 0 17204 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1604681595
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1604681595
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_211
timestamp 1604681595
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604681595
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604681595
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_11
timestamp 1604681595
transform 1 0 2116 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_10
timestamp 1604681595
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_18
timestamp 1604681595
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_14
timestamp 1604681595
transform 1 0 2392 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 2668 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 2944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2576 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 2852 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_23
timestamp 1604681595
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_22
timestamp 1604681595
transform 1 0 3128 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_36
timestamp 1604681595
transform 1 0 4416 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4600 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3680 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_34_51
timestamp 1604681595
transform 1 0 5796 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1604681595
transform 1 0 5428 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_47
timestamp 1604681595
transform 1 0 5428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 5888 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_54
timestamp 1604681595
transform 1 0 6072 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_55
timestamp 1604681595
transform 1 0 6164 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6716 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8648 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_81
timestamp 1604681595
transform 1 0 8556 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_84
timestamp 1604681595
transform 1 0 8832 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_88
timestamp 1604681595
transform 1 0 9200 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_85
timestamp 1604681595
transform 1 0 8924 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9568 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_101
timestamp 1604681595
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10028 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_33_109
timestamp 1604681595
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_105
timestamp 1604681595
transform 1 0 10764 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10948 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 11316 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_116
timestamp 1604681595
transform 1 0 11776 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 12512 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_127
timestamp 1604681595
transform 1 0 12788 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_133
timestamp 1604681595
transform 1 0 13340 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_129
timestamp 1604681595
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_137
timestamp 1604681595
transform 1 0 13708 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_137
timestamp 1604681595
transform 1 0 13708 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14260 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13800 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1604681595
transform 1 0 16284 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_157
timestamp 1604681595
transform 1 0 15548 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_157
timestamp 1604681595
transform 1 0 15548 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1604681595
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_180
timestamp 1604681595
transform 1 0 17664 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_169
timestamp 1604681595
transform 1 0 16652 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_181
timestamp 1604681595
transform 1 0 17756 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_193
timestamp 1604681595
transform 1 0 18860 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_205
timestamp 1604681595
transform 1 0 19964 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1604681595
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2852 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 2668 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_10
timestamp 1604681595
transform 1 0 2024 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_38
timestamp 1604681595
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_42
timestamp 1604681595
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 5336 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_50
timestamp 1604681595
transform 1 0 5704 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1604681595
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_58
timestamp 1604681595
transform 1 0 6440 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7452 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8464 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_66
timestamp 1604681595
transform 1 0 7176 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_78
timestamp 1604681595
transform 1 0 8280 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_82
timestamp 1604681595
transform 1 0 8648 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9476 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10488 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_86
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_100
timestamp 1604681595
transform 1 0 10304 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_104
timestamp 1604681595
transform 1 0 10672 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10856 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_114
timestamp 1604681595
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1604681595
transform 1 0 12696 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 13708 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13156 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13524 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_129
timestamp 1604681595
transform 1 0 12972 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_133
timestamp 1604681595
transform 1 0 13340 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604681595
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604681595
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_180
timestamp 1604681595
transform 1 0 17664 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1604681595
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 2760 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2576 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_10
timestamp 1604681595
transform 1 0 2024 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_14
timestamp 1604681595
transform 1 0 2392 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 3312 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_22
timestamp 1604681595
transform 1 0 3128 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_26
timestamp 1604681595
transform 1 0 3496 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_41
timestamp 1604681595
transform 1 0 4876 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 5520 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5888 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_46
timestamp 1604681595
transform 1 0 5336 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_50
timestamp 1604681595
transform 1 0 5704 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_54
timestamp 1604681595
transform 1 0 6072 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_65
timestamp 1604681595
transform 1 0 7084 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_71
timestamp 1604681595
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1604681595
transform 1 0 8648 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10212 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_86
timestamp 1604681595
transform 1 0 9016 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_118
timestamp 1604681595
transform 1 0 11960 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_124
timestamp 1604681595
transform 1 0 12512 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13800 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14168 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_136
timestamp 1604681595
transform 1 0 13616 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_140
timestamp 1604681595
transform 1 0 13984 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_144
timestamp 1604681595
transform 1 0 14352 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1604681595
transform 1 0 16284 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_152
timestamp 1604681595
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_157
timestamp 1604681595
transform 1 0 15548 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1604681595
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_180
timestamp 1604681595
transform 1 0 17664 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_192
timestamp 1604681595
transform 1 0 18768 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_204
timestamp 1604681595
transform 1 0 19872 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_212
timestamp 1604681595
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604681595
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2760 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2208 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_10
timestamp 1604681595
transform 1 0 2024 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_14
timestamp 1604681595
transform 1 0 2392 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_31
timestamp 1604681595
transform 1 0 3956 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1604681595
transform 1 0 4232 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_40
timestamp 1604681595
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1604681595
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604681595
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7176 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6992 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9476 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9108 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_85
timestamp 1604681595
transform 1 0 8924 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_89
timestamp 1604681595
transform 1 0 9292 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_93
timestamp 1604681595
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_106
timestamp 1604681595
transform 1 0 10856 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_110
timestamp 1604681595
transform 1 0 11224 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1604681595
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13708 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_126
timestamp 1604681595
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_130
timestamp 1604681595
transform 1 0 13064 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_134
timestamp 1604681595
transform 1 0 13432 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15640 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_156
timestamp 1604681595
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_160
timestamp 1604681595
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_164
timestamp 1604681595
transform 1 0 16192 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_176
timestamp 1604681595
transform 1 0 17296 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_182
timestamp 1604681595
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__90__A
timestamp 1604681595
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_196
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_201
timestamp 1604681595
transform 1 0 19596 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_213
timestamp 1604681595
transform 1 0 20700 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1604681595
transform 1 0 21804 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_237
timestamp 1604681595
transform 1 0 22908 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_243
timestamp 1604681595
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1604681595
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 2852 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_11
timestamp 1604681595
transform 1 0 2116 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_23
timestamp 1604681595
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_51
timestamp 1604681595
transform 1 0 5796 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7084 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6900 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10028 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_84
timestamp 1604681595
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_116
timestamp 1604681595
transform 1 0 11776 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12696 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_38_145
timestamp 1604681595
transform 1 0 14444 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_173
timestamp 1604681595
transform 1 0 17020 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_185
timestamp 1604681595
transform 1 0 18124 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _90_
timestamp 1604681595
transform 1 0 19412 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1604681595
transform 1 0 19228 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_203
timestamp 1604681595
transform 1 0 19780 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_211
timestamp 1604681595
transform 1 0 20516 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1604681595
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1604681595
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_251
timestamp 1604681595
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1604681595
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_11
timestamp 1604681595
transform 1 0 2116 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_17
timestamp 1604681595
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_13
timestamp 1604681595
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 2852 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_23
timestamp 1604681595
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_25
timestamp 1604681595
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_21
timestamp 1604681595
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_36
timestamp 1604681595
transform 1 0 4416 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4784 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 3772 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_40_42
timestamp 1604681595
transform 1 0 4968 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_52
timestamp 1604681595
transform 1 0 5888 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_48
timestamp 1604681595
transform 1 0 5520 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5704 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_56
timestamp 1604681595
transform 1 0 6256 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6072 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_31.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_40_67
timestamp 1604681595
transform 1 0 7268 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_63
timestamp 1604681595
transform 1 0 6900 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_68
timestamp 1604681595
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 7084 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7452 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7544 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7636 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7728 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10120 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10212 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9936 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_91
timestamp 1604681595
transform 1 0 9476 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_95
timestamp 1604681595
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_112
timestamp 1604681595
transform 1 0 11408 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_108
timestamp 1604681595
transform 1 0 11040 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_117
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12604 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1604681595
transform 1 0 14168 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12880 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 13616 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_127
timestamp 1604681595
transform 1 0 12788 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_134
timestamp 1604681595
transform 1 0 13432 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_138
timestamp 1604681595
transform 1 0 13800 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_145
timestamp 1604681595
transform 1 0 14444 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _98_
timestamp 1604681595
transform 1 0 15364 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__98__A
timestamp 1604681595
transform 1 0 15916 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__95__A
timestamp 1604681595
transform 1 0 16284 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_147
timestamp 1604681595
transform 1 0 14628 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_159
timestamp 1604681595
transform 1 0 15732 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_163
timestamp 1604681595
transform 1 0 16100 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_172
timestamp 1604681595
transform 1 0 16928 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_175
timestamp 1604681595
transform 1 0 17204 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_171
timestamp 1604681595
transform 1 0 16836 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__96__A
timestamp 1604681595
transform 1 0 17020 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _96_
timestamp 1604681595
transform 1 0 16468 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _95_
timestamp 1604681595
transform 1 0 16560 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_184
timestamp 1604681595
transform 1 0 18032 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_182
timestamp 1604681595
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_179
timestamp 1604681595
transform 1 0 17572 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__94__A
timestamp 1604681595
transform 1 0 17664 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _94_
timestamp 1604681595
transform 1 0 17664 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _93_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_192
timestamp 1604681595
transform 1 0 18768 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_192
timestamp 1604681595
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_188
timestamp 1604681595
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__91__A
timestamp 1604681595
transform 1 0 18952 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__93__A
timestamp 1604681595
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _92_
timestamp 1604681595
transform 1 0 19136 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _91_
timestamp 1604681595
transform 1 0 18860 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_204
timestamp 1604681595
transform 1 0 19872 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_200
timestamp 1604681595
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__92__A
timestamp 1604681595
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _89_
timestamp 1604681595
transform 1 0 20240 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1604681595
transform 1 0 19228 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1604681595
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1604681595
transform 1 0 20332 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_216
timestamp 1604681595
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_212
timestamp 1604681595
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__88__A
timestamp 1604681595
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__89__A
timestamp 1604681595
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_224
timestamp 1604681595
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__87__A
timestamp 1604681595
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_219
timestamp 1604681595
transform 1 0 21252 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_228
timestamp 1604681595
transform 1 0 22080 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_231
timestamp 1604681595
transform 1 0 22356 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_243
timestamp 1604681595
transform 1 0 23460 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1604681595
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1604681595
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_255
timestamp 1604681595
transform 1 0 24564 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_267
timestamp 1604681595
transform 1 0 25668 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 2668 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1604681595
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1604681595
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_19
timestamp 1604681595
transform 1 0 2852 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3404 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_34
timestamp 1604681595
transform 1 0 4232 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_38
timestamp 1604681595
transform 1 0 4600 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_42
timestamp 1604681595
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_53
timestamp 1604681595
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604681595
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7728 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 7360 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 8464 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_66
timestamp 1604681595
transform 1 0 7176 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_70
timestamp 1604681595
transform 1 0 7544 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_78
timestamp 1604681595
transform 1 0 8280 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_82
timestamp 1604681595
transform 1 0 8648 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10672 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10488 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 9752 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 8832 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_90
timestamp 1604681595
transform 1 0 9384 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_96
timestamp 1604681595
transform 1 0 9936 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_100
timestamp 1604681595
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_113
timestamp 1604681595
transform 1 0 11500 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_132
timestamp 1604681595
transform 1 0 13248 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_144
timestamp 1604681595
transform 1 0 14352 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_156
timestamp 1604681595
transform 1 0 15456 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_168
timestamp 1604681595
transform 1 0 16560 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_180
timestamp 1604681595
transform 1 0 17664 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_7
timestamp 1604681595
transform 1 0 1748 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_19
timestamp 1604681595
transform 1 0 2852 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4784 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5796 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_49
timestamp 1604681595
transform 1 0 5612 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_53
timestamp 1604681595
transform 1 0 5980 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_61
timestamp 1604681595
transform 1 0 6716 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 8556 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_67
timestamp 1604681595
transform 1 0 7268 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_79
timestamp 1604681595
transform 1 0 8372 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_83
timestamp 1604681595
transform 1 0 8740 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10672 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_91
timestamp 1604681595
transform 1 0 9476 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_98
timestamp 1604681595
transform 1 0 10120 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1604681595
transform 1 0 11132 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_121
timestamp 1604681595
transform 1 0 12236 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_128
timestamp 1604681595
transform 1 0 12880 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_140
timestamp 1604681595
transform 1 0 13984 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_152
timestamp 1604681595
transform 1 0 15088 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 13910 0 13966 480 6 ccff_head
port 0 nsew default input
rlabel metal2 s 23202 0 23258 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 16056 480 16176 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 22720 480 22840 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 23400 480 23520 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 23944 480 24064 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 24624 480 24744 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 25168 480 25288 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 26392 480 26512 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 27616 480 27736 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 11058 27520 11114 28000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 11702 27520 11758 28000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 12806 27520 12862 28000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 13358 27520 13414 28000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15106 27520 15162 28000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15658 27520 15714 28000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 5354 27520 5410 28000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 5998 27520 6054 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 6550 27520 6606 28000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 8206 27520 8262 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 8850 27520 8906 28000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 9402 27520 9458 28000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 9954 27520 10010 28000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 16210 27520 16266 28000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 21914 27520 21970 28000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 23110 27520 23166 28000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 23662 27520 23718 28000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 16762 27520 16818 28000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 18510 27520 18566 28000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 19614 27520 19670 28000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 20258 27520 20314 28000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 20810 27520 20866 28000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 left_bottom_grid_pin_11_
port 82 nsew default input
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_1_
port 83 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_3_
port 84 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_5_
port 85 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_7_
port 86 nsew default input
rlabel metal3 s 0 2592 480 2712 6 left_bottom_grid_pin_9_
port 87 nsew default input
rlabel metal2 s 4618 0 4674 480 6 prog_clk
port 88 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_42_
port 89 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_43_
port 90 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_44_
port 91 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_45_
port 92 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_46_
port 93 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_47_
port 94 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 top_left_grid_pin_48_
port 95 nsew default input
rlabel metal2 s 4250 27520 4306 28000 6 top_left_grid_pin_49_
port 96 nsew default input
rlabel metal2 s 27618 27520 27674 28000 6 top_right_grid_pin_1_
port 97 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 98 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 99 nsew default input
<< properties >>
string FIXED_BBOX 0 0 27679 28000
<< end >>
